magic
tech gf180mcuD
magscale 1 5
timestamp 1701904170
<< obsm1 >>
rect 672 1538 279328 174078
<< metal2 >>
rect 27888 0 27944 400
rect 83888 0 83944 400
rect 139888 0 139944 400
rect 195888 0 195944 400
rect 251888 0 251944 400
<< obsm2 >>
rect 854 430 279146 174067
rect 854 400 27858 430
rect 27974 400 83858 430
rect 83974 400 139858 430
rect 139974 400 195858 430
rect 195974 400 251858 430
rect 251974 400 279146 430
<< metal3 >>
rect 0 171696 400 171752
rect 279600 171696 280000 171752
rect 0 164416 400 164472
rect 279600 164416 280000 164472
rect 0 157136 400 157192
rect 279600 157136 280000 157192
rect 0 149856 400 149912
rect 279600 149856 280000 149912
rect 0 142576 400 142632
rect 279600 142576 280000 142632
rect 0 135296 400 135352
rect 279600 135296 280000 135352
rect 0 128016 400 128072
rect 279600 128016 280000 128072
rect 0 120736 400 120792
rect 279600 120736 280000 120792
rect 0 113456 400 113512
rect 279600 113456 280000 113512
rect 0 106176 400 106232
rect 279600 106176 280000 106232
rect 0 98896 400 98952
rect 279600 98896 280000 98952
rect 0 91616 400 91672
rect 279600 91616 280000 91672
rect 0 84336 400 84392
rect 279600 84336 280000 84392
rect 0 77056 400 77112
rect 279600 77056 280000 77112
rect 0 69776 400 69832
rect 279600 69776 280000 69832
rect 0 62496 400 62552
rect 279600 62496 280000 62552
rect 0 55216 400 55272
rect 279600 55216 280000 55272
rect 0 47936 400 47992
rect 279600 47936 280000 47992
rect 0 40656 400 40712
rect 279600 40656 280000 40712
rect 0 33376 400 33432
rect 279600 33376 280000 33432
rect 0 26096 400 26152
rect 279600 26096 280000 26152
rect 0 18816 400 18872
rect 279600 18816 280000 18872
rect 0 11536 400 11592
rect 279600 11536 280000 11592
rect 0 4256 400 4312
rect 279600 4256 280000 4312
<< obsm3 >>
rect 400 171782 279600 174062
rect 430 171666 279570 171782
rect 400 164502 279600 171666
rect 430 164386 279570 164502
rect 400 157222 279600 164386
rect 430 157106 279570 157222
rect 400 149942 279600 157106
rect 430 149826 279570 149942
rect 400 142662 279600 149826
rect 430 142546 279570 142662
rect 400 135382 279600 142546
rect 430 135266 279570 135382
rect 400 128102 279600 135266
rect 430 127986 279570 128102
rect 400 120822 279600 127986
rect 430 120706 279570 120822
rect 400 113542 279600 120706
rect 430 113426 279570 113542
rect 400 106262 279600 113426
rect 430 106146 279570 106262
rect 400 98982 279600 106146
rect 430 98866 279570 98982
rect 400 91702 279600 98866
rect 430 91586 279570 91702
rect 400 84422 279600 91586
rect 430 84306 279570 84422
rect 400 77142 279600 84306
rect 430 77026 279570 77142
rect 400 69862 279600 77026
rect 430 69746 279570 69862
rect 400 62582 279600 69746
rect 430 62466 279570 62582
rect 400 55302 279600 62466
rect 430 55186 279570 55302
rect 400 48022 279600 55186
rect 430 47906 279570 48022
rect 400 40742 279600 47906
rect 430 40626 279570 40742
rect 400 33462 279600 40626
rect 430 33346 279570 33462
rect 400 26182 279600 33346
rect 430 26066 279570 26182
rect 400 18902 279600 26066
rect 430 18786 279570 18902
rect 400 11622 279600 18786
rect 430 11506 279570 11622
rect 400 4342 279600 11506
rect 430 4226 279570 4342
rect 400 1554 279600 4226
<< metal4 >>
rect 2224 1538 2384 174078
rect 9904 1538 10064 174078
rect 17584 1538 17744 174078
rect 25264 1538 25424 174078
rect 32944 1538 33104 174078
rect 40624 1538 40784 174078
rect 48304 1538 48464 174078
rect 55984 1538 56144 174078
rect 63664 1538 63824 174078
rect 71344 1538 71504 174078
rect 79024 1538 79184 174078
rect 86704 1538 86864 174078
rect 94384 1538 94544 174078
rect 102064 1538 102224 174078
rect 109744 1538 109904 174078
rect 117424 1538 117584 174078
rect 125104 1538 125264 174078
rect 132784 1538 132944 174078
rect 140464 1538 140624 174078
rect 148144 1538 148304 174078
rect 155824 1538 155984 174078
rect 163504 1538 163664 174078
rect 171184 1538 171344 174078
rect 178864 1538 179024 174078
rect 186544 1538 186704 174078
rect 194224 1538 194384 174078
rect 201904 1538 202064 174078
rect 209584 1538 209744 174078
rect 217264 1538 217424 174078
rect 224944 1538 225104 174078
rect 232624 1538 232784 174078
rect 240304 1538 240464 174078
rect 247984 1538 248144 174078
rect 255664 1538 255824 174078
rect 263344 1538 263504 174078
rect 271024 1538 271184 174078
rect 278704 1538 278864 174078
<< labels >>
rlabel metal3 s 279600 4256 280000 4312 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 128016 400 128072 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 0 106176 400 106232 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 0 84336 400 84392 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 0 62496 400 62552 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 0 40656 400 40712 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 0 18816 400 18872 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 279600 26096 280000 26152 6 io_in[1]
port 8 nsew signal input
rlabel metal3 s 279600 47936 280000 47992 6 io_in[2]
port 9 nsew signal input
rlabel metal3 s 279600 69776 280000 69832 6 io_in[3]
port 10 nsew signal input
rlabel metal3 s 279600 91616 280000 91672 6 io_in[4]
port 11 nsew signal input
rlabel metal3 s 279600 113456 280000 113512 6 io_in[5]
port 12 nsew signal input
rlabel metal3 s 279600 135296 280000 135352 6 io_in[6]
port 13 nsew signal input
rlabel metal3 s 279600 157136 280000 157192 6 io_in[7]
port 14 nsew signal input
rlabel metal3 s 0 171696 400 171752 6 io_in[8]
port 15 nsew signal input
rlabel metal3 s 0 149856 400 149912 6 io_in[9]
port 16 nsew signal input
rlabel metal3 s 279600 18816 280000 18872 6 io_oeb[0]
port 17 nsew signal output
rlabel metal3 s 0 113456 400 113512 6 io_oeb[10]
port 18 nsew signal output
rlabel metal3 s 0 91616 400 91672 6 io_oeb[11]
port 19 nsew signal output
rlabel metal3 s 0 69776 400 69832 6 io_oeb[12]
port 20 nsew signal output
rlabel metal3 s 0 47936 400 47992 6 io_oeb[13]
port 21 nsew signal output
rlabel metal3 s 0 26096 400 26152 6 io_oeb[14]
port 22 nsew signal output
rlabel metal3 s 0 4256 400 4312 6 io_oeb[15]
port 23 nsew signal output
rlabel metal3 s 279600 40656 280000 40712 6 io_oeb[1]
port 24 nsew signal output
rlabel metal3 s 279600 62496 280000 62552 6 io_oeb[2]
port 25 nsew signal output
rlabel metal3 s 279600 84336 280000 84392 6 io_oeb[3]
port 26 nsew signal output
rlabel metal3 s 279600 106176 280000 106232 6 io_oeb[4]
port 27 nsew signal output
rlabel metal3 s 279600 128016 280000 128072 6 io_oeb[5]
port 28 nsew signal output
rlabel metal3 s 279600 149856 280000 149912 6 io_oeb[6]
port 29 nsew signal output
rlabel metal3 s 279600 171696 280000 171752 6 io_oeb[7]
port 30 nsew signal output
rlabel metal3 s 0 157136 400 157192 6 io_oeb[8]
port 31 nsew signal output
rlabel metal3 s 0 135296 400 135352 6 io_oeb[9]
port 32 nsew signal output
rlabel metal3 s 279600 11536 280000 11592 6 io_out[0]
port 33 nsew signal output
rlabel metal3 s 0 120736 400 120792 6 io_out[10]
port 34 nsew signal output
rlabel metal3 s 0 98896 400 98952 6 io_out[11]
port 35 nsew signal output
rlabel metal3 s 0 77056 400 77112 6 io_out[12]
port 36 nsew signal output
rlabel metal3 s 0 55216 400 55272 6 io_out[13]
port 37 nsew signal output
rlabel metal3 s 0 33376 400 33432 6 io_out[14]
port 38 nsew signal output
rlabel metal3 s 0 11536 400 11592 6 io_out[15]
port 39 nsew signal output
rlabel metal3 s 279600 33376 280000 33432 6 io_out[1]
port 40 nsew signal output
rlabel metal3 s 279600 55216 280000 55272 6 io_out[2]
port 41 nsew signal output
rlabel metal3 s 279600 77056 280000 77112 6 io_out[3]
port 42 nsew signal output
rlabel metal3 s 279600 98896 280000 98952 6 io_out[4]
port 43 nsew signal output
rlabel metal3 s 279600 120736 280000 120792 6 io_out[5]
port 44 nsew signal output
rlabel metal3 s 279600 142576 280000 142632 6 io_out[6]
port 45 nsew signal output
rlabel metal3 s 279600 164416 280000 164472 6 io_out[7]
port 46 nsew signal output
rlabel metal3 s 0 164416 400 164472 6 io_out[8]
port 47 nsew signal output
rlabel metal3 s 0 142576 400 142632 6 io_out[9]
port 48 nsew signal output
rlabel metal2 s 139888 0 139944 400 6 irq[0]
port 49 nsew signal output
rlabel metal2 s 195888 0 195944 400 6 irq[1]
port 50 nsew signal output
rlabel metal2 s 251888 0 251944 400 6 irq[2]
port 51 nsew signal output
rlabel metal4 s 2224 1538 2384 174078 6 vdd
port 52 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 174078 6 vdd
port 52 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 174078 6 vdd
port 52 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 174078 6 vdd
port 52 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 174078 6 vdd
port 52 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 174078 6 vdd
port 52 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 174078 6 vdd
port 52 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 174078 6 vdd
port 52 nsew power bidirectional
rlabel metal4 s 125104 1538 125264 174078 6 vdd
port 52 nsew power bidirectional
rlabel metal4 s 140464 1538 140624 174078 6 vdd
port 52 nsew power bidirectional
rlabel metal4 s 155824 1538 155984 174078 6 vdd
port 52 nsew power bidirectional
rlabel metal4 s 171184 1538 171344 174078 6 vdd
port 52 nsew power bidirectional
rlabel metal4 s 186544 1538 186704 174078 6 vdd
port 52 nsew power bidirectional
rlabel metal4 s 201904 1538 202064 174078 6 vdd
port 52 nsew power bidirectional
rlabel metal4 s 217264 1538 217424 174078 6 vdd
port 52 nsew power bidirectional
rlabel metal4 s 232624 1538 232784 174078 6 vdd
port 52 nsew power bidirectional
rlabel metal4 s 247984 1538 248144 174078 6 vdd
port 52 nsew power bidirectional
rlabel metal4 s 263344 1538 263504 174078 6 vdd
port 52 nsew power bidirectional
rlabel metal4 s 278704 1538 278864 174078 6 vdd
port 52 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 174078 6 vss
port 53 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 174078 6 vss
port 53 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 174078 6 vss
port 53 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 174078 6 vss
port 53 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 174078 6 vss
port 53 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 174078 6 vss
port 53 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 174078 6 vss
port 53 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 174078 6 vss
port 53 nsew ground bidirectional
rlabel metal4 s 132784 1538 132944 174078 6 vss
port 53 nsew ground bidirectional
rlabel metal4 s 148144 1538 148304 174078 6 vss
port 53 nsew ground bidirectional
rlabel metal4 s 163504 1538 163664 174078 6 vss
port 53 nsew ground bidirectional
rlabel metal4 s 178864 1538 179024 174078 6 vss
port 53 nsew ground bidirectional
rlabel metal4 s 194224 1538 194384 174078 6 vss
port 53 nsew ground bidirectional
rlabel metal4 s 209584 1538 209744 174078 6 vss
port 53 nsew ground bidirectional
rlabel metal4 s 224944 1538 225104 174078 6 vss
port 53 nsew ground bidirectional
rlabel metal4 s 240304 1538 240464 174078 6 vss
port 53 nsew ground bidirectional
rlabel metal4 s 255664 1538 255824 174078 6 vss
port 53 nsew ground bidirectional
rlabel metal4 s 271024 1538 271184 174078 6 vss
port 53 nsew ground bidirectional
rlabel metal2 s 27888 0 27944 400 6 wb_clk_i
port 54 nsew signal input
rlabel metal2 s 83888 0 83944 400 6 wb_rst_i
port 55 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 280000 176000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 14848882
string GDS_FILE /home/gonsolo/work/caravel/gfmpw1/openlane/user_proj_example/runs/23_12_07_00_06/results/signoff/user_proj_example.magic.gds
string GDS_START 51278
<< end >>

