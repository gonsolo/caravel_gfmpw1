magic
tech gf180mcuD
magscale 1 5
timestamp 1701904763
<< metal2 >>
rect 5516 297780 5628 298500
rect 16548 297780 16660 298500
rect 27580 297780 27692 298500
rect 38612 297780 38724 298500
rect 49644 297780 49756 298500
rect 60676 297780 60788 298500
rect 71708 297780 71820 298500
rect 82740 297780 82852 298500
rect 93772 297780 93884 298500
rect 104804 297780 104916 298500
rect 115836 297780 115948 298500
rect 126868 297780 126980 298500
rect 137900 297780 138012 298500
rect 148932 297780 149044 298500
rect 159964 297780 160076 298500
rect 170996 297780 171108 298500
rect 182028 297780 182140 298500
rect 193060 297780 193172 298500
rect 204092 297780 204204 298500
rect 215124 297780 215236 298500
rect 226156 297780 226268 298500
rect 237188 297780 237300 298500
rect 248220 297780 248332 298500
rect 259252 297780 259364 298500
rect 270284 297780 270396 298500
rect 281316 297780 281428 298500
rect 292348 297780 292460 298500
rect 5782 240 5866 266
rect 5684 238 5866 240
rect 5684 196 5810 238
rect 5684 -480 5796 196
rect 5838 42 5866 238
rect 6566 240 6650 266
rect 6566 238 6748 240
rect 6566 98 6594 238
rect 6622 196 6748 238
rect 6566 65 6594 70
rect 5838 9 5866 14
rect 6636 -480 6748 196
rect 7588 -480 7700 240
rect 8540 -480 8652 240
rect 9492 -480 9604 240
rect 10444 -480 10556 240
rect 11396 -480 11508 240
rect 12348 -480 12460 240
rect 13300 -480 13412 240
rect 14252 -480 14364 240
rect 15204 -480 15316 240
rect 16156 -480 16268 240
rect 17108 -480 17220 240
rect 18060 -480 18172 240
rect 19012 -480 19124 240
rect 19964 -480 20076 240
rect 20916 -480 21028 240
rect 21868 -480 21980 240
rect 22820 -480 22932 240
rect 23772 -480 23884 240
rect 24724 -480 24836 240
rect 25676 -480 25788 240
rect 26628 -480 26740 240
rect 27580 -480 27692 240
rect 28532 -480 28644 240
rect 29484 -480 29596 240
rect 30436 -480 30548 240
rect 31388 -480 31500 240
rect 32340 -480 32452 240
rect 33292 -480 33404 240
rect 33894 42 33922 1540
rect 33894 9 33922 14
rect 34244 -480 34356 240
rect 35196 -480 35308 240
rect 36148 -480 36260 240
rect 37100 -480 37212 240
rect 38052 -480 38164 240
rect 39004 -480 39116 240
rect 39956 -480 40068 240
rect 40908 -480 41020 240
rect 41860 -480 41972 240
rect 42812 -480 42924 240
rect 43764 -480 43876 240
rect 44716 -480 44828 240
rect 45668 -480 45780 240
rect 46620 -480 46732 240
rect 47572 -480 47684 240
rect 48524 -480 48636 240
rect 49476 -480 49588 240
rect 50428 -480 50540 240
rect 51380 -480 51492 240
rect 52332 -480 52444 240
rect 53284 -480 53396 240
rect 54236 -480 54348 240
rect 55188 -480 55300 240
rect 56140 -480 56252 240
rect 57092 -480 57204 240
rect 58044 -480 58156 240
rect 58996 -480 59108 240
rect 59948 -480 60060 240
rect 60900 -480 61012 240
rect 61852 -480 61964 240
rect 62804 -480 62916 240
rect 63756 -480 63868 240
rect 64708 -480 64820 240
rect 65660 -480 65772 240
rect 66612 -480 66724 240
rect 67564 -480 67676 240
rect 68516 -480 68628 240
rect 69468 -480 69580 240
rect 70420 -480 70532 240
rect 71372 -480 71484 240
rect 72324 -480 72436 240
rect 73276 -480 73388 240
rect 74228 -480 74340 240
rect 75180 -480 75292 240
rect 76132 -480 76244 240
rect 77084 -480 77196 240
rect 78036 -480 78148 240
rect 78988 -480 79100 240
rect 79940 -480 80052 240
rect 80892 -480 81004 240
rect 81844 -480 81956 240
rect 82796 -480 82908 240
rect 83748 -480 83860 240
rect 84700 -480 84812 240
rect 85652 -480 85764 240
rect 86604 -480 86716 240
rect 87556 -480 87668 240
rect 88508 -480 88620 240
rect 89460 -480 89572 240
rect 89894 98 89922 1540
rect 89894 65 89922 70
rect 90412 -480 90524 240
rect 91364 -480 91476 240
rect 92316 -480 92428 240
rect 93268 -480 93380 240
rect 94220 -480 94332 240
rect 95172 -480 95284 240
rect 96124 -480 96236 240
rect 97076 -480 97188 240
rect 98028 -480 98140 240
rect 98980 -480 99092 240
rect 99932 -480 100044 240
rect 100884 -480 100996 240
rect 101836 -480 101948 240
rect 102788 -480 102900 240
rect 103740 -480 103852 240
rect 104692 -480 104804 240
rect 105644 -480 105756 240
rect 106596 -480 106708 240
rect 107548 -480 107660 240
rect 108500 -480 108612 240
rect 109452 -480 109564 240
rect 110404 -480 110516 240
rect 111356 -480 111468 240
rect 112308 -480 112420 240
rect 113260 -480 113372 240
rect 114212 -480 114324 240
rect 115164 -480 115276 240
rect 116116 -480 116228 240
rect 117068 -480 117180 240
rect 118020 -480 118132 240
rect 118972 -480 119084 240
rect 119924 -480 120036 240
rect 120876 -480 120988 240
rect 121828 -480 121940 240
rect 122780 -480 122892 240
rect 123732 -480 123844 240
rect 124684 -480 124796 240
rect 125636 -480 125748 240
rect 126588 -480 126700 240
rect 127540 -480 127652 240
rect 128492 -480 128604 240
rect 129444 -480 129556 240
rect 130396 -480 130508 240
rect 131348 -480 131460 240
rect 132300 -480 132412 240
rect 133252 -480 133364 240
rect 134204 -480 134316 240
rect 135156 -480 135268 240
rect 136108 -480 136220 240
rect 137060 -480 137172 240
rect 138012 -480 138124 240
rect 138964 -480 139076 240
rect 139916 -480 140028 240
rect 140868 -480 140980 240
rect 141820 -480 141932 240
rect 142772 -480 142884 240
rect 143724 -480 143836 240
rect 144676 -480 144788 240
rect 145628 -480 145740 240
rect 145894 42 145922 1540
rect 201908 1526 202258 1554
rect 145894 9 145922 14
rect 146580 -480 146692 240
rect 147532 -480 147644 240
rect 148484 -480 148596 240
rect 149436 -480 149548 240
rect 150388 -480 150500 240
rect 151340 -480 151452 240
rect 152292 -480 152404 240
rect 153244 -480 153356 240
rect 154196 -480 154308 240
rect 155148 -480 155260 240
rect 156100 -480 156212 240
rect 157052 -480 157164 240
rect 158004 -480 158116 240
rect 158956 -480 159068 240
rect 159908 -480 160020 240
rect 160860 -480 160972 240
rect 161812 -480 161924 240
rect 162764 -480 162876 240
rect 163716 -480 163828 240
rect 164668 -480 164780 240
rect 165620 -480 165732 240
rect 166572 -480 166684 240
rect 167524 -480 167636 240
rect 168476 -480 168588 240
rect 169428 -480 169540 240
rect 170380 -480 170492 240
rect 171332 -480 171444 240
rect 172284 -480 172396 240
rect 173236 -480 173348 240
rect 174188 -480 174300 240
rect 175140 -480 175252 240
rect 176092 -480 176204 240
rect 177044 -480 177156 240
rect 177996 -480 178108 240
rect 178948 -480 179060 240
rect 179900 -480 180012 240
rect 180852 -480 180964 240
rect 181804 -480 181916 240
rect 182756 -480 182868 240
rect 183708 -480 183820 240
rect 184660 -480 184772 240
rect 185612 -480 185724 240
rect 186564 -480 186676 240
rect 187516 -480 187628 240
rect 188468 -480 188580 240
rect 189420 -480 189532 240
rect 190372 -480 190484 240
rect 191324 -480 191436 240
rect 192276 -480 192388 240
rect 193228 -480 193340 240
rect 194180 -480 194292 240
rect 195132 -480 195244 240
rect 196084 -480 196196 240
rect 197036 -480 197148 240
rect 197988 -480 198100 240
rect 198940 -480 199052 240
rect 199892 -480 200004 240
rect 200844 -480 200956 240
rect 201796 -480 201908 240
rect 202230 98 202258 1526
rect 202230 65 202258 70
rect 202748 -480 202860 240
rect 203700 -480 203812 240
rect 204652 -480 204764 240
rect 205604 -480 205716 240
rect 206556 -480 206668 240
rect 207508 -480 207620 240
rect 208460 -480 208572 240
rect 209412 -480 209524 240
rect 210364 -480 210476 240
rect 211316 -480 211428 240
rect 212268 -480 212380 240
rect 213220 -480 213332 240
rect 214172 -480 214284 240
rect 215124 -480 215236 240
rect 216076 -480 216188 240
rect 217028 -480 217140 240
rect 217980 -480 218092 240
rect 218932 -480 219044 240
rect 219884 -480 219996 240
rect 220836 -480 220948 240
rect 221788 -480 221900 240
rect 222740 -480 222852 240
rect 223692 -480 223804 240
rect 224644 -480 224756 240
rect 225596 -480 225708 240
rect 226548 -480 226660 240
rect 227500 -480 227612 240
rect 228452 -480 228564 240
rect 229404 -480 229516 240
rect 230356 -480 230468 240
rect 231308 -480 231420 240
rect 232260 -480 232372 240
rect 233212 -480 233324 240
rect 234164 -480 234276 240
rect 235116 -480 235228 240
rect 236068 -480 236180 240
rect 237020 -480 237132 240
rect 237972 -480 238084 240
rect 238924 -480 239036 240
rect 239876 -480 239988 240
rect 240828 -480 240940 240
rect 241780 -480 241892 240
rect 242732 -480 242844 240
rect 243684 -480 243796 240
rect 244636 -480 244748 240
rect 245588 -480 245700 240
rect 246540 -480 246652 240
rect 247492 -480 247604 240
rect 248444 -480 248556 240
rect 249396 -480 249508 240
rect 250348 -480 250460 240
rect 251300 -480 251412 240
rect 252252 -480 252364 240
rect 253204 -480 253316 240
rect 254156 -480 254268 240
rect 255108 -480 255220 240
rect 256060 -480 256172 240
rect 257012 -480 257124 240
rect 257894 154 257922 1540
rect 290262 240 290346 266
rect 291214 240 291298 266
rect 292166 240 292250 266
rect 257894 121 257922 126
rect 257964 -480 258076 240
rect 258916 -480 259028 240
rect 259868 -480 259980 240
rect 260820 -480 260932 240
rect 261772 -480 261884 240
rect 262724 -480 262836 240
rect 263676 -480 263788 240
rect 264628 -480 264740 240
rect 265580 -480 265692 240
rect 266532 -480 266644 240
rect 267484 -480 267596 240
rect 268436 -480 268548 240
rect 269388 -480 269500 240
rect 270340 -480 270452 240
rect 271292 -480 271404 240
rect 272244 -480 272356 240
rect 273196 -480 273308 240
rect 274148 -480 274260 240
rect 275100 -480 275212 240
rect 276052 -480 276164 240
rect 277004 -480 277116 240
rect 277956 -480 278068 240
rect 278908 -480 279020 240
rect 279860 -480 279972 240
rect 280812 -480 280924 240
rect 281764 -480 281876 240
rect 282716 -480 282828 240
rect 283668 -480 283780 240
rect 284620 -480 284732 240
rect 285572 -480 285684 240
rect 286524 -480 286636 240
rect 287476 -480 287588 240
rect 288428 -480 288540 240
rect 289380 -480 289492 240
rect 290262 238 290444 240
rect 290262 42 290290 238
rect 290318 196 290444 238
rect 290262 9 290290 14
rect 290332 -480 290444 196
rect 291214 238 291396 240
rect 291214 98 291242 238
rect 291270 196 291396 238
rect 291214 65 291242 70
rect 291284 -480 291396 196
rect 292166 238 292348 240
rect 292166 154 292194 238
rect 292222 196 292348 238
rect 292166 121 292194 126
rect 292236 -480 292348 196
<< via2 >>
rect 6566 70 6594 98
rect 5838 14 5866 42
rect 33894 14 33922 42
rect 89894 70 89922 98
rect 145894 14 145922 42
rect 202230 70 202258 98
rect 257894 126 257922 154
rect 290262 14 290290 42
rect 291214 70 291242 98
rect 292166 126 292194 154
<< metal3 >>
rect 297780 294308 298500 294420
rect -480 293580 240 293692
rect 297780 287700 298500 287812
rect -480 286524 240 286636
rect 297780 281092 298500 281204
rect -480 279468 240 279580
rect 297780 274484 298500 274596
rect -480 272412 240 272524
rect 297780 267876 298500 267988
rect -480 265356 240 265468
rect 297780 261268 298500 261380
rect -480 258300 240 258412
rect 297780 254660 298500 254772
rect -480 251244 240 251356
rect 297780 248052 298500 248164
rect -480 244188 240 244300
rect 297780 241444 298500 241556
rect -480 237132 240 237244
rect 297780 234836 298500 234948
rect -480 230076 240 230188
rect 297780 228228 298500 228340
rect -480 223020 240 223132
rect 297780 221620 298500 221732
rect -480 215964 240 216076
rect 297780 215012 298500 215124
rect -480 208908 240 209020
rect 297780 208404 298500 208516
rect -480 201852 240 201964
rect 297780 201796 298500 201908
rect 297780 195188 298500 195300
rect -480 194796 240 194908
rect 297780 188580 298500 188692
rect -480 187740 240 187852
rect 297780 181972 298500 182084
rect -480 180684 240 180796
rect 297780 175364 298500 175476
rect -480 173628 240 173740
rect 3761 173222 3766 173250
rect 3794 173222 6020 173250
rect 285964 173222 287686 173250
rect 287714 173222 287719 173250
rect 297780 168756 298500 168868
rect 196 166684 3766 166698
rect -480 166670 3766 166684
rect 3794 166670 3799 166698
rect -480 166572 240 166670
rect 3761 165942 3766 165970
rect 3794 165942 6020 165970
rect 285964 165942 287742 165970
rect 287770 165942 287775 165970
rect 297780 162148 298500 162260
rect -480 159586 240 159628
rect -480 159558 3766 159586
rect 3794 159558 3799 159586
rect -480 159516 240 159558
rect 3761 158662 3766 158690
rect 3794 158662 6020 158690
rect 285964 158662 287798 158690
rect 287826 158662 287831 158690
rect 297780 155554 298500 155652
rect 287681 155526 287686 155554
rect 287714 155540 298500 155554
rect 287714 155526 297836 155540
rect 196 152572 3766 152586
rect -480 152558 3766 152572
rect 3794 152558 3799 152586
rect -480 152460 240 152558
rect 3761 151382 3766 151410
rect 3794 151382 6020 151410
rect 285964 151382 287686 151410
rect 287714 151382 287719 151410
rect 297780 148946 298500 149044
rect 287737 148918 287742 148946
rect 287770 148932 298500 148946
rect 287770 148918 297836 148932
rect 196 145516 3766 145530
rect -480 145502 3766 145516
rect 3794 145502 3799 145530
rect -480 145404 240 145502
rect 3761 144102 3766 144130
rect 3794 144102 6020 144130
rect 285964 144102 287742 144130
rect 287770 144102 287775 144130
rect 297780 142338 298500 142436
rect 287793 142310 287798 142338
rect 287826 142324 298500 142338
rect 287826 142310 297836 142324
rect 196 138460 3766 138474
rect -480 138446 3766 138460
rect 3794 138446 3799 138474
rect -480 138348 240 138446
rect 3089 136822 3094 136850
rect 3122 136822 6020 136850
rect 285964 136822 287798 136850
rect 287826 136822 287831 136850
rect 297780 135730 298500 135828
rect 287681 135702 287686 135730
rect 287714 135716 298500 135730
rect 287714 135702 297836 135716
rect 196 131404 3094 131418
rect -480 131390 3094 131404
rect 3122 131390 3127 131418
rect -480 131292 240 131390
rect 3761 129542 3766 129570
rect 3794 129542 6020 129570
rect 285964 129542 287686 129570
rect 287714 129542 287719 129570
rect 297780 129122 298500 129220
rect 287737 129094 287742 129122
rect 287770 129108 298500 129122
rect 287770 129094 297836 129108
rect -480 124306 240 124348
rect -480 124278 3766 124306
rect 3794 124278 3799 124306
rect -480 124236 240 124278
rect 297780 122514 298500 122612
rect 287793 122486 287798 122514
rect 287826 122500 298500 122514
rect 287826 122486 297836 122500
rect 3089 122262 3094 122290
rect 3122 122262 6020 122290
rect 285964 122262 287910 122290
rect 287938 122262 287943 122290
rect 196 117292 3094 117306
rect -480 117278 3094 117292
rect 3122 117278 3127 117306
rect -480 117180 240 117278
rect 297780 115962 298500 116004
rect 287681 115934 287686 115962
rect 287714 115934 298500 115962
rect 297780 115892 298500 115934
rect 2081 114982 2086 115010
rect 2114 114982 6020 115010
rect 285964 114982 287742 115010
rect 287770 114982 287775 115010
rect 196 110236 2086 110250
rect -480 110222 2086 110236
rect 2114 110222 2119 110250
rect -480 110124 240 110222
rect 297780 109298 298500 109396
rect 287905 109270 287910 109298
rect 287938 109284 298500 109298
rect 287938 109270 297836 109284
rect 3089 107702 3094 107730
rect 3122 107702 6020 107730
rect 285964 107702 287686 107730
rect 287714 107702 287719 107730
rect 196 103180 3094 103194
rect -480 103166 3094 103180
rect 3122 103166 3127 103194
rect -480 103068 240 103166
rect 297780 102690 298500 102788
rect 287737 102662 287742 102690
rect 287770 102676 298500 102690
rect 287770 102662 297836 102676
rect 2081 100422 2086 100450
rect 2114 100422 6020 100450
rect 285964 100422 287742 100450
rect 287770 100422 287775 100450
rect 196 96124 2086 96138
rect -480 96110 2086 96124
rect 2114 96110 2119 96138
rect -480 96012 240 96110
rect 297780 96082 298500 96180
rect 287681 96054 287686 96082
rect 287714 96068 298500 96082
rect 287714 96054 297836 96068
rect 2473 93142 2478 93170
rect 2506 93142 6020 93170
rect 285964 93142 287798 93170
rect 287826 93142 287831 93170
rect 297780 89474 298500 89572
rect 287737 89446 287742 89474
rect 287770 89460 298500 89474
rect 287770 89446 297836 89460
rect -480 89026 240 89068
rect -480 88998 2478 89026
rect 2506 88998 2511 89026
rect -480 88956 240 88998
rect 2081 85862 2086 85890
rect 2114 85862 6020 85890
rect 285964 85862 287686 85890
rect 287714 85862 287719 85890
rect 297780 82866 298500 82964
rect 287793 82838 287798 82866
rect 287826 82852 298500 82866
rect 287826 82838 297836 82852
rect 196 82012 2086 82026
rect -480 81998 2086 82012
rect 2114 81998 2119 82026
rect -480 81900 240 81998
rect 3761 78582 3766 78610
rect 3794 78582 6020 78610
rect 285964 78582 287742 78610
rect 287770 78582 287775 78610
rect 297780 76258 298500 76356
rect 287681 76230 287686 76258
rect 287714 76244 298500 76258
rect 287714 76230 297836 76244
rect 196 74956 3766 74970
rect -480 74942 3766 74956
rect 3794 74942 3799 74970
rect -480 74844 240 74942
rect 3761 71302 3766 71330
rect 3794 71302 6020 71330
rect 285964 71302 287798 71330
rect 287826 71302 287831 71330
rect 297780 69650 298500 69748
rect 287737 69622 287742 69650
rect 287770 69636 298500 69650
rect 287770 69622 297836 69636
rect 196 67900 3766 67914
rect -480 67886 3766 67900
rect 3794 67886 3799 67914
rect -480 67788 240 67886
rect 3369 64022 3374 64050
rect 3402 64022 6020 64050
rect 285964 64022 287686 64050
rect 287714 64022 287719 64050
rect 297780 63042 298500 63140
rect 287793 63014 287798 63042
rect 287826 63028 298500 63042
rect 287826 63014 297836 63028
rect 196 60844 3374 60858
rect -480 60830 3374 60844
rect 3402 60830 3407 60858
rect -480 60732 240 60830
rect 3369 56742 3374 56770
rect 3402 56742 6020 56770
rect 285964 56742 295246 56770
rect 295274 56742 295279 56770
rect 297780 56434 298500 56532
rect 287681 56406 287686 56434
rect 287714 56420 298500 56434
rect 287714 56406 297836 56420
rect -480 53746 240 53788
rect -480 53718 3374 53746
rect 3402 53718 3407 53746
rect -480 53676 240 53718
rect 295241 49910 295246 49938
rect 295274 49924 297836 49938
rect 295274 49910 298500 49924
rect 297780 49812 298500 49910
rect 3761 49462 3766 49490
rect 3794 49462 6020 49490
rect 285964 49462 293566 49490
rect 293594 49462 293599 49490
rect 196 46732 3766 46746
rect -480 46718 3766 46732
rect 3794 46718 3799 46746
rect -480 46620 240 46718
rect 297780 43218 298500 43316
rect 293561 43190 293566 43218
rect 293594 43204 298500 43218
rect 293594 43190 297836 43204
rect 3761 42182 3766 42210
rect 3794 42182 6020 42210
rect 285964 42182 293566 42210
rect 293594 42182 293599 42210
rect 196 39676 3766 39690
rect -480 39662 3766 39676
rect 3794 39662 3799 39690
rect -480 39564 240 39662
rect 297780 36610 298500 36708
rect 293561 36582 293566 36610
rect 293594 36596 298500 36610
rect 293594 36582 297836 36596
rect 3369 34902 3374 34930
rect 3402 34902 6020 34930
rect 285964 34902 293174 34930
rect 293202 34902 293207 34930
rect 196 32620 3374 32634
rect -480 32606 3374 32620
rect 3402 32606 3407 32634
rect -480 32508 240 32606
rect 297780 30002 298500 30100
rect 293169 29974 293174 30002
rect 293202 29988 298500 30002
rect 293202 29974 297836 29988
rect 2473 27622 2478 27650
rect 2506 27622 6020 27650
rect 285964 27622 293566 27650
rect 293594 27622 293599 27650
rect 196 25564 2478 25578
rect -480 25550 2478 25564
rect 2506 25550 2511 25578
rect -480 25452 240 25550
rect 297780 23394 298500 23492
rect 293561 23366 293566 23394
rect 293594 23380 298500 23394
rect 293594 23366 297836 23380
rect 3369 20342 3374 20370
rect 3402 20342 6020 20370
rect 285964 20342 293566 20370
rect 293594 20342 293599 20370
rect -480 18466 240 18508
rect -480 18438 3374 18466
rect 3402 18438 3407 18466
rect -480 18396 240 18438
rect 297780 16842 298500 16884
rect 293561 16814 293566 16842
rect 293594 16814 298500 16842
rect 297780 16772 298500 16814
rect 2081 13062 2086 13090
rect 2114 13062 6020 13090
rect 285964 13062 293566 13090
rect 293594 13062 293599 13090
rect 196 11452 2086 11466
rect -480 11438 2086 11452
rect 2114 11438 2119 11466
rect -480 11340 240 11438
rect 297780 10178 298500 10276
rect 293561 10150 293566 10178
rect 293594 10164 298500 10178
rect 293594 10150 297836 10164
rect 3369 5782 3374 5810
rect 3402 5782 6020 5810
rect 285964 5782 295638 5810
rect 295666 5782 295671 5810
rect 196 4396 3374 4410
rect -480 4382 3374 4396
rect 3402 4382 3407 4410
rect -480 4284 240 4382
rect 295633 3654 295638 3682
rect 295666 3668 297836 3682
rect 295666 3654 298500 3668
rect 297780 3556 298500 3654
rect 257889 126 257894 154
rect 257922 126 292166 154
rect 292194 126 292199 154
rect 6561 70 6566 98
rect 6594 70 89894 98
rect 89922 70 89927 98
rect 202225 70 202230 98
rect 202258 70 291214 98
rect 291242 70 291247 98
rect 5828 14 5838 42
rect 5866 14 33894 42
rect 33922 14 33927 42
rect 145889 14 145894 42
rect 145922 14 290262 42
rect 290290 14 290295 42
<< via3 >>
rect 3766 173222 3794 173250
rect 287686 173222 287714 173250
rect 3766 166670 3794 166698
rect 3766 165942 3794 165970
rect 287742 165942 287770 165970
rect 3766 159558 3794 159586
rect 3766 158662 3794 158690
rect 287798 158662 287826 158690
rect 287686 155526 287714 155554
rect 3766 152558 3794 152586
rect 3766 151382 3794 151410
rect 287686 151382 287714 151410
rect 287742 148918 287770 148946
rect 3766 145502 3794 145530
rect 3766 144102 3794 144130
rect 287742 144102 287770 144130
rect 287798 142310 287826 142338
rect 3766 138446 3794 138474
rect 3094 136822 3122 136850
rect 287798 136822 287826 136850
rect 287686 135702 287714 135730
rect 3094 131390 3122 131418
rect 3766 129542 3794 129570
rect 287686 129542 287714 129570
rect 287742 129094 287770 129122
rect 3766 124278 3794 124306
rect 287798 122486 287826 122514
rect 3094 122262 3122 122290
rect 287910 122262 287938 122290
rect 3094 117278 3122 117306
rect 287686 115934 287714 115962
rect 2086 114982 2114 115010
rect 287742 114982 287770 115010
rect 2086 110222 2114 110250
rect 287910 109270 287938 109298
rect 3094 107702 3122 107730
rect 287686 107702 287714 107730
rect 3094 103166 3122 103194
rect 287742 102662 287770 102690
rect 2086 100422 2114 100450
rect 287742 100422 287770 100450
rect 2086 96110 2114 96138
rect 287686 96054 287714 96082
rect 2478 93142 2506 93170
rect 287798 93142 287826 93170
rect 287742 89446 287770 89474
rect 2478 88998 2506 89026
rect 2086 85862 2114 85890
rect 287686 85862 287714 85890
rect 287798 82838 287826 82866
rect 2086 81998 2114 82026
rect 3766 78582 3794 78610
rect 287742 78582 287770 78610
rect 287686 76230 287714 76258
rect 3766 74942 3794 74970
rect 3766 71302 3794 71330
rect 287798 71302 287826 71330
rect 287742 69622 287770 69650
rect 3766 67886 3794 67914
rect 3374 64022 3402 64050
rect 287686 64022 287714 64050
rect 287798 63014 287826 63042
rect 3374 60830 3402 60858
rect 3374 56742 3402 56770
rect 295246 56742 295274 56770
rect 287686 56406 287714 56434
rect 3374 53718 3402 53746
rect 295246 49910 295274 49938
rect 3766 49462 3794 49490
rect 293566 49462 293594 49490
rect 3766 46718 3794 46746
rect 293566 43190 293594 43218
rect 3766 42182 3794 42210
rect 293566 42182 293594 42210
rect 3766 39662 3794 39690
rect 293566 36582 293594 36610
rect 3374 34902 3402 34930
rect 293174 34902 293202 34930
rect 3374 32606 3402 32634
rect 293174 29974 293202 30002
rect 2478 27622 2506 27650
rect 293566 27622 293594 27650
rect 2478 25550 2506 25578
rect 293566 23366 293594 23394
rect 3374 20342 3402 20370
rect 293566 20342 293594 20370
rect 3374 18438 3402 18466
rect 293566 16814 293594 16842
rect 2086 13062 2114 13090
rect 293566 13062 293594 13090
rect 2086 11438 2114 11466
rect 293566 10150 293594 10178
rect 3374 5782 3402 5810
rect 295638 5782 295666 5810
rect 3374 4382 3402 4410
rect 295638 3654 295666 3682
<< metal4 >>
rect -958 299086 -648 299134
rect -958 299058 -910 299086
rect -882 299058 -848 299086
rect -820 299058 -786 299086
rect -758 299058 -724 299086
rect -696 299058 -648 299086
rect -958 299024 -648 299058
rect -958 298996 -910 299024
rect -882 298996 -848 299024
rect -820 298996 -786 299024
rect -758 298996 -724 299024
rect -696 298996 -648 299024
rect -958 298962 -648 298996
rect -958 298934 -910 298962
rect -882 298934 -848 298962
rect -820 298934 -786 298962
rect -758 298934 -724 298962
rect -696 298934 -648 298962
rect -958 298900 -648 298934
rect -958 298872 -910 298900
rect -882 298872 -848 298900
rect -820 298872 -786 298900
rect -758 298872 -724 298900
rect -696 298872 -648 298900
rect -958 293175 -648 298872
rect -958 293147 -910 293175
rect -882 293147 -848 293175
rect -820 293147 -786 293175
rect -758 293147 -724 293175
rect -696 293147 -648 293175
rect -958 293113 -648 293147
rect -958 293085 -910 293113
rect -882 293085 -848 293113
rect -820 293085 -786 293113
rect -758 293085 -724 293113
rect -696 293085 -648 293113
rect -958 293051 -648 293085
rect -958 293023 -910 293051
rect -882 293023 -848 293051
rect -820 293023 -786 293051
rect -758 293023 -724 293051
rect -696 293023 -648 293051
rect -958 292989 -648 293023
rect -958 292961 -910 292989
rect -882 292961 -848 292989
rect -820 292961 -786 292989
rect -758 292961 -724 292989
rect -696 292961 -648 292989
rect -958 284175 -648 292961
rect -958 284147 -910 284175
rect -882 284147 -848 284175
rect -820 284147 -786 284175
rect -758 284147 -724 284175
rect -696 284147 -648 284175
rect -958 284113 -648 284147
rect -958 284085 -910 284113
rect -882 284085 -848 284113
rect -820 284085 -786 284113
rect -758 284085 -724 284113
rect -696 284085 -648 284113
rect -958 284051 -648 284085
rect -958 284023 -910 284051
rect -882 284023 -848 284051
rect -820 284023 -786 284051
rect -758 284023 -724 284051
rect -696 284023 -648 284051
rect -958 283989 -648 284023
rect -958 283961 -910 283989
rect -882 283961 -848 283989
rect -820 283961 -786 283989
rect -758 283961 -724 283989
rect -696 283961 -648 283989
rect -958 275175 -648 283961
rect -958 275147 -910 275175
rect -882 275147 -848 275175
rect -820 275147 -786 275175
rect -758 275147 -724 275175
rect -696 275147 -648 275175
rect -958 275113 -648 275147
rect -958 275085 -910 275113
rect -882 275085 -848 275113
rect -820 275085 -786 275113
rect -758 275085 -724 275113
rect -696 275085 -648 275113
rect -958 275051 -648 275085
rect -958 275023 -910 275051
rect -882 275023 -848 275051
rect -820 275023 -786 275051
rect -758 275023 -724 275051
rect -696 275023 -648 275051
rect -958 274989 -648 275023
rect -958 274961 -910 274989
rect -882 274961 -848 274989
rect -820 274961 -786 274989
rect -758 274961 -724 274989
rect -696 274961 -648 274989
rect -958 266175 -648 274961
rect -958 266147 -910 266175
rect -882 266147 -848 266175
rect -820 266147 -786 266175
rect -758 266147 -724 266175
rect -696 266147 -648 266175
rect -958 266113 -648 266147
rect -958 266085 -910 266113
rect -882 266085 -848 266113
rect -820 266085 -786 266113
rect -758 266085 -724 266113
rect -696 266085 -648 266113
rect -958 266051 -648 266085
rect -958 266023 -910 266051
rect -882 266023 -848 266051
rect -820 266023 -786 266051
rect -758 266023 -724 266051
rect -696 266023 -648 266051
rect -958 265989 -648 266023
rect -958 265961 -910 265989
rect -882 265961 -848 265989
rect -820 265961 -786 265989
rect -758 265961 -724 265989
rect -696 265961 -648 265989
rect -958 257175 -648 265961
rect -958 257147 -910 257175
rect -882 257147 -848 257175
rect -820 257147 -786 257175
rect -758 257147 -724 257175
rect -696 257147 -648 257175
rect -958 257113 -648 257147
rect -958 257085 -910 257113
rect -882 257085 -848 257113
rect -820 257085 -786 257113
rect -758 257085 -724 257113
rect -696 257085 -648 257113
rect -958 257051 -648 257085
rect -958 257023 -910 257051
rect -882 257023 -848 257051
rect -820 257023 -786 257051
rect -758 257023 -724 257051
rect -696 257023 -648 257051
rect -958 256989 -648 257023
rect -958 256961 -910 256989
rect -882 256961 -848 256989
rect -820 256961 -786 256989
rect -758 256961 -724 256989
rect -696 256961 -648 256989
rect -958 248175 -648 256961
rect -958 248147 -910 248175
rect -882 248147 -848 248175
rect -820 248147 -786 248175
rect -758 248147 -724 248175
rect -696 248147 -648 248175
rect -958 248113 -648 248147
rect -958 248085 -910 248113
rect -882 248085 -848 248113
rect -820 248085 -786 248113
rect -758 248085 -724 248113
rect -696 248085 -648 248113
rect -958 248051 -648 248085
rect -958 248023 -910 248051
rect -882 248023 -848 248051
rect -820 248023 -786 248051
rect -758 248023 -724 248051
rect -696 248023 -648 248051
rect -958 247989 -648 248023
rect -958 247961 -910 247989
rect -882 247961 -848 247989
rect -820 247961 -786 247989
rect -758 247961 -724 247989
rect -696 247961 -648 247989
rect -958 239175 -648 247961
rect -958 239147 -910 239175
rect -882 239147 -848 239175
rect -820 239147 -786 239175
rect -758 239147 -724 239175
rect -696 239147 -648 239175
rect -958 239113 -648 239147
rect -958 239085 -910 239113
rect -882 239085 -848 239113
rect -820 239085 -786 239113
rect -758 239085 -724 239113
rect -696 239085 -648 239113
rect -958 239051 -648 239085
rect -958 239023 -910 239051
rect -882 239023 -848 239051
rect -820 239023 -786 239051
rect -758 239023 -724 239051
rect -696 239023 -648 239051
rect -958 238989 -648 239023
rect -958 238961 -910 238989
rect -882 238961 -848 238989
rect -820 238961 -786 238989
rect -758 238961 -724 238989
rect -696 238961 -648 238989
rect -958 230175 -648 238961
rect -958 230147 -910 230175
rect -882 230147 -848 230175
rect -820 230147 -786 230175
rect -758 230147 -724 230175
rect -696 230147 -648 230175
rect -958 230113 -648 230147
rect -958 230085 -910 230113
rect -882 230085 -848 230113
rect -820 230085 -786 230113
rect -758 230085 -724 230113
rect -696 230085 -648 230113
rect -958 230051 -648 230085
rect -958 230023 -910 230051
rect -882 230023 -848 230051
rect -820 230023 -786 230051
rect -758 230023 -724 230051
rect -696 230023 -648 230051
rect -958 229989 -648 230023
rect -958 229961 -910 229989
rect -882 229961 -848 229989
rect -820 229961 -786 229989
rect -758 229961 -724 229989
rect -696 229961 -648 229989
rect -958 221175 -648 229961
rect -958 221147 -910 221175
rect -882 221147 -848 221175
rect -820 221147 -786 221175
rect -758 221147 -724 221175
rect -696 221147 -648 221175
rect -958 221113 -648 221147
rect -958 221085 -910 221113
rect -882 221085 -848 221113
rect -820 221085 -786 221113
rect -758 221085 -724 221113
rect -696 221085 -648 221113
rect -958 221051 -648 221085
rect -958 221023 -910 221051
rect -882 221023 -848 221051
rect -820 221023 -786 221051
rect -758 221023 -724 221051
rect -696 221023 -648 221051
rect -958 220989 -648 221023
rect -958 220961 -910 220989
rect -882 220961 -848 220989
rect -820 220961 -786 220989
rect -758 220961 -724 220989
rect -696 220961 -648 220989
rect -958 212175 -648 220961
rect -958 212147 -910 212175
rect -882 212147 -848 212175
rect -820 212147 -786 212175
rect -758 212147 -724 212175
rect -696 212147 -648 212175
rect -958 212113 -648 212147
rect -958 212085 -910 212113
rect -882 212085 -848 212113
rect -820 212085 -786 212113
rect -758 212085 -724 212113
rect -696 212085 -648 212113
rect -958 212051 -648 212085
rect -958 212023 -910 212051
rect -882 212023 -848 212051
rect -820 212023 -786 212051
rect -758 212023 -724 212051
rect -696 212023 -648 212051
rect -958 211989 -648 212023
rect -958 211961 -910 211989
rect -882 211961 -848 211989
rect -820 211961 -786 211989
rect -758 211961 -724 211989
rect -696 211961 -648 211989
rect -958 203175 -648 211961
rect -958 203147 -910 203175
rect -882 203147 -848 203175
rect -820 203147 -786 203175
rect -758 203147 -724 203175
rect -696 203147 -648 203175
rect -958 203113 -648 203147
rect -958 203085 -910 203113
rect -882 203085 -848 203113
rect -820 203085 -786 203113
rect -758 203085 -724 203113
rect -696 203085 -648 203113
rect -958 203051 -648 203085
rect -958 203023 -910 203051
rect -882 203023 -848 203051
rect -820 203023 -786 203051
rect -758 203023 -724 203051
rect -696 203023 -648 203051
rect -958 202989 -648 203023
rect -958 202961 -910 202989
rect -882 202961 -848 202989
rect -820 202961 -786 202989
rect -758 202961 -724 202989
rect -696 202961 -648 202989
rect -958 194175 -648 202961
rect -958 194147 -910 194175
rect -882 194147 -848 194175
rect -820 194147 -786 194175
rect -758 194147 -724 194175
rect -696 194147 -648 194175
rect -958 194113 -648 194147
rect -958 194085 -910 194113
rect -882 194085 -848 194113
rect -820 194085 -786 194113
rect -758 194085 -724 194113
rect -696 194085 -648 194113
rect -958 194051 -648 194085
rect -958 194023 -910 194051
rect -882 194023 -848 194051
rect -820 194023 -786 194051
rect -758 194023 -724 194051
rect -696 194023 -648 194051
rect -958 193989 -648 194023
rect -958 193961 -910 193989
rect -882 193961 -848 193989
rect -820 193961 -786 193989
rect -758 193961 -724 193989
rect -696 193961 -648 193989
rect -958 185175 -648 193961
rect -958 185147 -910 185175
rect -882 185147 -848 185175
rect -820 185147 -786 185175
rect -758 185147 -724 185175
rect -696 185147 -648 185175
rect -958 185113 -648 185147
rect -958 185085 -910 185113
rect -882 185085 -848 185113
rect -820 185085 -786 185113
rect -758 185085 -724 185113
rect -696 185085 -648 185113
rect -958 185051 -648 185085
rect -958 185023 -910 185051
rect -882 185023 -848 185051
rect -820 185023 -786 185051
rect -758 185023 -724 185051
rect -696 185023 -648 185051
rect -958 184989 -648 185023
rect -958 184961 -910 184989
rect -882 184961 -848 184989
rect -820 184961 -786 184989
rect -758 184961 -724 184989
rect -696 184961 -648 184989
rect -958 176175 -648 184961
rect -958 176147 -910 176175
rect -882 176147 -848 176175
rect -820 176147 -786 176175
rect -758 176147 -724 176175
rect -696 176147 -648 176175
rect -958 176113 -648 176147
rect -958 176085 -910 176113
rect -882 176085 -848 176113
rect -820 176085 -786 176113
rect -758 176085 -724 176113
rect -696 176085 -648 176113
rect -958 176051 -648 176085
rect -958 176023 -910 176051
rect -882 176023 -848 176051
rect -820 176023 -786 176051
rect -758 176023 -724 176051
rect -696 176023 -648 176051
rect -958 175989 -648 176023
rect -958 175961 -910 175989
rect -882 175961 -848 175989
rect -820 175961 -786 175989
rect -758 175961 -724 175989
rect -696 175961 -648 175989
rect -958 167175 -648 175961
rect -958 167147 -910 167175
rect -882 167147 -848 167175
rect -820 167147 -786 167175
rect -758 167147 -724 167175
rect -696 167147 -648 167175
rect -958 167113 -648 167147
rect -958 167085 -910 167113
rect -882 167085 -848 167113
rect -820 167085 -786 167113
rect -758 167085 -724 167113
rect -696 167085 -648 167113
rect -958 167051 -648 167085
rect -958 167023 -910 167051
rect -882 167023 -848 167051
rect -820 167023 -786 167051
rect -758 167023 -724 167051
rect -696 167023 -648 167051
rect -958 166989 -648 167023
rect -958 166961 -910 166989
rect -882 166961 -848 166989
rect -820 166961 -786 166989
rect -758 166961 -724 166989
rect -696 166961 -648 166989
rect -958 158175 -648 166961
rect -958 158147 -910 158175
rect -882 158147 -848 158175
rect -820 158147 -786 158175
rect -758 158147 -724 158175
rect -696 158147 -648 158175
rect -958 158113 -648 158147
rect -958 158085 -910 158113
rect -882 158085 -848 158113
rect -820 158085 -786 158113
rect -758 158085 -724 158113
rect -696 158085 -648 158113
rect -958 158051 -648 158085
rect -958 158023 -910 158051
rect -882 158023 -848 158051
rect -820 158023 -786 158051
rect -758 158023 -724 158051
rect -696 158023 -648 158051
rect -958 157989 -648 158023
rect -958 157961 -910 157989
rect -882 157961 -848 157989
rect -820 157961 -786 157989
rect -758 157961 -724 157989
rect -696 157961 -648 157989
rect -958 149175 -648 157961
rect -958 149147 -910 149175
rect -882 149147 -848 149175
rect -820 149147 -786 149175
rect -758 149147 -724 149175
rect -696 149147 -648 149175
rect -958 149113 -648 149147
rect -958 149085 -910 149113
rect -882 149085 -848 149113
rect -820 149085 -786 149113
rect -758 149085 -724 149113
rect -696 149085 -648 149113
rect -958 149051 -648 149085
rect -958 149023 -910 149051
rect -882 149023 -848 149051
rect -820 149023 -786 149051
rect -758 149023 -724 149051
rect -696 149023 -648 149051
rect -958 148989 -648 149023
rect -958 148961 -910 148989
rect -882 148961 -848 148989
rect -820 148961 -786 148989
rect -758 148961 -724 148989
rect -696 148961 -648 148989
rect -958 140175 -648 148961
rect -958 140147 -910 140175
rect -882 140147 -848 140175
rect -820 140147 -786 140175
rect -758 140147 -724 140175
rect -696 140147 -648 140175
rect -958 140113 -648 140147
rect -958 140085 -910 140113
rect -882 140085 -848 140113
rect -820 140085 -786 140113
rect -758 140085 -724 140113
rect -696 140085 -648 140113
rect -958 140051 -648 140085
rect -958 140023 -910 140051
rect -882 140023 -848 140051
rect -820 140023 -786 140051
rect -758 140023 -724 140051
rect -696 140023 -648 140051
rect -958 139989 -648 140023
rect -958 139961 -910 139989
rect -882 139961 -848 139989
rect -820 139961 -786 139989
rect -758 139961 -724 139989
rect -696 139961 -648 139989
rect -958 131175 -648 139961
rect -958 131147 -910 131175
rect -882 131147 -848 131175
rect -820 131147 -786 131175
rect -758 131147 -724 131175
rect -696 131147 -648 131175
rect -958 131113 -648 131147
rect -958 131085 -910 131113
rect -882 131085 -848 131113
rect -820 131085 -786 131113
rect -758 131085 -724 131113
rect -696 131085 -648 131113
rect -958 131051 -648 131085
rect -958 131023 -910 131051
rect -882 131023 -848 131051
rect -820 131023 -786 131051
rect -758 131023 -724 131051
rect -696 131023 -648 131051
rect -958 130989 -648 131023
rect -958 130961 -910 130989
rect -882 130961 -848 130989
rect -820 130961 -786 130989
rect -758 130961 -724 130989
rect -696 130961 -648 130989
rect -958 122175 -648 130961
rect -958 122147 -910 122175
rect -882 122147 -848 122175
rect -820 122147 -786 122175
rect -758 122147 -724 122175
rect -696 122147 -648 122175
rect -958 122113 -648 122147
rect -958 122085 -910 122113
rect -882 122085 -848 122113
rect -820 122085 -786 122113
rect -758 122085 -724 122113
rect -696 122085 -648 122113
rect -958 122051 -648 122085
rect -958 122023 -910 122051
rect -882 122023 -848 122051
rect -820 122023 -786 122051
rect -758 122023 -724 122051
rect -696 122023 -648 122051
rect -958 121989 -648 122023
rect -958 121961 -910 121989
rect -882 121961 -848 121989
rect -820 121961 -786 121989
rect -758 121961 -724 121989
rect -696 121961 -648 121989
rect -958 113175 -648 121961
rect -958 113147 -910 113175
rect -882 113147 -848 113175
rect -820 113147 -786 113175
rect -758 113147 -724 113175
rect -696 113147 -648 113175
rect -958 113113 -648 113147
rect -958 113085 -910 113113
rect -882 113085 -848 113113
rect -820 113085 -786 113113
rect -758 113085 -724 113113
rect -696 113085 -648 113113
rect -958 113051 -648 113085
rect -958 113023 -910 113051
rect -882 113023 -848 113051
rect -820 113023 -786 113051
rect -758 113023 -724 113051
rect -696 113023 -648 113051
rect -958 112989 -648 113023
rect -958 112961 -910 112989
rect -882 112961 -848 112989
rect -820 112961 -786 112989
rect -758 112961 -724 112989
rect -696 112961 -648 112989
rect -958 104175 -648 112961
rect -958 104147 -910 104175
rect -882 104147 -848 104175
rect -820 104147 -786 104175
rect -758 104147 -724 104175
rect -696 104147 -648 104175
rect -958 104113 -648 104147
rect -958 104085 -910 104113
rect -882 104085 -848 104113
rect -820 104085 -786 104113
rect -758 104085 -724 104113
rect -696 104085 -648 104113
rect -958 104051 -648 104085
rect -958 104023 -910 104051
rect -882 104023 -848 104051
rect -820 104023 -786 104051
rect -758 104023 -724 104051
rect -696 104023 -648 104051
rect -958 103989 -648 104023
rect -958 103961 -910 103989
rect -882 103961 -848 103989
rect -820 103961 -786 103989
rect -758 103961 -724 103989
rect -696 103961 -648 103989
rect -958 95175 -648 103961
rect -958 95147 -910 95175
rect -882 95147 -848 95175
rect -820 95147 -786 95175
rect -758 95147 -724 95175
rect -696 95147 -648 95175
rect -958 95113 -648 95147
rect -958 95085 -910 95113
rect -882 95085 -848 95113
rect -820 95085 -786 95113
rect -758 95085 -724 95113
rect -696 95085 -648 95113
rect -958 95051 -648 95085
rect -958 95023 -910 95051
rect -882 95023 -848 95051
rect -820 95023 -786 95051
rect -758 95023 -724 95051
rect -696 95023 -648 95051
rect -958 94989 -648 95023
rect -958 94961 -910 94989
rect -882 94961 -848 94989
rect -820 94961 -786 94989
rect -758 94961 -724 94989
rect -696 94961 -648 94989
rect -958 86175 -648 94961
rect -958 86147 -910 86175
rect -882 86147 -848 86175
rect -820 86147 -786 86175
rect -758 86147 -724 86175
rect -696 86147 -648 86175
rect -958 86113 -648 86147
rect -958 86085 -910 86113
rect -882 86085 -848 86113
rect -820 86085 -786 86113
rect -758 86085 -724 86113
rect -696 86085 -648 86113
rect -958 86051 -648 86085
rect -958 86023 -910 86051
rect -882 86023 -848 86051
rect -820 86023 -786 86051
rect -758 86023 -724 86051
rect -696 86023 -648 86051
rect -958 85989 -648 86023
rect -958 85961 -910 85989
rect -882 85961 -848 85989
rect -820 85961 -786 85989
rect -758 85961 -724 85989
rect -696 85961 -648 85989
rect -958 77175 -648 85961
rect -958 77147 -910 77175
rect -882 77147 -848 77175
rect -820 77147 -786 77175
rect -758 77147 -724 77175
rect -696 77147 -648 77175
rect -958 77113 -648 77147
rect -958 77085 -910 77113
rect -882 77085 -848 77113
rect -820 77085 -786 77113
rect -758 77085 -724 77113
rect -696 77085 -648 77113
rect -958 77051 -648 77085
rect -958 77023 -910 77051
rect -882 77023 -848 77051
rect -820 77023 -786 77051
rect -758 77023 -724 77051
rect -696 77023 -648 77051
rect -958 76989 -648 77023
rect -958 76961 -910 76989
rect -882 76961 -848 76989
rect -820 76961 -786 76989
rect -758 76961 -724 76989
rect -696 76961 -648 76989
rect -958 68175 -648 76961
rect -958 68147 -910 68175
rect -882 68147 -848 68175
rect -820 68147 -786 68175
rect -758 68147 -724 68175
rect -696 68147 -648 68175
rect -958 68113 -648 68147
rect -958 68085 -910 68113
rect -882 68085 -848 68113
rect -820 68085 -786 68113
rect -758 68085 -724 68113
rect -696 68085 -648 68113
rect -958 68051 -648 68085
rect -958 68023 -910 68051
rect -882 68023 -848 68051
rect -820 68023 -786 68051
rect -758 68023 -724 68051
rect -696 68023 -648 68051
rect -958 67989 -648 68023
rect -958 67961 -910 67989
rect -882 67961 -848 67989
rect -820 67961 -786 67989
rect -758 67961 -724 67989
rect -696 67961 -648 67989
rect -958 59175 -648 67961
rect -958 59147 -910 59175
rect -882 59147 -848 59175
rect -820 59147 -786 59175
rect -758 59147 -724 59175
rect -696 59147 -648 59175
rect -958 59113 -648 59147
rect -958 59085 -910 59113
rect -882 59085 -848 59113
rect -820 59085 -786 59113
rect -758 59085 -724 59113
rect -696 59085 -648 59113
rect -958 59051 -648 59085
rect -958 59023 -910 59051
rect -882 59023 -848 59051
rect -820 59023 -786 59051
rect -758 59023 -724 59051
rect -696 59023 -648 59051
rect -958 58989 -648 59023
rect -958 58961 -910 58989
rect -882 58961 -848 58989
rect -820 58961 -786 58989
rect -758 58961 -724 58989
rect -696 58961 -648 58989
rect -958 50175 -648 58961
rect -958 50147 -910 50175
rect -882 50147 -848 50175
rect -820 50147 -786 50175
rect -758 50147 -724 50175
rect -696 50147 -648 50175
rect -958 50113 -648 50147
rect -958 50085 -910 50113
rect -882 50085 -848 50113
rect -820 50085 -786 50113
rect -758 50085 -724 50113
rect -696 50085 -648 50113
rect -958 50051 -648 50085
rect -958 50023 -910 50051
rect -882 50023 -848 50051
rect -820 50023 -786 50051
rect -758 50023 -724 50051
rect -696 50023 -648 50051
rect -958 49989 -648 50023
rect -958 49961 -910 49989
rect -882 49961 -848 49989
rect -820 49961 -786 49989
rect -758 49961 -724 49989
rect -696 49961 -648 49989
rect -958 41175 -648 49961
rect -958 41147 -910 41175
rect -882 41147 -848 41175
rect -820 41147 -786 41175
rect -758 41147 -724 41175
rect -696 41147 -648 41175
rect -958 41113 -648 41147
rect -958 41085 -910 41113
rect -882 41085 -848 41113
rect -820 41085 -786 41113
rect -758 41085 -724 41113
rect -696 41085 -648 41113
rect -958 41051 -648 41085
rect -958 41023 -910 41051
rect -882 41023 -848 41051
rect -820 41023 -786 41051
rect -758 41023 -724 41051
rect -696 41023 -648 41051
rect -958 40989 -648 41023
rect -958 40961 -910 40989
rect -882 40961 -848 40989
rect -820 40961 -786 40989
rect -758 40961 -724 40989
rect -696 40961 -648 40989
rect -958 32175 -648 40961
rect -958 32147 -910 32175
rect -882 32147 -848 32175
rect -820 32147 -786 32175
rect -758 32147 -724 32175
rect -696 32147 -648 32175
rect -958 32113 -648 32147
rect -958 32085 -910 32113
rect -882 32085 -848 32113
rect -820 32085 -786 32113
rect -758 32085 -724 32113
rect -696 32085 -648 32113
rect -958 32051 -648 32085
rect -958 32023 -910 32051
rect -882 32023 -848 32051
rect -820 32023 -786 32051
rect -758 32023 -724 32051
rect -696 32023 -648 32051
rect -958 31989 -648 32023
rect -958 31961 -910 31989
rect -882 31961 -848 31989
rect -820 31961 -786 31989
rect -758 31961 -724 31989
rect -696 31961 -648 31989
rect -958 23175 -648 31961
rect -958 23147 -910 23175
rect -882 23147 -848 23175
rect -820 23147 -786 23175
rect -758 23147 -724 23175
rect -696 23147 -648 23175
rect -958 23113 -648 23147
rect -958 23085 -910 23113
rect -882 23085 -848 23113
rect -820 23085 -786 23113
rect -758 23085 -724 23113
rect -696 23085 -648 23113
rect -958 23051 -648 23085
rect -958 23023 -910 23051
rect -882 23023 -848 23051
rect -820 23023 -786 23051
rect -758 23023 -724 23051
rect -696 23023 -648 23051
rect -958 22989 -648 23023
rect -958 22961 -910 22989
rect -882 22961 -848 22989
rect -820 22961 -786 22989
rect -758 22961 -724 22989
rect -696 22961 -648 22989
rect -958 14175 -648 22961
rect -958 14147 -910 14175
rect -882 14147 -848 14175
rect -820 14147 -786 14175
rect -758 14147 -724 14175
rect -696 14147 -648 14175
rect -958 14113 -648 14147
rect -958 14085 -910 14113
rect -882 14085 -848 14113
rect -820 14085 -786 14113
rect -758 14085 -724 14113
rect -696 14085 -648 14113
rect -958 14051 -648 14085
rect -958 14023 -910 14051
rect -882 14023 -848 14051
rect -820 14023 -786 14051
rect -758 14023 -724 14051
rect -696 14023 -648 14051
rect -958 13989 -648 14023
rect -958 13961 -910 13989
rect -882 13961 -848 13989
rect -820 13961 -786 13989
rect -758 13961 -724 13989
rect -696 13961 -648 13989
rect -958 5175 -648 13961
rect -958 5147 -910 5175
rect -882 5147 -848 5175
rect -820 5147 -786 5175
rect -758 5147 -724 5175
rect -696 5147 -648 5175
rect -958 5113 -648 5147
rect -958 5085 -910 5113
rect -882 5085 -848 5113
rect -820 5085 -786 5113
rect -758 5085 -724 5113
rect -696 5085 -648 5113
rect -958 5051 -648 5085
rect -958 5023 -910 5051
rect -882 5023 -848 5051
rect -820 5023 -786 5051
rect -758 5023 -724 5051
rect -696 5023 -648 5051
rect -958 4989 -648 5023
rect -958 4961 -910 4989
rect -882 4961 -848 4989
rect -820 4961 -786 4989
rect -758 4961 -724 4989
rect -696 4961 -648 4989
rect -958 -560 -648 4961
rect -478 298606 -168 298654
rect -478 298578 -430 298606
rect -402 298578 -368 298606
rect -340 298578 -306 298606
rect -278 298578 -244 298606
rect -216 298578 -168 298606
rect -478 298544 -168 298578
rect -478 298516 -430 298544
rect -402 298516 -368 298544
rect -340 298516 -306 298544
rect -278 298516 -244 298544
rect -216 298516 -168 298544
rect -478 298482 -168 298516
rect -478 298454 -430 298482
rect -402 298454 -368 298482
rect -340 298454 -306 298482
rect -278 298454 -244 298482
rect -216 298454 -168 298482
rect -478 298420 -168 298454
rect -478 298392 -430 298420
rect -402 298392 -368 298420
rect -340 298392 -306 298420
rect -278 298392 -244 298420
rect -216 298392 -168 298420
rect -478 290175 -168 298392
rect -478 290147 -430 290175
rect -402 290147 -368 290175
rect -340 290147 -306 290175
rect -278 290147 -244 290175
rect -216 290147 -168 290175
rect -478 290113 -168 290147
rect -478 290085 -430 290113
rect -402 290085 -368 290113
rect -340 290085 -306 290113
rect -278 290085 -244 290113
rect -216 290085 -168 290113
rect -478 290051 -168 290085
rect -478 290023 -430 290051
rect -402 290023 -368 290051
rect -340 290023 -306 290051
rect -278 290023 -244 290051
rect -216 290023 -168 290051
rect -478 289989 -168 290023
rect -478 289961 -430 289989
rect -402 289961 -368 289989
rect -340 289961 -306 289989
rect -278 289961 -244 289989
rect -216 289961 -168 289989
rect -478 281175 -168 289961
rect -478 281147 -430 281175
rect -402 281147 -368 281175
rect -340 281147 -306 281175
rect -278 281147 -244 281175
rect -216 281147 -168 281175
rect -478 281113 -168 281147
rect -478 281085 -430 281113
rect -402 281085 -368 281113
rect -340 281085 -306 281113
rect -278 281085 -244 281113
rect -216 281085 -168 281113
rect -478 281051 -168 281085
rect -478 281023 -430 281051
rect -402 281023 -368 281051
rect -340 281023 -306 281051
rect -278 281023 -244 281051
rect -216 281023 -168 281051
rect -478 280989 -168 281023
rect -478 280961 -430 280989
rect -402 280961 -368 280989
rect -340 280961 -306 280989
rect -278 280961 -244 280989
rect -216 280961 -168 280989
rect -478 272175 -168 280961
rect -478 272147 -430 272175
rect -402 272147 -368 272175
rect -340 272147 -306 272175
rect -278 272147 -244 272175
rect -216 272147 -168 272175
rect -478 272113 -168 272147
rect -478 272085 -430 272113
rect -402 272085 -368 272113
rect -340 272085 -306 272113
rect -278 272085 -244 272113
rect -216 272085 -168 272113
rect -478 272051 -168 272085
rect -478 272023 -430 272051
rect -402 272023 -368 272051
rect -340 272023 -306 272051
rect -278 272023 -244 272051
rect -216 272023 -168 272051
rect -478 271989 -168 272023
rect -478 271961 -430 271989
rect -402 271961 -368 271989
rect -340 271961 -306 271989
rect -278 271961 -244 271989
rect -216 271961 -168 271989
rect -478 263175 -168 271961
rect -478 263147 -430 263175
rect -402 263147 -368 263175
rect -340 263147 -306 263175
rect -278 263147 -244 263175
rect -216 263147 -168 263175
rect -478 263113 -168 263147
rect -478 263085 -430 263113
rect -402 263085 -368 263113
rect -340 263085 -306 263113
rect -278 263085 -244 263113
rect -216 263085 -168 263113
rect -478 263051 -168 263085
rect -478 263023 -430 263051
rect -402 263023 -368 263051
rect -340 263023 -306 263051
rect -278 263023 -244 263051
rect -216 263023 -168 263051
rect -478 262989 -168 263023
rect -478 262961 -430 262989
rect -402 262961 -368 262989
rect -340 262961 -306 262989
rect -278 262961 -244 262989
rect -216 262961 -168 262989
rect -478 254175 -168 262961
rect -478 254147 -430 254175
rect -402 254147 -368 254175
rect -340 254147 -306 254175
rect -278 254147 -244 254175
rect -216 254147 -168 254175
rect -478 254113 -168 254147
rect -478 254085 -430 254113
rect -402 254085 -368 254113
rect -340 254085 -306 254113
rect -278 254085 -244 254113
rect -216 254085 -168 254113
rect -478 254051 -168 254085
rect -478 254023 -430 254051
rect -402 254023 -368 254051
rect -340 254023 -306 254051
rect -278 254023 -244 254051
rect -216 254023 -168 254051
rect -478 253989 -168 254023
rect -478 253961 -430 253989
rect -402 253961 -368 253989
rect -340 253961 -306 253989
rect -278 253961 -244 253989
rect -216 253961 -168 253989
rect -478 245175 -168 253961
rect -478 245147 -430 245175
rect -402 245147 -368 245175
rect -340 245147 -306 245175
rect -278 245147 -244 245175
rect -216 245147 -168 245175
rect -478 245113 -168 245147
rect -478 245085 -430 245113
rect -402 245085 -368 245113
rect -340 245085 -306 245113
rect -278 245085 -244 245113
rect -216 245085 -168 245113
rect -478 245051 -168 245085
rect -478 245023 -430 245051
rect -402 245023 -368 245051
rect -340 245023 -306 245051
rect -278 245023 -244 245051
rect -216 245023 -168 245051
rect -478 244989 -168 245023
rect -478 244961 -430 244989
rect -402 244961 -368 244989
rect -340 244961 -306 244989
rect -278 244961 -244 244989
rect -216 244961 -168 244989
rect -478 236175 -168 244961
rect -478 236147 -430 236175
rect -402 236147 -368 236175
rect -340 236147 -306 236175
rect -278 236147 -244 236175
rect -216 236147 -168 236175
rect -478 236113 -168 236147
rect -478 236085 -430 236113
rect -402 236085 -368 236113
rect -340 236085 -306 236113
rect -278 236085 -244 236113
rect -216 236085 -168 236113
rect -478 236051 -168 236085
rect -478 236023 -430 236051
rect -402 236023 -368 236051
rect -340 236023 -306 236051
rect -278 236023 -244 236051
rect -216 236023 -168 236051
rect -478 235989 -168 236023
rect -478 235961 -430 235989
rect -402 235961 -368 235989
rect -340 235961 -306 235989
rect -278 235961 -244 235989
rect -216 235961 -168 235989
rect -478 227175 -168 235961
rect -478 227147 -430 227175
rect -402 227147 -368 227175
rect -340 227147 -306 227175
rect -278 227147 -244 227175
rect -216 227147 -168 227175
rect -478 227113 -168 227147
rect -478 227085 -430 227113
rect -402 227085 -368 227113
rect -340 227085 -306 227113
rect -278 227085 -244 227113
rect -216 227085 -168 227113
rect -478 227051 -168 227085
rect -478 227023 -430 227051
rect -402 227023 -368 227051
rect -340 227023 -306 227051
rect -278 227023 -244 227051
rect -216 227023 -168 227051
rect -478 226989 -168 227023
rect -478 226961 -430 226989
rect -402 226961 -368 226989
rect -340 226961 -306 226989
rect -278 226961 -244 226989
rect -216 226961 -168 226989
rect -478 218175 -168 226961
rect -478 218147 -430 218175
rect -402 218147 -368 218175
rect -340 218147 -306 218175
rect -278 218147 -244 218175
rect -216 218147 -168 218175
rect -478 218113 -168 218147
rect -478 218085 -430 218113
rect -402 218085 -368 218113
rect -340 218085 -306 218113
rect -278 218085 -244 218113
rect -216 218085 -168 218113
rect -478 218051 -168 218085
rect -478 218023 -430 218051
rect -402 218023 -368 218051
rect -340 218023 -306 218051
rect -278 218023 -244 218051
rect -216 218023 -168 218051
rect -478 217989 -168 218023
rect -478 217961 -430 217989
rect -402 217961 -368 217989
rect -340 217961 -306 217989
rect -278 217961 -244 217989
rect -216 217961 -168 217989
rect -478 209175 -168 217961
rect -478 209147 -430 209175
rect -402 209147 -368 209175
rect -340 209147 -306 209175
rect -278 209147 -244 209175
rect -216 209147 -168 209175
rect -478 209113 -168 209147
rect -478 209085 -430 209113
rect -402 209085 -368 209113
rect -340 209085 -306 209113
rect -278 209085 -244 209113
rect -216 209085 -168 209113
rect -478 209051 -168 209085
rect -478 209023 -430 209051
rect -402 209023 -368 209051
rect -340 209023 -306 209051
rect -278 209023 -244 209051
rect -216 209023 -168 209051
rect -478 208989 -168 209023
rect -478 208961 -430 208989
rect -402 208961 -368 208989
rect -340 208961 -306 208989
rect -278 208961 -244 208989
rect -216 208961 -168 208989
rect -478 200175 -168 208961
rect -478 200147 -430 200175
rect -402 200147 -368 200175
rect -340 200147 -306 200175
rect -278 200147 -244 200175
rect -216 200147 -168 200175
rect -478 200113 -168 200147
rect -478 200085 -430 200113
rect -402 200085 -368 200113
rect -340 200085 -306 200113
rect -278 200085 -244 200113
rect -216 200085 -168 200113
rect -478 200051 -168 200085
rect -478 200023 -430 200051
rect -402 200023 -368 200051
rect -340 200023 -306 200051
rect -278 200023 -244 200051
rect -216 200023 -168 200051
rect -478 199989 -168 200023
rect -478 199961 -430 199989
rect -402 199961 -368 199989
rect -340 199961 -306 199989
rect -278 199961 -244 199989
rect -216 199961 -168 199989
rect -478 191175 -168 199961
rect -478 191147 -430 191175
rect -402 191147 -368 191175
rect -340 191147 -306 191175
rect -278 191147 -244 191175
rect -216 191147 -168 191175
rect -478 191113 -168 191147
rect -478 191085 -430 191113
rect -402 191085 -368 191113
rect -340 191085 -306 191113
rect -278 191085 -244 191113
rect -216 191085 -168 191113
rect -478 191051 -168 191085
rect -478 191023 -430 191051
rect -402 191023 -368 191051
rect -340 191023 -306 191051
rect -278 191023 -244 191051
rect -216 191023 -168 191051
rect -478 190989 -168 191023
rect -478 190961 -430 190989
rect -402 190961 -368 190989
rect -340 190961 -306 190989
rect -278 190961 -244 190989
rect -216 190961 -168 190989
rect -478 182175 -168 190961
rect -478 182147 -430 182175
rect -402 182147 -368 182175
rect -340 182147 -306 182175
rect -278 182147 -244 182175
rect -216 182147 -168 182175
rect -478 182113 -168 182147
rect -478 182085 -430 182113
rect -402 182085 -368 182113
rect -340 182085 -306 182113
rect -278 182085 -244 182113
rect -216 182085 -168 182113
rect -478 182051 -168 182085
rect -478 182023 -430 182051
rect -402 182023 -368 182051
rect -340 182023 -306 182051
rect -278 182023 -244 182051
rect -216 182023 -168 182051
rect -478 181989 -168 182023
rect -478 181961 -430 181989
rect -402 181961 -368 181989
rect -340 181961 -306 181989
rect -278 181961 -244 181989
rect -216 181961 -168 181989
rect -478 173175 -168 181961
rect -478 173147 -430 173175
rect -402 173147 -368 173175
rect -340 173147 -306 173175
rect -278 173147 -244 173175
rect -216 173147 -168 173175
rect -478 173113 -168 173147
rect -478 173085 -430 173113
rect -402 173085 -368 173113
rect -340 173085 -306 173113
rect -278 173085 -244 173113
rect -216 173085 -168 173113
rect -478 173051 -168 173085
rect -478 173023 -430 173051
rect -402 173023 -368 173051
rect -340 173023 -306 173051
rect -278 173023 -244 173051
rect -216 173023 -168 173051
rect -478 172989 -168 173023
rect -478 172961 -430 172989
rect -402 172961 -368 172989
rect -340 172961 -306 172989
rect -278 172961 -244 172989
rect -216 172961 -168 172989
rect -478 164175 -168 172961
rect -478 164147 -430 164175
rect -402 164147 -368 164175
rect -340 164147 -306 164175
rect -278 164147 -244 164175
rect -216 164147 -168 164175
rect -478 164113 -168 164147
rect -478 164085 -430 164113
rect -402 164085 -368 164113
rect -340 164085 -306 164113
rect -278 164085 -244 164113
rect -216 164085 -168 164113
rect -478 164051 -168 164085
rect -478 164023 -430 164051
rect -402 164023 -368 164051
rect -340 164023 -306 164051
rect -278 164023 -244 164051
rect -216 164023 -168 164051
rect -478 163989 -168 164023
rect -478 163961 -430 163989
rect -402 163961 -368 163989
rect -340 163961 -306 163989
rect -278 163961 -244 163989
rect -216 163961 -168 163989
rect -478 155175 -168 163961
rect -478 155147 -430 155175
rect -402 155147 -368 155175
rect -340 155147 -306 155175
rect -278 155147 -244 155175
rect -216 155147 -168 155175
rect -478 155113 -168 155147
rect -478 155085 -430 155113
rect -402 155085 -368 155113
rect -340 155085 -306 155113
rect -278 155085 -244 155113
rect -216 155085 -168 155113
rect -478 155051 -168 155085
rect -478 155023 -430 155051
rect -402 155023 -368 155051
rect -340 155023 -306 155051
rect -278 155023 -244 155051
rect -216 155023 -168 155051
rect -478 154989 -168 155023
rect -478 154961 -430 154989
rect -402 154961 -368 154989
rect -340 154961 -306 154989
rect -278 154961 -244 154989
rect -216 154961 -168 154989
rect -478 146175 -168 154961
rect -478 146147 -430 146175
rect -402 146147 -368 146175
rect -340 146147 -306 146175
rect -278 146147 -244 146175
rect -216 146147 -168 146175
rect -478 146113 -168 146147
rect -478 146085 -430 146113
rect -402 146085 -368 146113
rect -340 146085 -306 146113
rect -278 146085 -244 146113
rect -216 146085 -168 146113
rect -478 146051 -168 146085
rect -478 146023 -430 146051
rect -402 146023 -368 146051
rect -340 146023 -306 146051
rect -278 146023 -244 146051
rect -216 146023 -168 146051
rect -478 145989 -168 146023
rect -478 145961 -430 145989
rect -402 145961 -368 145989
rect -340 145961 -306 145989
rect -278 145961 -244 145989
rect -216 145961 -168 145989
rect -478 137175 -168 145961
rect -478 137147 -430 137175
rect -402 137147 -368 137175
rect -340 137147 -306 137175
rect -278 137147 -244 137175
rect -216 137147 -168 137175
rect -478 137113 -168 137147
rect -478 137085 -430 137113
rect -402 137085 -368 137113
rect -340 137085 -306 137113
rect -278 137085 -244 137113
rect -216 137085 -168 137113
rect -478 137051 -168 137085
rect -478 137023 -430 137051
rect -402 137023 -368 137051
rect -340 137023 -306 137051
rect -278 137023 -244 137051
rect -216 137023 -168 137051
rect -478 136989 -168 137023
rect -478 136961 -430 136989
rect -402 136961 -368 136989
rect -340 136961 -306 136989
rect -278 136961 -244 136989
rect -216 136961 -168 136989
rect -478 128175 -168 136961
rect -478 128147 -430 128175
rect -402 128147 -368 128175
rect -340 128147 -306 128175
rect -278 128147 -244 128175
rect -216 128147 -168 128175
rect -478 128113 -168 128147
rect -478 128085 -430 128113
rect -402 128085 -368 128113
rect -340 128085 -306 128113
rect -278 128085 -244 128113
rect -216 128085 -168 128113
rect -478 128051 -168 128085
rect -478 128023 -430 128051
rect -402 128023 -368 128051
rect -340 128023 -306 128051
rect -278 128023 -244 128051
rect -216 128023 -168 128051
rect -478 127989 -168 128023
rect -478 127961 -430 127989
rect -402 127961 -368 127989
rect -340 127961 -306 127989
rect -278 127961 -244 127989
rect -216 127961 -168 127989
rect -478 119175 -168 127961
rect -478 119147 -430 119175
rect -402 119147 -368 119175
rect -340 119147 -306 119175
rect -278 119147 -244 119175
rect -216 119147 -168 119175
rect -478 119113 -168 119147
rect -478 119085 -430 119113
rect -402 119085 -368 119113
rect -340 119085 -306 119113
rect -278 119085 -244 119113
rect -216 119085 -168 119113
rect -478 119051 -168 119085
rect -478 119023 -430 119051
rect -402 119023 -368 119051
rect -340 119023 -306 119051
rect -278 119023 -244 119051
rect -216 119023 -168 119051
rect -478 118989 -168 119023
rect -478 118961 -430 118989
rect -402 118961 -368 118989
rect -340 118961 -306 118989
rect -278 118961 -244 118989
rect -216 118961 -168 118989
rect -478 110175 -168 118961
rect 2709 298606 3019 299134
rect 2709 298578 2757 298606
rect 2785 298578 2819 298606
rect 2847 298578 2881 298606
rect 2909 298578 2943 298606
rect 2971 298578 3019 298606
rect 2709 298544 3019 298578
rect 2709 298516 2757 298544
rect 2785 298516 2819 298544
rect 2847 298516 2881 298544
rect 2909 298516 2943 298544
rect 2971 298516 3019 298544
rect 2709 298482 3019 298516
rect 2709 298454 2757 298482
rect 2785 298454 2819 298482
rect 2847 298454 2881 298482
rect 2909 298454 2943 298482
rect 2971 298454 3019 298482
rect 2709 298420 3019 298454
rect 2709 298392 2757 298420
rect 2785 298392 2819 298420
rect 2847 298392 2881 298420
rect 2909 298392 2943 298420
rect 2971 298392 3019 298420
rect 2709 290175 3019 298392
rect 2709 290147 2757 290175
rect 2785 290147 2819 290175
rect 2847 290147 2881 290175
rect 2909 290147 2943 290175
rect 2971 290147 3019 290175
rect 2709 290113 3019 290147
rect 2709 290085 2757 290113
rect 2785 290085 2819 290113
rect 2847 290085 2881 290113
rect 2909 290085 2943 290113
rect 2971 290085 3019 290113
rect 2709 290051 3019 290085
rect 2709 290023 2757 290051
rect 2785 290023 2819 290051
rect 2847 290023 2881 290051
rect 2909 290023 2943 290051
rect 2971 290023 3019 290051
rect 2709 289989 3019 290023
rect 2709 289961 2757 289989
rect 2785 289961 2819 289989
rect 2847 289961 2881 289989
rect 2909 289961 2943 289989
rect 2971 289961 3019 289989
rect 2709 281175 3019 289961
rect 2709 281147 2757 281175
rect 2785 281147 2819 281175
rect 2847 281147 2881 281175
rect 2909 281147 2943 281175
rect 2971 281147 3019 281175
rect 2709 281113 3019 281147
rect 2709 281085 2757 281113
rect 2785 281085 2819 281113
rect 2847 281085 2881 281113
rect 2909 281085 2943 281113
rect 2971 281085 3019 281113
rect 2709 281051 3019 281085
rect 2709 281023 2757 281051
rect 2785 281023 2819 281051
rect 2847 281023 2881 281051
rect 2909 281023 2943 281051
rect 2971 281023 3019 281051
rect 2709 280989 3019 281023
rect 2709 280961 2757 280989
rect 2785 280961 2819 280989
rect 2847 280961 2881 280989
rect 2909 280961 2943 280989
rect 2971 280961 3019 280989
rect 2709 272175 3019 280961
rect 2709 272147 2757 272175
rect 2785 272147 2819 272175
rect 2847 272147 2881 272175
rect 2909 272147 2943 272175
rect 2971 272147 3019 272175
rect 2709 272113 3019 272147
rect 2709 272085 2757 272113
rect 2785 272085 2819 272113
rect 2847 272085 2881 272113
rect 2909 272085 2943 272113
rect 2971 272085 3019 272113
rect 2709 272051 3019 272085
rect 2709 272023 2757 272051
rect 2785 272023 2819 272051
rect 2847 272023 2881 272051
rect 2909 272023 2943 272051
rect 2971 272023 3019 272051
rect 2709 271989 3019 272023
rect 2709 271961 2757 271989
rect 2785 271961 2819 271989
rect 2847 271961 2881 271989
rect 2909 271961 2943 271989
rect 2971 271961 3019 271989
rect 2709 263175 3019 271961
rect 2709 263147 2757 263175
rect 2785 263147 2819 263175
rect 2847 263147 2881 263175
rect 2909 263147 2943 263175
rect 2971 263147 3019 263175
rect 2709 263113 3019 263147
rect 2709 263085 2757 263113
rect 2785 263085 2819 263113
rect 2847 263085 2881 263113
rect 2909 263085 2943 263113
rect 2971 263085 3019 263113
rect 2709 263051 3019 263085
rect 2709 263023 2757 263051
rect 2785 263023 2819 263051
rect 2847 263023 2881 263051
rect 2909 263023 2943 263051
rect 2971 263023 3019 263051
rect 2709 262989 3019 263023
rect 2709 262961 2757 262989
rect 2785 262961 2819 262989
rect 2847 262961 2881 262989
rect 2909 262961 2943 262989
rect 2971 262961 3019 262989
rect 2709 254175 3019 262961
rect 2709 254147 2757 254175
rect 2785 254147 2819 254175
rect 2847 254147 2881 254175
rect 2909 254147 2943 254175
rect 2971 254147 3019 254175
rect 2709 254113 3019 254147
rect 2709 254085 2757 254113
rect 2785 254085 2819 254113
rect 2847 254085 2881 254113
rect 2909 254085 2943 254113
rect 2971 254085 3019 254113
rect 2709 254051 3019 254085
rect 2709 254023 2757 254051
rect 2785 254023 2819 254051
rect 2847 254023 2881 254051
rect 2909 254023 2943 254051
rect 2971 254023 3019 254051
rect 2709 253989 3019 254023
rect 2709 253961 2757 253989
rect 2785 253961 2819 253989
rect 2847 253961 2881 253989
rect 2909 253961 2943 253989
rect 2971 253961 3019 253989
rect 2709 245175 3019 253961
rect 2709 245147 2757 245175
rect 2785 245147 2819 245175
rect 2847 245147 2881 245175
rect 2909 245147 2943 245175
rect 2971 245147 3019 245175
rect 2709 245113 3019 245147
rect 2709 245085 2757 245113
rect 2785 245085 2819 245113
rect 2847 245085 2881 245113
rect 2909 245085 2943 245113
rect 2971 245085 3019 245113
rect 2709 245051 3019 245085
rect 2709 245023 2757 245051
rect 2785 245023 2819 245051
rect 2847 245023 2881 245051
rect 2909 245023 2943 245051
rect 2971 245023 3019 245051
rect 2709 244989 3019 245023
rect 2709 244961 2757 244989
rect 2785 244961 2819 244989
rect 2847 244961 2881 244989
rect 2909 244961 2943 244989
rect 2971 244961 3019 244989
rect 2709 236175 3019 244961
rect 2709 236147 2757 236175
rect 2785 236147 2819 236175
rect 2847 236147 2881 236175
rect 2909 236147 2943 236175
rect 2971 236147 3019 236175
rect 2709 236113 3019 236147
rect 2709 236085 2757 236113
rect 2785 236085 2819 236113
rect 2847 236085 2881 236113
rect 2909 236085 2943 236113
rect 2971 236085 3019 236113
rect 2709 236051 3019 236085
rect 2709 236023 2757 236051
rect 2785 236023 2819 236051
rect 2847 236023 2881 236051
rect 2909 236023 2943 236051
rect 2971 236023 3019 236051
rect 2709 235989 3019 236023
rect 2709 235961 2757 235989
rect 2785 235961 2819 235989
rect 2847 235961 2881 235989
rect 2909 235961 2943 235989
rect 2971 235961 3019 235989
rect 2709 227175 3019 235961
rect 2709 227147 2757 227175
rect 2785 227147 2819 227175
rect 2847 227147 2881 227175
rect 2909 227147 2943 227175
rect 2971 227147 3019 227175
rect 2709 227113 3019 227147
rect 2709 227085 2757 227113
rect 2785 227085 2819 227113
rect 2847 227085 2881 227113
rect 2909 227085 2943 227113
rect 2971 227085 3019 227113
rect 2709 227051 3019 227085
rect 2709 227023 2757 227051
rect 2785 227023 2819 227051
rect 2847 227023 2881 227051
rect 2909 227023 2943 227051
rect 2971 227023 3019 227051
rect 2709 226989 3019 227023
rect 2709 226961 2757 226989
rect 2785 226961 2819 226989
rect 2847 226961 2881 226989
rect 2909 226961 2943 226989
rect 2971 226961 3019 226989
rect 2709 218175 3019 226961
rect 2709 218147 2757 218175
rect 2785 218147 2819 218175
rect 2847 218147 2881 218175
rect 2909 218147 2943 218175
rect 2971 218147 3019 218175
rect 2709 218113 3019 218147
rect 2709 218085 2757 218113
rect 2785 218085 2819 218113
rect 2847 218085 2881 218113
rect 2909 218085 2943 218113
rect 2971 218085 3019 218113
rect 2709 218051 3019 218085
rect 2709 218023 2757 218051
rect 2785 218023 2819 218051
rect 2847 218023 2881 218051
rect 2909 218023 2943 218051
rect 2971 218023 3019 218051
rect 2709 217989 3019 218023
rect 2709 217961 2757 217989
rect 2785 217961 2819 217989
rect 2847 217961 2881 217989
rect 2909 217961 2943 217989
rect 2971 217961 3019 217989
rect 2709 209175 3019 217961
rect 2709 209147 2757 209175
rect 2785 209147 2819 209175
rect 2847 209147 2881 209175
rect 2909 209147 2943 209175
rect 2971 209147 3019 209175
rect 2709 209113 3019 209147
rect 2709 209085 2757 209113
rect 2785 209085 2819 209113
rect 2847 209085 2881 209113
rect 2909 209085 2943 209113
rect 2971 209085 3019 209113
rect 2709 209051 3019 209085
rect 2709 209023 2757 209051
rect 2785 209023 2819 209051
rect 2847 209023 2881 209051
rect 2909 209023 2943 209051
rect 2971 209023 3019 209051
rect 2709 208989 3019 209023
rect 2709 208961 2757 208989
rect 2785 208961 2819 208989
rect 2847 208961 2881 208989
rect 2909 208961 2943 208989
rect 2971 208961 3019 208989
rect 2709 200175 3019 208961
rect 2709 200147 2757 200175
rect 2785 200147 2819 200175
rect 2847 200147 2881 200175
rect 2909 200147 2943 200175
rect 2971 200147 3019 200175
rect 2709 200113 3019 200147
rect 2709 200085 2757 200113
rect 2785 200085 2819 200113
rect 2847 200085 2881 200113
rect 2909 200085 2943 200113
rect 2971 200085 3019 200113
rect 2709 200051 3019 200085
rect 2709 200023 2757 200051
rect 2785 200023 2819 200051
rect 2847 200023 2881 200051
rect 2909 200023 2943 200051
rect 2971 200023 3019 200051
rect 2709 199989 3019 200023
rect 2709 199961 2757 199989
rect 2785 199961 2819 199989
rect 2847 199961 2881 199989
rect 2909 199961 2943 199989
rect 2971 199961 3019 199989
rect 2709 191175 3019 199961
rect 2709 191147 2757 191175
rect 2785 191147 2819 191175
rect 2847 191147 2881 191175
rect 2909 191147 2943 191175
rect 2971 191147 3019 191175
rect 2709 191113 3019 191147
rect 2709 191085 2757 191113
rect 2785 191085 2819 191113
rect 2847 191085 2881 191113
rect 2909 191085 2943 191113
rect 2971 191085 3019 191113
rect 2709 191051 3019 191085
rect 2709 191023 2757 191051
rect 2785 191023 2819 191051
rect 2847 191023 2881 191051
rect 2909 191023 2943 191051
rect 2971 191023 3019 191051
rect 2709 190989 3019 191023
rect 2709 190961 2757 190989
rect 2785 190961 2819 190989
rect 2847 190961 2881 190989
rect 2909 190961 2943 190989
rect 2971 190961 3019 190989
rect 2709 182175 3019 190961
rect 2709 182147 2757 182175
rect 2785 182147 2819 182175
rect 2847 182147 2881 182175
rect 2909 182147 2943 182175
rect 2971 182147 3019 182175
rect 2709 182113 3019 182147
rect 2709 182085 2757 182113
rect 2785 182085 2819 182113
rect 2847 182085 2881 182113
rect 2909 182085 2943 182113
rect 2971 182085 3019 182113
rect 2709 182051 3019 182085
rect 2709 182023 2757 182051
rect 2785 182023 2819 182051
rect 2847 182023 2881 182051
rect 2909 182023 2943 182051
rect 2971 182023 3019 182051
rect 2709 181989 3019 182023
rect 2709 181961 2757 181989
rect 2785 181961 2819 181989
rect 2847 181961 2881 181989
rect 2909 181961 2943 181989
rect 2971 181961 3019 181989
rect 2709 173175 3019 181961
rect 4569 299086 4879 299134
rect 4569 299058 4617 299086
rect 4645 299058 4679 299086
rect 4707 299058 4741 299086
rect 4769 299058 4803 299086
rect 4831 299058 4879 299086
rect 4569 299024 4879 299058
rect 4569 298996 4617 299024
rect 4645 298996 4679 299024
rect 4707 298996 4741 299024
rect 4769 298996 4803 299024
rect 4831 298996 4879 299024
rect 4569 298962 4879 298996
rect 4569 298934 4617 298962
rect 4645 298934 4679 298962
rect 4707 298934 4741 298962
rect 4769 298934 4803 298962
rect 4831 298934 4879 298962
rect 4569 298900 4879 298934
rect 4569 298872 4617 298900
rect 4645 298872 4679 298900
rect 4707 298872 4741 298900
rect 4769 298872 4803 298900
rect 4831 298872 4879 298900
rect 4569 293175 4879 298872
rect 4569 293147 4617 293175
rect 4645 293147 4679 293175
rect 4707 293147 4741 293175
rect 4769 293147 4803 293175
rect 4831 293147 4879 293175
rect 4569 293113 4879 293147
rect 4569 293085 4617 293113
rect 4645 293085 4679 293113
rect 4707 293085 4741 293113
rect 4769 293085 4803 293113
rect 4831 293085 4879 293113
rect 4569 293051 4879 293085
rect 4569 293023 4617 293051
rect 4645 293023 4679 293051
rect 4707 293023 4741 293051
rect 4769 293023 4803 293051
rect 4831 293023 4879 293051
rect 4569 292989 4879 293023
rect 4569 292961 4617 292989
rect 4645 292961 4679 292989
rect 4707 292961 4741 292989
rect 4769 292961 4803 292989
rect 4831 292961 4879 292989
rect 4569 284175 4879 292961
rect 4569 284147 4617 284175
rect 4645 284147 4679 284175
rect 4707 284147 4741 284175
rect 4769 284147 4803 284175
rect 4831 284147 4879 284175
rect 4569 284113 4879 284147
rect 4569 284085 4617 284113
rect 4645 284085 4679 284113
rect 4707 284085 4741 284113
rect 4769 284085 4803 284113
rect 4831 284085 4879 284113
rect 4569 284051 4879 284085
rect 4569 284023 4617 284051
rect 4645 284023 4679 284051
rect 4707 284023 4741 284051
rect 4769 284023 4803 284051
rect 4831 284023 4879 284051
rect 4569 283989 4879 284023
rect 4569 283961 4617 283989
rect 4645 283961 4679 283989
rect 4707 283961 4741 283989
rect 4769 283961 4803 283989
rect 4831 283961 4879 283989
rect 4569 275175 4879 283961
rect 4569 275147 4617 275175
rect 4645 275147 4679 275175
rect 4707 275147 4741 275175
rect 4769 275147 4803 275175
rect 4831 275147 4879 275175
rect 4569 275113 4879 275147
rect 4569 275085 4617 275113
rect 4645 275085 4679 275113
rect 4707 275085 4741 275113
rect 4769 275085 4803 275113
rect 4831 275085 4879 275113
rect 4569 275051 4879 275085
rect 4569 275023 4617 275051
rect 4645 275023 4679 275051
rect 4707 275023 4741 275051
rect 4769 275023 4803 275051
rect 4831 275023 4879 275051
rect 4569 274989 4879 275023
rect 4569 274961 4617 274989
rect 4645 274961 4679 274989
rect 4707 274961 4741 274989
rect 4769 274961 4803 274989
rect 4831 274961 4879 274989
rect 4569 266175 4879 274961
rect 4569 266147 4617 266175
rect 4645 266147 4679 266175
rect 4707 266147 4741 266175
rect 4769 266147 4803 266175
rect 4831 266147 4879 266175
rect 4569 266113 4879 266147
rect 4569 266085 4617 266113
rect 4645 266085 4679 266113
rect 4707 266085 4741 266113
rect 4769 266085 4803 266113
rect 4831 266085 4879 266113
rect 4569 266051 4879 266085
rect 4569 266023 4617 266051
rect 4645 266023 4679 266051
rect 4707 266023 4741 266051
rect 4769 266023 4803 266051
rect 4831 266023 4879 266051
rect 4569 265989 4879 266023
rect 4569 265961 4617 265989
rect 4645 265961 4679 265989
rect 4707 265961 4741 265989
rect 4769 265961 4803 265989
rect 4831 265961 4879 265989
rect 4569 257175 4879 265961
rect 4569 257147 4617 257175
rect 4645 257147 4679 257175
rect 4707 257147 4741 257175
rect 4769 257147 4803 257175
rect 4831 257147 4879 257175
rect 4569 257113 4879 257147
rect 4569 257085 4617 257113
rect 4645 257085 4679 257113
rect 4707 257085 4741 257113
rect 4769 257085 4803 257113
rect 4831 257085 4879 257113
rect 4569 257051 4879 257085
rect 4569 257023 4617 257051
rect 4645 257023 4679 257051
rect 4707 257023 4741 257051
rect 4769 257023 4803 257051
rect 4831 257023 4879 257051
rect 4569 256989 4879 257023
rect 4569 256961 4617 256989
rect 4645 256961 4679 256989
rect 4707 256961 4741 256989
rect 4769 256961 4803 256989
rect 4831 256961 4879 256989
rect 4569 248175 4879 256961
rect 4569 248147 4617 248175
rect 4645 248147 4679 248175
rect 4707 248147 4741 248175
rect 4769 248147 4803 248175
rect 4831 248147 4879 248175
rect 4569 248113 4879 248147
rect 4569 248085 4617 248113
rect 4645 248085 4679 248113
rect 4707 248085 4741 248113
rect 4769 248085 4803 248113
rect 4831 248085 4879 248113
rect 4569 248051 4879 248085
rect 4569 248023 4617 248051
rect 4645 248023 4679 248051
rect 4707 248023 4741 248051
rect 4769 248023 4803 248051
rect 4831 248023 4879 248051
rect 4569 247989 4879 248023
rect 4569 247961 4617 247989
rect 4645 247961 4679 247989
rect 4707 247961 4741 247989
rect 4769 247961 4803 247989
rect 4831 247961 4879 247989
rect 4569 239175 4879 247961
rect 4569 239147 4617 239175
rect 4645 239147 4679 239175
rect 4707 239147 4741 239175
rect 4769 239147 4803 239175
rect 4831 239147 4879 239175
rect 4569 239113 4879 239147
rect 4569 239085 4617 239113
rect 4645 239085 4679 239113
rect 4707 239085 4741 239113
rect 4769 239085 4803 239113
rect 4831 239085 4879 239113
rect 4569 239051 4879 239085
rect 4569 239023 4617 239051
rect 4645 239023 4679 239051
rect 4707 239023 4741 239051
rect 4769 239023 4803 239051
rect 4831 239023 4879 239051
rect 4569 238989 4879 239023
rect 4569 238961 4617 238989
rect 4645 238961 4679 238989
rect 4707 238961 4741 238989
rect 4769 238961 4803 238989
rect 4831 238961 4879 238989
rect 4569 230175 4879 238961
rect 4569 230147 4617 230175
rect 4645 230147 4679 230175
rect 4707 230147 4741 230175
rect 4769 230147 4803 230175
rect 4831 230147 4879 230175
rect 4569 230113 4879 230147
rect 4569 230085 4617 230113
rect 4645 230085 4679 230113
rect 4707 230085 4741 230113
rect 4769 230085 4803 230113
rect 4831 230085 4879 230113
rect 4569 230051 4879 230085
rect 4569 230023 4617 230051
rect 4645 230023 4679 230051
rect 4707 230023 4741 230051
rect 4769 230023 4803 230051
rect 4831 230023 4879 230051
rect 4569 229989 4879 230023
rect 4569 229961 4617 229989
rect 4645 229961 4679 229989
rect 4707 229961 4741 229989
rect 4769 229961 4803 229989
rect 4831 229961 4879 229989
rect 4569 221175 4879 229961
rect 4569 221147 4617 221175
rect 4645 221147 4679 221175
rect 4707 221147 4741 221175
rect 4769 221147 4803 221175
rect 4831 221147 4879 221175
rect 4569 221113 4879 221147
rect 4569 221085 4617 221113
rect 4645 221085 4679 221113
rect 4707 221085 4741 221113
rect 4769 221085 4803 221113
rect 4831 221085 4879 221113
rect 4569 221051 4879 221085
rect 4569 221023 4617 221051
rect 4645 221023 4679 221051
rect 4707 221023 4741 221051
rect 4769 221023 4803 221051
rect 4831 221023 4879 221051
rect 4569 220989 4879 221023
rect 4569 220961 4617 220989
rect 4645 220961 4679 220989
rect 4707 220961 4741 220989
rect 4769 220961 4803 220989
rect 4831 220961 4879 220989
rect 4569 212175 4879 220961
rect 4569 212147 4617 212175
rect 4645 212147 4679 212175
rect 4707 212147 4741 212175
rect 4769 212147 4803 212175
rect 4831 212147 4879 212175
rect 4569 212113 4879 212147
rect 4569 212085 4617 212113
rect 4645 212085 4679 212113
rect 4707 212085 4741 212113
rect 4769 212085 4803 212113
rect 4831 212085 4879 212113
rect 4569 212051 4879 212085
rect 4569 212023 4617 212051
rect 4645 212023 4679 212051
rect 4707 212023 4741 212051
rect 4769 212023 4803 212051
rect 4831 212023 4879 212051
rect 4569 211989 4879 212023
rect 4569 211961 4617 211989
rect 4645 211961 4679 211989
rect 4707 211961 4741 211989
rect 4769 211961 4803 211989
rect 4831 211961 4879 211989
rect 4569 203175 4879 211961
rect 4569 203147 4617 203175
rect 4645 203147 4679 203175
rect 4707 203147 4741 203175
rect 4769 203147 4803 203175
rect 4831 203147 4879 203175
rect 4569 203113 4879 203147
rect 4569 203085 4617 203113
rect 4645 203085 4679 203113
rect 4707 203085 4741 203113
rect 4769 203085 4803 203113
rect 4831 203085 4879 203113
rect 4569 203051 4879 203085
rect 4569 203023 4617 203051
rect 4645 203023 4679 203051
rect 4707 203023 4741 203051
rect 4769 203023 4803 203051
rect 4831 203023 4879 203051
rect 4569 202989 4879 203023
rect 4569 202961 4617 202989
rect 4645 202961 4679 202989
rect 4707 202961 4741 202989
rect 4769 202961 4803 202989
rect 4831 202961 4879 202989
rect 4569 194175 4879 202961
rect 4569 194147 4617 194175
rect 4645 194147 4679 194175
rect 4707 194147 4741 194175
rect 4769 194147 4803 194175
rect 4831 194147 4879 194175
rect 4569 194113 4879 194147
rect 4569 194085 4617 194113
rect 4645 194085 4679 194113
rect 4707 194085 4741 194113
rect 4769 194085 4803 194113
rect 4831 194085 4879 194113
rect 4569 194051 4879 194085
rect 4569 194023 4617 194051
rect 4645 194023 4679 194051
rect 4707 194023 4741 194051
rect 4769 194023 4803 194051
rect 4831 194023 4879 194051
rect 4569 193989 4879 194023
rect 4569 193961 4617 193989
rect 4645 193961 4679 193989
rect 4707 193961 4741 193989
rect 4769 193961 4803 193989
rect 4831 193961 4879 193989
rect 4569 185175 4879 193961
rect 4569 185147 4617 185175
rect 4645 185147 4679 185175
rect 4707 185147 4741 185175
rect 4769 185147 4803 185175
rect 4831 185147 4879 185175
rect 4569 185113 4879 185147
rect 4569 185085 4617 185113
rect 4645 185085 4679 185113
rect 4707 185085 4741 185113
rect 4769 185085 4803 185113
rect 4831 185085 4879 185113
rect 4569 185051 4879 185085
rect 4569 185023 4617 185051
rect 4645 185023 4679 185051
rect 4707 185023 4741 185051
rect 4769 185023 4803 185051
rect 4831 185023 4879 185051
rect 4569 184989 4879 185023
rect 4569 184961 4617 184989
rect 4645 184961 4679 184989
rect 4707 184961 4741 184989
rect 4769 184961 4803 184989
rect 4831 184961 4879 184989
rect 4569 176175 4879 184961
rect 4569 176147 4617 176175
rect 4645 176147 4679 176175
rect 4707 176147 4741 176175
rect 4769 176147 4803 176175
rect 4831 176147 4879 176175
rect 4569 176113 4879 176147
rect 4569 176085 4617 176113
rect 4645 176085 4679 176113
rect 4707 176085 4741 176113
rect 4769 176085 4803 176113
rect 4831 176085 4879 176113
rect 4569 176051 4879 176085
rect 4569 176023 4617 176051
rect 4645 176023 4679 176051
rect 4707 176023 4741 176051
rect 4769 176023 4803 176051
rect 4831 176023 4879 176051
rect 4569 175989 4879 176023
rect 4569 175961 4617 175989
rect 4645 175961 4679 175989
rect 4707 175961 4741 175989
rect 4769 175961 4803 175989
rect 4831 175961 4879 175989
rect 2709 173147 2757 173175
rect 2785 173147 2819 173175
rect 2847 173147 2881 173175
rect 2909 173147 2943 173175
rect 2971 173147 3019 173175
rect 2709 173113 3019 173147
rect 2709 173085 2757 173113
rect 2785 173085 2819 173113
rect 2847 173085 2881 173113
rect 2909 173085 2943 173113
rect 2971 173085 3019 173113
rect 2709 173051 3019 173085
rect 2709 173023 2757 173051
rect 2785 173023 2819 173051
rect 2847 173023 2881 173051
rect 2909 173023 2943 173051
rect 2971 173023 3019 173051
rect 2709 172989 3019 173023
rect 2709 172961 2757 172989
rect 2785 172961 2819 172989
rect 2847 172961 2881 172989
rect 2909 172961 2943 172989
rect 2971 172961 3019 172989
rect 2709 164175 3019 172961
rect 3766 173250 3794 173255
rect 3766 166698 3794 173222
rect 3766 166665 3794 166670
rect 4569 167175 4879 175961
rect 18069 298606 18379 299134
rect 18069 298578 18117 298606
rect 18145 298578 18179 298606
rect 18207 298578 18241 298606
rect 18269 298578 18303 298606
rect 18331 298578 18379 298606
rect 18069 298544 18379 298578
rect 18069 298516 18117 298544
rect 18145 298516 18179 298544
rect 18207 298516 18241 298544
rect 18269 298516 18303 298544
rect 18331 298516 18379 298544
rect 18069 298482 18379 298516
rect 18069 298454 18117 298482
rect 18145 298454 18179 298482
rect 18207 298454 18241 298482
rect 18269 298454 18303 298482
rect 18331 298454 18379 298482
rect 18069 298420 18379 298454
rect 18069 298392 18117 298420
rect 18145 298392 18179 298420
rect 18207 298392 18241 298420
rect 18269 298392 18303 298420
rect 18331 298392 18379 298420
rect 18069 290175 18379 298392
rect 18069 290147 18117 290175
rect 18145 290147 18179 290175
rect 18207 290147 18241 290175
rect 18269 290147 18303 290175
rect 18331 290147 18379 290175
rect 18069 290113 18379 290147
rect 18069 290085 18117 290113
rect 18145 290085 18179 290113
rect 18207 290085 18241 290113
rect 18269 290085 18303 290113
rect 18331 290085 18379 290113
rect 18069 290051 18379 290085
rect 18069 290023 18117 290051
rect 18145 290023 18179 290051
rect 18207 290023 18241 290051
rect 18269 290023 18303 290051
rect 18331 290023 18379 290051
rect 18069 289989 18379 290023
rect 18069 289961 18117 289989
rect 18145 289961 18179 289989
rect 18207 289961 18241 289989
rect 18269 289961 18303 289989
rect 18331 289961 18379 289989
rect 18069 281175 18379 289961
rect 18069 281147 18117 281175
rect 18145 281147 18179 281175
rect 18207 281147 18241 281175
rect 18269 281147 18303 281175
rect 18331 281147 18379 281175
rect 18069 281113 18379 281147
rect 18069 281085 18117 281113
rect 18145 281085 18179 281113
rect 18207 281085 18241 281113
rect 18269 281085 18303 281113
rect 18331 281085 18379 281113
rect 18069 281051 18379 281085
rect 18069 281023 18117 281051
rect 18145 281023 18179 281051
rect 18207 281023 18241 281051
rect 18269 281023 18303 281051
rect 18331 281023 18379 281051
rect 18069 280989 18379 281023
rect 18069 280961 18117 280989
rect 18145 280961 18179 280989
rect 18207 280961 18241 280989
rect 18269 280961 18303 280989
rect 18331 280961 18379 280989
rect 18069 272175 18379 280961
rect 18069 272147 18117 272175
rect 18145 272147 18179 272175
rect 18207 272147 18241 272175
rect 18269 272147 18303 272175
rect 18331 272147 18379 272175
rect 18069 272113 18379 272147
rect 18069 272085 18117 272113
rect 18145 272085 18179 272113
rect 18207 272085 18241 272113
rect 18269 272085 18303 272113
rect 18331 272085 18379 272113
rect 18069 272051 18379 272085
rect 18069 272023 18117 272051
rect 18145 272023 18179 272051
rect 18207 272023 18241 272051
rect 18269 272023 18303 272051
rect 18331 272023 18379 272051
rect 18069 271989 18379 272023
rect 18069 271961 18117 271989
rect 18145 271961 18179 271989
rect 18207 271961 18241 271989
rect 18269 271961 18303 271989
rect 18331 271961 18379 271989
rect 18069 263175 18379 271961
rect 18069 263147 18117 263175
rect 18145 263147 18179 263175
rect 18207 263147 18241 263175
rect 18269 263147 18303 263175
rect 18331 263147 18379 263175
rect 18069 263113 18379 263147
rect 18069 263085 18117 263113
rect 18145 263085 18179 263113
rect 18207 263085 18241 263113
rect 18269 263085 18303 263113
rect 18331 263085 18379 263113
rect 18069 263051 18379 263085
rect 18069 263023 18117 263051
rect 18145 263023 18179 263051
rect 18207 263023 18241 263051
rect 18269 263023 18303 263051
rect 18331 263023 18379 263051
rect 18069 262989 18379 263023
rect 18069 262961 18117 262989
rect 18145 262961 18179 262989
rect 18207 262961 18241 262989
rect 18269 262961 18303 262989
rect 18331 262961 18379 262989
rect 18069 254175 18379 262961
rect 18069 254147 18117 254175
rect 18145 254147 18179 254175
rect 18207 254147 18241 254175
rect 18269 254147 18303 254175
rect 18331 254147 18379 254175
rect 18069 254113 18379 254147
rect 18069 254085 18117 254113
rect 18145 254085 18179 254113
rect 18207 254085 18241 254113
rect 18269 254085 18303 254113
rect 18331 254085 18379 254113
rect 18069 254051 18379 254085
rect 18069 254023 18117 254051
rect 18145 254023 18179 254051
rect 18207 254023 18241 254051
rect 18269 254023 18303 254051
rect 18331 254023 18379 254051
rect 18069 253989 18379 254023
rect 18069 253961 18117 253989
rect 18145 253961 18179 253989
rect 18207 253961 18241 253989
rect 18269 253961 18303 253989
rect 18331 253961 18379 253989
rect 18069 245175 18379 253961
rect 18069 245147 18117 245175
rect 18145 245147 18179 245175
rect 18207 245147 18241 245175
rect 18269 245147 18303 245175
rect 18331 245147 18379 245175
rect 18069 245113 18379 245147
rect 18069 245085 18117 245113
rect 18145 245085 18179 245113
rect 18207 245085 18241 245113
rect 18269 245085 18303 245113
rect 18331 245085 18379 245113
rect 18069 245051 18379 245085
rect 18069 245023 18117 245051
rect 18145 245023 18179 245051
rect 18207 245023 18241 245051
rect 18269 245023 18303 245051
rect 18331 245023 18379 245051
rect 18069 244989 18379 245023
rect 18069 244961 18117 244989
rect 18145 244961 18179 244989
rect 18207 244961 18241 244989
rect 18269 244961 18303 244989
rect 18331 244961 18379 244989
rect 18069 236175 18379 244961
rect 18069 236147 18117 236175
rect 18145 236147 18179 236175
rect 18207 236147 18241 236175
rect 18269 236147 18303 236175
rect 18331 236147 18379 236175
rect 18069 236113 18379 236147
rect 18069 236085 18117 236113
rect 18145 236085 18179 236113
rect 18207 236085 18241 236113
rect 18269 236085 18303 236113
rect 18331 236085 18379 236113
rect 18069 236051 18379 236085
rect 18069 236023 18117 236051
rect 18145 236023 18179 236051
rect 18207 236023 18241 236051
rect 18269 236023 18303 236051
rect 18331 236023 18379 236051
rect 18069 235989 18379 236023
rect 18069 235961 18117 235989
rect 18145 235961 18179 235989
rect 18207 235961 18241 235989
rect 18269 235961 18303 235989
rect 18331 235961 18379 235989
rect 18069 227175 18379 235961
rect 18069 227147 18117 227175
rect 18145 227147 18179 227175
rect 18207 227147 18241 227175
rect 18269 227147 18303 227175
rect 18331 227147 18379 227175
rect 18069 227113 18379 227147
rect 18069 227085 18117 227113
rect 18145 227085 18179 227113
rect 18207 227085 18241 227113
rect 18269 227085 18303 227113
rect 18331 227085 18379 227113
rect 18069 227051 18379 227085
rect 18069 227023 18117 227051
rect 18145 227023 18179 227051
rect 18207 227023 18241 227051
rect 18269 227023 18303 227051
rect 18331 227023 18379 227051
rect 18069 226989 18379 227023
rect 18069 226961 18117 226989
rect 18145 226961 18179 226989
rect 18207 226961 18241 226989
rect 18269 226961 18303 226989
rect 18331 226961 18379 226989
rect 18069 218175 18379 226961
rect 18069 218147 18117 218175
rect 18145 218147 18179 218175
rect 18207 218147 18241 218175
rect 18269 218147 18303 218175
rect 18331 218147 18379 218175
rect 18069 218113 18379 218147
rect 18069 218085 18117 218113
rect 18145 218085 18179 218113
rect 18207 218085 18241 218113
rect 18269 218085 18303 218113
rect 18331 218085 18379 218113
rect 18069 218051 18379 218085
rect 18069 218023 18117 218051
rect 18145 218023 18179 218051
rect 18207 218023 18241 218051
rect 18269 218023 18303 218051
rect 18331 218023 18379 218051
rect 18069 217989 18379 218023
rect 18069 217961 18117 217989
rect 18145 217961 18179 217989
rect 18207 217961 18241 217989
rect 18269 217961 18303 217989
rect 18331 217961 18379 217989
rect 18069 209175 18379 217961
rect 18069 209147 18117 209175
rect 18145 209147 18179 209175
rect 18207 209147 18241 209175
rect 18269 209147 18303 209175
rect 18331 209147 18379 209175
rect 18069 209113 18379 209147
rect 18069 209085 18117 209113
rect 18145 209085 18179 209113
rect 18207 209085 18241 209113
rect 18269 209085 18303 209113
rect 18331 209085 18379 209113
rect 18069 209051 18379 209085
rect 18069 209023 18117 209051
rect 18145 209023 18179 209051
rect 18207 209023 18241 209051
rect 18269 209023 18303 209051
rect 18331 209023 18379 209051
rect 18069 208989 18379 209023
rect 18069 208961 18117 208989
rect 18145 208961 18179 208989
rect 18207 208961 18241 208989
rect 18269 208961 18303 208989
rect 18331 208961 18379 208989
rect 18069 200175 18379 208961
rect 18069 200147 18117 200175
rect 18145 200147 18179 200175
rect 18207 200147 18241 200175
rect 18269 200147 18303 200175
rect 18331 200147 18379 200175
rect 18069 200113 18379 200147
rect 18069 200085 18117 200113
rect 18145 200085 18179 200113
rect 18207 200085 18241 200113
rect 18269 200085 18303 200113
rect 18331 200085 18379 200113
rect 18069 200051 18379 200085
rect 18069 200023 18117 200051
rect 18145 200023 18179 200051
rect 18207 200023 18241 200051
rect 18269 200023 18303 200051
rect 18331 200023 18379 200051
rect 18069 199989 18379 200023
rect 18069 199961 18117 199989
rect 18145 199961 18179 199989
rect 18207 199961 18241 199989
rect 18269 199961 18303 199989
rect 18331 199961 18379 199989
rect 18069 191175 18379 199961
rect 18069 191147 18117 191175
rect 18145 191147 18179 191175
rect 18207 191147 18241 191175
rect 18269 191147 18303 191175
rect 18331 191147 18379 191175
rect 18069 191113 18379 191147
rect 18069 191085 18117 191113
rect 18145 191085 18179 191113
rect 18207 191085 18241 191113
rect 18269 191085 18303 191113
rect 18331 191085 18379 191113
rect 18069 191051 18379 191085
rect 18069 191023 18117 191051
rect 18145 191023 18179 191051
rect 18207 191023 18241 191051
rect 18269 191023 18303 191051
rect 18331 191023 18379 191051
rect 18069 190989 18379 191023
rect 18069 190961 18117 190989
rect 18145 190961 18179 190989
rect 18207 190961 18241 190989
rect 18269 190961 18303 190989
rect 18331 190961 18379 190989
rect 18069 182175 18379 190961
rect 18069 182147 18117 182175
rect 18145 182147 18179 182175
rect 18207 182147 18241 182175
rect 18269 182147 18303 182175
rect 18331 182147 18379 182175
rect 18069 182113 18379 182147
rect 18069 182085 18117 182113
rect 18145 182085 18179 182113
rect 18207 182085 18241 182113
rect 18269 182085 18303 182113
rect 18331 182085 18379 182113
rect 18069 182051 18379 182085
rect 18069 182023 18117 182051
rect 18145 182023 18179 182051
rect 18207 182023 18241 182051
rect 18269 182023 18303 182051
rect 18331 182023 18379 182051
rect 18069 181989 18379 182023
rect 18069 181961 18117 181989
rect 18145 181961 18179 181989
rect 18207 181961 18241 181989
rect 18269 181961 18303 181989
rect 18331 181961 18379 181989
rect 8224 173175 8384 173192
rect 8224 173147 8259 173175
rect 8287 173147 8321 173175
rect 8349 173147 8384 173175
rect 8224 173113 8384 173147
rect 8224 173085 8259 173113
rect 8287 173085 8321 173113
rect 8349 173085 8384 173113
rect 8224 173051 8384 173085
rect 8224 173023 8259 173051
rect 8287 173023 8321 173051
rect 8349 173023 8384 173051
rect 8224 172989 8384 173023
rect 8224 172961 8259 172989
rect 8287 172961 8321 172989
rect 8349 172961 8384 172989
rect 8224 172944 8384 172961
rect 18069 173175 18379 181961
rect 18069 173147 18117 173175
rect 18145 173147 18179 173175
rect 18207 173147 18241 173175
rect 18269 173147 18303 173175
rect 18331 173147 18379 173175
rect 18069 173113 18379 173147
rect 18069 173085 18117 173113
rect 18145 173085 18179 173113
rect 18207 173085 18241 173113
rect 18269 173085 18303 173113
rect 18331 173085 18379 173113
rect 18069 173051 18379 173085
rect 18069 173023 18117 173051
rect 18145 173023 18179 173051
rect 18207 173023 18241 173051
rect 18269 173023 18303 173051
rect 18331 173023 18379 173051
rect 18069 172989 18379 173023
rect 18069 172961 18117 172989
rect 18145 172961 18179 172989
rect 18207 172961 18241 172989
rect 18269 172961 18303 172989
rect 18331 172961 18379 172989
rect 4569 167147 4617 167175
rect 4645 167147 4679 167175
rect 4707 167147 4741 167175
rect 4769 167147 4803 167175
rect 4831 167147 4879 167175
rect 4569 167113 4879 167147
rect 4569 167085 4617 167113
rect 4645 167085 4679 167113
rect 4707 167085 4741 167113
rect 4769 167085 4803 167113
rect 4831 167085 4879 167113
rect 4569 167051 4879 167085
rect 4569 167023 4617 167051
rect 4645 167023 4679 167051
rect 4707 167023 4741 167051
rect 4769 167023 4803 167051
rect 4831 167023 4879 167051
rect 4569 166989 4879 167023
rect 4569 166961 4617 166989
rect 4645 166961 4679 166989
rect 4707 166961 4741 166989
rect 4769 166961 4803 166989
rect 4831 166961 4879 166989
rect 2709 164147 2757 164175
rect 2785 164147 2819 164175
rect 2847 164147 2881 164175
rect 2909 164147 2943 164175
rect 2971 164147 3019 164175
rect 2709 164113 3019 164147
rect 2709 164085 2757 164113
rect 2785 164085 2819 164113
rect 2847 164085 2881 164113
rect 2909 164085 2943 164113
rect 2971 164085 3019 164113
rect 2709 164051 3019 164085
rect 2709 164023 2757 164051
rect 2785 164023 2819 164051
rect 2847 164023 2881 164051
rect 2909 164023 2943 164051
rect 2971 164023 3019 164051
rect 2709 163989 3019 164023
rect 2709 163961 2757 163989
rect 2785 163961 2819 163989
rect 2847 163961 2881 163989
rect 2909 163961 2943 163989
rect 2971 163961 3019 163989
rect 2709 155175 3019 163961
rect 3766 165970 3794 165975
rect 3766 159586 3794 165942
rect 3766 159553 3794 159558
rect 2709 155147 2757 155175
rect 2785 155147 2819 155175
rect 2847 155147 2881 155175
rect 2909 155147 2943 155175
rect 2971 155147 3019 155175
rect 2709 155113 3019 155147
rect 2709 155085 2757 155113
rect 2785 155085 2819 155113
rect 2847 155085 2881 155113
rect 2909 155085 2943 155113
rect 2971 155085 3019 155113
rect 2709 155051 3019 155085
rect 2709 155023 2757 155051
rect 2785 155023 2819 155051
rect 2847 155023 2881 155051
rect 2909 155023 2943 155051
rect 2971 155023 3019 155051
rect 2709 154989 3019 155023
rect 2709 154961 2757 154989
rect 2785 154961 2819 154989
rect 2847 154961 2881 154989
rect 2909 154961 2943 154989
rect 2971 154961 3019 154989
rect 2709 146175 3019 154961
rect 3766 158690 3794 158695
rect 3766 152586 3794 158662
rect 3766 152553 3794 152558
rect 4569 158175 4879 166961
rect 15904 167175 16064 167192
rect 15904 167147 15939 167175
rect 15967 167147 16001 167175
rect 16029 167147 16064 167175
rect 15904 167113 16064 167147
rect 15904 167085 15939 167113
rect 15967 167085 16001 167113
rect 16029 167085 16064 167113
rect 15904 167051 16064 167085
rect 15904 167023 15939 167051
rect 15967 167023 16001 167051
rect 16029 167023 16064 167051
rect 15904 166989 16064 167023
rect 15904 166961 15939 166989
rect 15967 166961 16001 166989
rect 16029 166961 16064 166989
rect 15904 166944 16064 166961
rect 8224 164175 8384 164192
rect 8224 164147 8259 164175
rect 8287 164147 8321 164175
rect 8349 164147 8384 164175
rect 8224 164113 8384 164147
rect 8224 164085 8259 164113
rect 8287 164085 8321 164113
rect 8349 164085 8384 164113
rect 8224 164051 8384 164085
rect 8224 164023 8259 164051
rect 8287 164023 8321 164051
rect 8349 164023 8384 164051
rect 8224 163989 8384 164023
rect 8224 163961 8259 163989
rect 8287 163961 8321 163989
rect 8349 163961 8384 163989
rect 8224 163944 8384 163961
rect 18069 164175 18379 172961
rect 18069 164147 18117 164175
rect 18145 164147 18179 164175
rect 18207 164147 18241 164175
rect 18269 164147 18303 164175
rect 18331 164147 18379 164175
rect 18069 164113 18379 164147
rect 18069 164085 18117 164113
rect 18145 164085 18179 164113
rect 18207 164085 18241 164113
rect 18269 164085 18303 164113
rect 18331 164085 18379 164113
rect 18069 164051 18379 164085
rect 18069 164023 18117 164051
rect 18145 164023 18179 164051
rect 18207 164023 18241 164051
rect 18269 164023 18303 164051
rect 18331 164023 18379 164051
rect 18069 163989 18379 164023
rect 18069 163961 18117 163989
rect 18145 163961 18179 163989
rect 18207 163961 18241 163989
rect 18269 163961 18303 163989
rect 18331 163961 18379 163989
rect 4569 158147 4617 158175
rect 4645 158147 4679 158175
rect 4707 158147 4741 158175
rect 4769 158147 4803 158175
rect 4831 158147 4879 158175
rect 4569 158113 4879 158147
rect 4569 158085 4617 158113
rect 4645 158085 4679 158113
rect 4707 158085 4741 158113
rect 4769 158085 4803 158113
rect 4831 158085 4879 158113
rect 4569 158051 4879 158085
rect 4569 158023 4617 158051
rect 4645 158023 4679 158051
rect 4707 158023 4741 158051
rect 4769 158023 4803 158051
rect 4831 158023 4879 158051
rect 4569 157989 4879 158023
rect 4569 157961 4617 157989
rect 4645 157961 4679 157989
rect 4707 157961 4741 157989
rect 4769 157961 4803 157989
rect 4831 157961 4879 157989
rect 2709 146147 2757 146175
rect 2785 146147 2819 146175
rect 2847 146147 2881 146175
rect 2909 146147 2943 146175
rect 2971 146147 3019 146175
rect 2709 146113 3019 146147
rect 2709 146085 2757 146113
rect 2785 146085 2819 146113
rect 2847 146085 2881 146113
rect 2909 146085 2943 146113
rect 2971 146085 3019 146113
rect 2709 146051 3019 146085
rect 2709 146023 2757 146051
rect 2785 146023 2819 146051
rect 2847 146023 2881 146051
rect 2909 146023 2943 146051
rect 2971 146023 3019 146051
rect 2709 145989 3019 146023
rect 2709 145961 2757 145989
rect 2785 145961 2819 145989
rect 2847 145961 2881 145989
rect 2909 145961 2943 145989
rect 2971 145961 3019 145989
rect 2709 137175 3019 145961
rect 3766 151410 3794 151415
rect 3766 145530 3794 151382
rect 3766 145497 3794 145502
rect 4569 149175 4879 157961
rect 15904 158175 16064 158192
rect 15904 158147 15939 158175
rect 15967 158147 16001 158175
rect 16029 158147 16064 158175
rect 15904 158113 16064 158147
rect 15904 158085 15939 158113
rect 15967 158085 16001 158113
rect 16029 158085 16064 158113
rect 15904 158051 16064 158085
rect 15904 158023 15939 158051
rect 15967 158023 16001 158051
rect 16029 158023 16064 158051
rect 15904 157989 16064 158023
rect 15904 157961 15939 157989
rect 15967 157961 16001 157989
rect 16029 157961 16064 157989
rect 15904 157944 16064 157961
rect 8224 155175 8384 155192
rect 8224 155147 8259 155175
rect 8287 155147 8321 155175
rect 8349 155147 8384 155175
rect 8224 155113 8384 155147
rect 8224 155085 8259 155113
rect 8287 155085 8321 155113
rect 8349 155085 8384 155113
rect 8224 155051 8384 155085
rect 8224 155023 8259 155051
rect 8287 155023 8321 155051
rect 8349 155023 8384 155051
rect 8224 154989 8384 155023
rect 8224 154961 8259 154989
rect 8287 154961 8321 154989
rect 8349 154961 8384 154989
rect 8224 154944 8384 154961
rect 18069 155175 18379 163961
rect 18069 155147 18117 155175
rect 18145 155147 18179 155175
rect 18207 155147 18241 155175
rect 18269 155147 18303 155175
rect 18331 155147 18379 155175
rect 18069 155113 18379 155147
rect 18069 155085 18117 155113
rect 18145 155085 18179 155113
rect 18207 155085 18241 155113
rect 18269 155085 18303 155113
rect 18331 155085 18379 155113
rect 18069 155051 18379 155085
rect 18069 155023 18117 155051
rect 18145 155023 18179 155051
rect 18207 155023 18241 155051
rect 18269 155023 18303 155051
rect 18331 155023 18379 155051
rect 18069 154989 18379 155023
rect 18069 154961 18117 154989
rect 18145 154961 18179 154989
rect 18207 154961 18241 154989
rect 18269 154961 18303 154989
rect 18331 154961 18379 154989
rect 4569 149147 4617 149175
rect 4645 149147 4679 149175
rect 4707 149147 4741 149175
rect 4769 149147 4803 149175
rect 4831 149147 4879 149175
rect 4569 149113 4879 149147
rect 4569 149085 4617 149113
rect 4645 149085 4679 149113
rect 4707 149085 4741 149113
rect 4769 149085 4803 149113
rect 4831 149085 4879 149113
rect 4569 149051 4879 149085
rect 4569 149023 4617 149051
rect 4645 149023 4679 149051
rect 4707 149023 4741 149051
rect 4769 149023 4803 149051
rect 4831 149023 4879 149051
rect 4569 148989 4879 149023
rect 4569 148961 4617 148989
rect 4645 148961 4679 148989
rect 4707 148961 4741 148989
rect 4769 148961 4803 148989
rect 4831 148961 4879 148989
rect 3766 144130 3794 144135
rect 3766 138474 3794 144102
rect 3766 138441 3794 138446
rect 4569 140175 4879 148961
rect 15904 149175 16064 149192
rect 15904 149147 15939 149175
rect 15967 149147 16001 149175
rect 16029 149147 16064 149175
rect 15904 149113 16064 149147
rect 15904 149085 15939 149113
rect 15967 149085 16001 149113
rect 16029 149085 16064 149113
rect 15904 149051 16064 149085
rect 15904 149023 15939 149051
rect 15967 149023 16001 149051
rect 16029 149023 16064 149051
rect 15904 148989 16064 149023
rect 15904 148961 15939 148989
rect 15967 148961 16001 148989
rect 16029 148961 16064 148989
rect 15904 148944 16064 148961
rect 8224 146175 8384 146192
rect 8224 146147 8259 146175
rect 8287 146147 8321 146175
rect 8349 146147 8384 146175
rect 8224 146113 8384 146147
rect 8224 146085 8259 146113
rect 8287 146085 8321 146113
rect 8349 146085 8384 146113
rect 8224 146051 8384 146085
rect 8224 146023 8259 146051
rect 8287 146023 8321 146051
rect 8349 146023 8384 146051
rect 8224 145989 8384 146023
rect 8224 145961 8259 145989
rect 8287 145961 8321 145989
rect 8349 145961 8384 145989
rect 8224 145944 8384 145961
rect 18069 146175 18379 154961
rect 18069 146147 18117 146175
rect 18145 146147 18179 146175
rect 18207 146147 18241 146175
rect 18269 146147 18303 146175
rect 18331 146147 18379 146175
rect 18069 146113 18379 146147
rect 18069 146085 18117 146113
rect 18145 146085 18179 146113
rect 18207 146085 18241 146113
rect 18269 146085 18303 146113
rect 18331 146085 18379 146113
rect 18069 146051 18379 146085
rect 18069 146023 18117 146051
rect 18145 146023 18179 146051
rect 18207 146023 18241 146051
rect 18269 146023 18303 146051
rect 18331 146023 18379 146051
rect 18069 145989 18379 146023
rect 18069 145961 18117 145989
rect 18145 145961 18179 145989
rect 18207 145961 18241 145989
rect 18269 145961 18303 145989
rect 18331 145961 18379 145989
rect 4569 140147 4617 140175
rect 4645 140147 4679 140175
rect 4707 140147 4741 140175
rect 4769 140147 4803 140175
rect 4831 140147 4879 140175
rect 4569 140113 4879 140147
rect 4569 140085 4617 140113
rect 4645 140085 4679 140113
rect 4707 140085 4741 140113
rect 4769 140085 4803 140113
rect 4831 140085 4879 140113
rect 4569 140051 4879 140085
rect 4569 140023 4617 140051
rect 4645 140023 4679 140051
rect 4707 140023 4741 140051
rect 4769 140023 4803 140051
rect 4831 140023 4879 140051
rect 4569 139989 4879 140023
rect 4569 139961 4617 139989
rect 4645 139961 4679 139989
rect 4707 139961 4741 139989
rect 4769 139961 4803 139989
rect 4831 139961 4879 139989
rect 2709 137147 2757 137175
rect 2785 137147 2819 137175
rect 2847 137147 2881 137175
rect 2909 137147 2943 137175
rect 2971 137147 3019 137175
rect 2709 137113 3019 137147
rect 2709 137085 2757 137113
rect 2785 137085 2819 137113
rect 2847 137085 2881 137113
rect 2909 137085 2943 137113
rect 2971 137085 3019 137113
rect 2709 137051 3019 137085
rect 2709 137023 2757 137051
rect 2785 137023 2819 137051
rect 2847 137023 2881 137051
rect 2909 137023 2943 137051
rect 2971 137023 3019 137051
rect 2709 136989 3019 137023
rect 2709 136961 2757 136989
rect 2785 136961 2819 136989
rect 2847 136961 2881 136989
rect 2909 136961 2943 136989
rect 2971 136961 3019 136989
rect 2709 128175 3019 136961
rect 3094 136850 3122 136855
rect 3094 131418 3122 136822
rect 3094 131385 3122 131390
rect 4569 131175 4879 139961
rect 15904 140175 16064 140192
rect 15904 140147 15939 140175
rect 15967 140147 16001 140175
rect 16029 140147 16064 140175
rect 15904 140113 16064 140147
rect 15904 140085 15939 140113
rect 15967 140085 16001 140113
rect 16029 140085 16064 140113
rect 15904 140051 16064 140085
rect 15904 140023 15939 140051
rect 15967 140023 16001 140051
rect 16029 140023 16064 140051
rect 15904 139989 16064 140023
rect 15904 139961 15939 139989
rect 15967 139961 16001 139989
rect 16029 139961 16064 139989
rect 15904 139944 16064 139961
rect 8224 137175 8384 137192
rect 8224 137147 8259 137175
rect 8287 137147 8321 137175
rect 8349 137147 8384 137175
rect 8224 137113 8384 137147
rect 8224 137085 8259 137113
rect 8287 137085 8321 137113
rect 8349 137085 8384 137113
rect 8224 137051 8384 137085
rect 8224 137023 8259 137051
rect 8287 137023 8321 137051
rect 8349 137023 8384 137051
rect 8224 136989 8384 137023
rect 8224 136961 8259 136989
rect 8287 136961 8321 136989
rect 8349 136961 8384 136989
rect 8224 136944 8384 136961
rect 18069 137175 18379 145961
rect 18069 137147 18117 137175
rect 18145 137147 18179 137175
rect 18207 137147 18241 137175
rect 18269 137147 18303 137175
rect 18331 137147 18379 137175
rect 18069 137113 18379 137147
rect 18069 137085 18117 137113
rect 18145 137085 18179 137113
rect 18207 137085 18241 137113
rect 18269 137085 18303 137113
rect 18331 137085 18379 137113
rect 18069 137051 18379 137085
rect 18069 137023 18117 137051
rect 18145 137023 18179 137051
rect 18207 137023 18241 137051
rect 18269 137023 18303 137051
rect 18331 137023 18379 137051
rect 18069 136989 18379 137023
rect 18069 136961 18117 136989
rect 18145 136961 18179 136989
rect 18207 136961 18241 136989
rect 18269 136961 18303 136989
rect 18331 136961 18379 136989
rect 4569 131147 4617 131175
rect 4645 131147 4679 131175
rect 4707 131147 4741 131175
rect 4769 131147 4803 131175
rect 4831 131147 4879 131175
rect 4569 131113 4879 131147
rect 4569 131085 4617 131113
rect 4645 131085 4679 131113
rect 4707 131085 4741 131113
rect 4769 131085 4803 131113
rect 4831 131085 4879 131113
rect 4569 131051 4879 131085
rect 4569 131023 4617 131051
rect 4645 131023 4679 131051
rect 4707 131023 4741 131051
rect 4769 131023 4803 131051
rect 4831 131023 4879 131051
rect 4569 130989 4879 131023
rect 4569 130961 4617 130989
rect 4645 130961 4679 130989
rect 4707 130961 4741 130989
rect 4769 130961 4803 130989
rect 4831 130961 4879 130989
rect 2709 128147 2757 128175
rect 2785 128147 2819 128175
rect 2847 128147 2881 128175
rect 2909 128147 2943 128175
rect 2971 128147 3019 128175
rect 2709 128113 3019 128147
rect 2709 128085 2757 128113
rect 2785 128085 2819 128113
rect 2847 128085 2881 128113
rect 2909 128085 2943 128113
rect 2971 128085 3019 128113
rect 2709 128051 3019 128085
rect 2709 128023 2757 128051
rect 2785 128023 2819 128051
rect 2847 128023 2881 128051
rect 2909 128023 2943 128051
rect 2971 128023 3019 128051
rect 2709 127989 3019 128023
rect 2709 127961 2757 127989
rect 2785 127961 2819 127989
rect 2847 127961 2881 127989
rect 2909 127961 2943 127989
rect 2971 127961 3019 127989
rect 2709 119175 3019 127961
rect 3766 129570 3794 129575
rect 3766 124306 3794 129542
rect 3766 124273 3794 124278
rect 2709 119147 2757 119175
rect 2785 119147 2819 119175
rect 2847 119147 2881 119175
rect 2909 119147 2943 119175
rect 2971 119147 3019 119175
rect 2709 119113 3019 119147
rect 2709 119085 2757 119113
rect 2785 119085 2819 119113
rect 2847 119085 2881 119113
rect 2909 119085 2943 119113
rect 2971 119085 3019 119113
rect 2709 119051 3019 119085
rect 2709 119023 2757 119051
rect 2785 119023 2819 119051
rect 2847 119023 2881 119051
rect 2909 119023 2943 119051
rect 2971 119023 3019 119051
rect 2709 118989 3019 119023
rect 2709 118961 2757 118989
rect 2785 118961 2819 118989
rect 2847 118961 2881 118989
rect 2909 118961 2943 118989
rect 2971 118961 3019 118989
rect 2086 115010 2114 115015
rect 2086 110250 2114 114982
rect 2086 110217 2114 110222
rect -478 110147 -430 110175
rect -402 110147 -368 110175
rect -340 110147 -306 110175
rect -278 110147 -244 110175
rect -216 110147 -168 110175
rect -478 110113 -168 110147
rect -478 110085 -430 110113
rect -402 110085 -368 110113
rect -340 110085 -306 110113
rect -278 110085 -244 110113
rect -216 110085 -168 110113
rect -478 110051 -168 110085
rect -478 110023 -430 110051
rect -402 110023 -368 110051
rect -340 110023 -306 110051
rect -278 110023 -244 110051
rect -216 110023 -168 110051
rect -478 109989 -168 110023
rect -478 109961 -430 109989
rect -402 109961 -368 109989
rect -340 109961 -306 109989
rect -278 109961 -244 109989
rect -216 109961 -168 109989
rect -478 101175 -168 109961
rect -478 101147 -430 101175
rect -402 101147 -368 101175
rect -340 101147 -306 101175
rect -278 101147 -244 101175
rect -216 101147 -168 101175
rect -478 101113 -168 101147
rect -478 101085 -430 101113
rect -402 101085 -368 101113
rect -340 101085 -306 101113
rect -278 101085 -244 101113
rect -216 101085 -168 101113
rect -478 101051 -168 101085
rect -478 101023 -430 101051
rect -402 101023 -368 101051
rect -340 101023 -306 101051
rect -278 101023 -244 101051
rect -216 101023 -168 101051
rect -478 100989 -168 101023
rect -478 100961 -430 100989
rect -402 100961 -368 100989
rect -340 100961 -306 100989
rect -278 100961 -244 100989
rect -216 100961 -168 100989
rect -478 92175 -168 100961
rect 2709 110175 3019 118961
rect 3094 122290 3122 122295
rect 3094 117306 3122 122262
rect 3094 117273 3122 117278
rect 4569 122175 4879 130961
rect 15904 131175 16064 131192
rect 15904 131147 15939 131175
rect 15967 131147 16001 131175
rect 16029 131147 16064 131175
rect 15904 131113 16064 131147
rect 15904 131085 15939 131113
rect 15967 131085 16001 131113
rect 16029 131085 16064 131113
rect 15904 131051 16064 131085
rect 15904 131023 15939 131051
rect 15967 131023 16001 131051
rect 16029 131023 16064 131051
rect 15904 130989 16064 131023
rect 15904 130961 15939 130989
rect 15967 130961 16001 130989
rect 16029 130961 16064 130989
rect 15904 130944 16064 130961
rect 8224 128175 8384 128192
rect 8224 128147 8259 128175
rect 8287 128147 8321 128175
rect 8349 128147 8384 128175
rect 8224 128113 8384 128147
rect 8224 128085 8259 128113
rect 8287 128085 8321 128113
rect 8349 128085 8384 128113
rect 8224 128051 8384 128085
rect 8224 128023 8259 128051
rect 8287 128023 8321 128051
rect 8349 128023 8384 128051
rect 8224 127989 8384 128023
rect 8224 127961 8259 127989
rect 8287 127961 8321 127989
rect 8349 127961 8384 127989
rect 8224 127944 8384 127961
rect 18069 128175 18379 136961
rect 18069 128147 18117 128175
rect 18145 128147 18179 128175
rect 18207 128147 18241 128175
rect 18269 128147 18303 128175
rect 18331 128147 18379 128175
rect 18069 128113 18379 128147
rect 18069 128085 18117 128113
rect 18145 128085 18179 128113
rect 18207 128085 18241 128113
rect 18269 128085 18303 128113
rect 18331 128085 18379 128113
rect 18069 128051 18379 128085
rect 18069 128023 18117 128051
rect 18145 128023 18179 128051
rect 18207 128023 18241 128051
rect 18269 128023 18303 128051
rect 18331 128023 18379 128051
rect 18069 127989 18379 128023
rect 18069 127961 18117 127989
rect 18145 127961 18179 127989
rect 18207 127961 18241 127989
rect 18269 127961 18303 127989
rect 18331 127961 18379 127989
rect 4569 122147 4617 122175
rect 4645 122147 4679 122175
rect 4707 122147 4741 122175
rect 4769 122147 4803 122175
rect 4831 122147 4879 122175
rect 4569 122113 4879 122147
rect 4569 122085 4617 122113
rect 4645 122085 4679 122113
rect 4707 122085 4741 122113
rect 4769 122085 4803 122113
rect 4831 122085 4879 122113
rect 4569 122051 4879 122085
rect 4569 122023 4617 122051
rect 4645 122023 4679 122051
rect 4707 122023 4741 122051
rect 4769 122023 4803 122051
rect 4831 122023 4879 122051
rect 4569 121989 4879 122023
rect 4569 121961 4617 121989
rect 4645 121961 4679 121989
rect 4707 121961 4741 121989
rect 4769 121961 4803 121989
rect 4831 121961 4879 121989
rect 2709 110147 2757 110175
rect 2785 110147 2819 110175
rect 2847 110147 2881 110175
rect 2909 110147 2943 110175
rect 2971 110147 3019 110175
rect 2709 110113 3019 110147
rect 2709 110085 2757 110113
rect 2785 110085 2819 110113
rect 2847 110085 2881 110113
rect 2909 110085 2943 110113
rect 2971 110085 3019 110113
rect 2709 110051 3019 110085
rect 2709 110023 2757 110051
rect 2785 110023 2819 110051
rect 2847 110023 2881 110051
rect 2909 110023 2943 110051
rect 2971 110023 3019 110051
rect 2709 109989 3019 110023
rect 2709 109961 2757 109989
rect 2785 109961 2819 109989
rect 2847 109961 2881 109989
rect 2909 109961 2943 109989
rect 2971 109961 3019 109989
rect 2709 101175 3019 109961
rect 4569 113175 4879 121961
rect 15904 122175 16064 122192
rect 15904 122147 15939 122175
rect 15967 122147 16001 122175
rect 16029 122147 16064 122175
rect 15904 122113 16064 122147
rect 15904 122085 15939 122113
rect 15967 122085 16001 122113
rect 16029 122085 16064 122113
rect 15904 122051 16064 122085
rect 15904 122023 15939 122051
rect 15967 122023 16001 122051
rect 16029 122023 16064 122051
rect 15904 121989 16064 122023
rect 15904 121961 15939 121989
rect 15967 121961 16001 121989
rect 16029 121961 16064 121989
rect 15904 121944 16064 121961
rect 8224 119175 8384 119192
rect 8224 119147 8259 119175
rect 8287 119147 8321 119175
rect 8349 119147 8384 119175
rect 8224 119113 8384 119147
rect 8224 119085 8259 119113
rect 8287 119085 8321 119113
rect 8349 119085 8384 119113
rect 8224 119051 8384 119085
rect 8224 119023 8259 119051
rect 8287 119023 8321 119051
rect 8349 119023 8384 119051
rect 8224 118989 8384 119023
rect 8224 118961 8259 118989
rect 8287 118961 8321 118989
rect 8349 118961 8384 118989
rect 8224 118944 8384 118961
rect 18069 119175 18379 127961
rect 18069 119147 18117 119175
rect 18145 119147 18179 119175
rect 18207 119147 18241 119175
rect 18269 119147 18303 119175
rect 18331 119147 18379 119175
rect 18069 119113 18379 119147
rect 18069 119085 18117 119113
rect 18145 119085 18179 119113
rect 18207 119085 18241 119113
rect 18269 119085 18303 119113
rect 18331 119085 18379 119113
rect 18069 119051 18379 119085
rect 18069 119023 18117 119051
rect 18145 119023 18179 119051
rect 18207 119023 18241 119051
rect 18269 119023 18303 119051
rect 18331 119023 18379 119051
rect 18069 118989 18379 119023
rect 18069 118961 18117 118989
rect 18145 118961 18179 118989
rect 18207 118961 18241 118989
rect 18269 118961 18303 118989
rect 18331 118961 18379 118989
rect 4569 113147 4617 113175
rect 4645 113147 4679 113175
rect 4707 113147 4741 113175
rect 4769 113147 4803 113175
rect 4831 113147 4879 113175
rect 4569 113113 4879 113147
rect 4569 113085 4617 113113
rect 4645 113085 4679 113113
rect 4707 113085 4741 113113
rect 4769 113085 4803 113113
rect 4831 113085 4879 113113
rect 4569 113051 4879 113085
rect 4569 113023 4617 113051
rect 4645 113023 4679 113051
rect 4707 113023 4741 113051
rect 4769 113023 4803 113051
rect 4831 113023 4879 113051
rect 4569 112989 4879 113023
rect 4569 112961 4617 112989
rect 4645 112961 4679 112989
rect 4707 112961 4741 112989
rect 4769 112961 4803 112989
rect 4831 112961 4879 112989
rect 3094 107730 3122 107735
rect 3094 103194 3122 107702
rect 3094 103161 3122 103166
rect 4569 104175 4879 112961
rect 15904 113175 16064 113192
rect 15904 113147 15939 113175
rect 15967 113147 16001 113175
rect 16029 113147 16064 113175
rect 15904 113113 16064 113147
rect 15904 113085 15939 113113
rect 15967 113085 16001 113113
rect 16029 113085 16064 113113
rect 15904 113051 16064 113085
rect 15904 113023 15939 113051
rect 15967 113023 16001 113051
rect 16029 113023 16064 113051
rect 15904 112989 16064 113023
rect 15904 112961 15939 112989
rect 15967 112961 16001 112989
rect 16029 112961 16064 112989
rect 15904 112944 16064 112961
rect 8224 110175 8384 110192
rect 8224 110147 8259 110175
rect 8287 110147 8321 110175
rect 8349 110147 8384 110175
rect 8224 110113 8384 110147
rect 8224 110085 8259 110113
rect 8287 110085 8321 110113
rect 8349 110085 8384 110113
rect 8224 110051 8384 110085
rect 8224 110023 8259 110051
rect 8287 110023 8321 110051
rect 8349 110023 8384 110051
rect 8224 109989 8384 110023
rect 8224 109961 8259 109989
rect 8287 109961 8321 109989
rect 8349 109961 8384 109989
rect 8224 109944 8384 109961
rect 18069 110175 18379 118961
rect 18069 110147 18117 110175
rect 18145 110147 18179 110175
rect 18207 110147 18241 110175
rect 18269 110147 18303 110175
rect 18331 110147 18379 110175
rect 18069 110113 18379 110147
rect 18069 110085 18117 110113
rect 18145 110085 18179 110113
rect 18207 110085 18241 110113
rect 18269 110085 18303 110113
rect 18331 110085 18379 110113
rect 18069 110051 18379 110085
rect 18069 110023 18117 110051
rect 18145 110023 18179 110051
rect 18207 110023 18241 110051
rect 18269 110023 18303 110051
rect 18331 110023 18379 110051
rect 18069 109989 18379 110023
rect 18069 109961 18117 109989
rect 18145 109961 18179 109989
rect 18207 109961 18241 109989
rect 18269 109961 18303 109989
rect 18331 109961 18379 109989
rect 4569 104147 4617 104175
rect 4645 104147 4679 104175
rect 4707 104147 4741 104175
rect 4769 104147 4803 104175
rect 4831 104147 4879 104175
rect 4569 104113 4879 104147
rect 4569 104085 4617 104113
rect 4645 104085 4679 104113
rect 4707 104085 4741 104113
rect 4769 104085 4803 104113
rect 4831 104085 4879 104113
rect 4569 104051 4879 104085
rect 4569 104023 4617 104051
rect 4645 104023 4679 104051
rect 4707 104023 4741 104051
rect 4769 104023 4803 104051
rect 4831 104023 4879 104051
rect 4569 103989 4879 104023
rect 4569 103961 4617 103989
rect 4645 103961 4679 103989
rect 4707 103961 4741 103989
rect 4769 103961 4803 103989
rect 4831 103961 4879 103989
rect 2709 101147 2757 101175
rect 2785 101147 2819 101175
rect 2847 101147 2881 101175
rect 2909 101147 2943 101175
rect 2971 101147 3019 101175
rect 2709 101113 3019 101147
rect 2709 101085 2757 101113
rect 2785 101085 2819 101113
rect 2847 101085 2881 101113
rect 2909 101085 2943 101113
rect 2971 101085 3019 101113
rect 2709 101051 3019 101085
rect 2709 101023 2757 101051
rect 2785 101023 2819 101051
rect 2847 101023 2881 101051
rect 2909 101023 2943 101051
rect 2971 101023 3019 101051
rect 2709 100989 3019 101023
rect 2709 100961 2757 100989
rect 2785 100961 2819 100989
rect 2847 100961 2881 100989
rect 2909 100961 2943 100989
rect 2971 100961 3019 100989
rect 2086 100450 2114 100455
rect 2086 96138 2114 100422
rect 2086 96105 2114 96110
rect -478 92147 -430 92175
rect -402 92147 -368 92175
rect -340 92147 -306 92175
rect -278 92147 -244 92175
rect -216 92147 -168 92175
rect -478 92113 -168 92147
rect -478 92085 -430 92113
rect -402 92085 -368 92113
rect -340 92085 -306 92113
rect -278 92085 -244 92113
rect -216 92085 -168 92113
rect -478 92051 -168 92085
rect -478 92023 -430 92051
rect -402 92023 -368 92051
rect -340 92023 -306 92051
rect -278 92023 -244 92051
rect -216 92023 -168 92051
rect -478 91989 -168 92023
rect -478 91961 -430 91989
rect -402 91961 -368 91989
rect -340 91961 -306 91989
rect -278 91961 -244 91989
rect -216 91961 -168 91989
rect -478 83175 -168 91961
rect 2478 93170 2506 93175
rect 2478 89026 2506 93142
rect 2478 88993 2506 88998
rect 2709 92175 3019 100961
rect 2709 92147 2757 92175
rect 2785 92147 2819 92175
rect 2847 92147 2881 92175
rect 2909 92147 2943 92175
rect 2971 92147 3019 92175
rect 2709 92113 3019 92147
rect 2709 92085 2757 92113
rect 2785 92085 2819 92113
rect 2847 92085 2881 92113
rect 2909 92085 2943 92113
rect 2971 92085 3019 92113
rect 2709 92051 3019 92085
rect 2709 92023 2757 92051
rect 2785 92023 2819 92051
rect 2847 92023 2881 92051
rect 2909 92023 2943 92051
rect 2971 92023 3019 92051
rect 2709 91989 3019 92023
rect 2709 91961 2757 91989
rect 2785 91961 2819 91989
rect 2847 91961 2881 91989
rect 2909 91961 2943 91989
rect 2971 91961 3019 91989
rect -478 83147 -430 83175
rect -402 83147 -368 83175
rect -340 83147 -306 83175
rect -278 83147 -244 83175
rect -216 83147 -168 83175
rect -478 83113 -168 83147
rect -478 83085 -430 83113
rect -402 83085 -368 83113
rect -340 83085 -306 83113
rect -278 83085 -244 83113
rect -216 83085 -168 83113
rect -478 83051 -168 83085
rect -478 83023 -430 83051
rect -402 83023 -368 83051
rect -340 83023 -306 83051
rect -278 83023 -244 83051
rect -216 83023 -168 83051
rect -478 82989 -168 83023
rect -478 82961 -430 82989
rect -402 82961 -368 82989
rect -340 82961 -306 82989
rect -278 82961 -244 82989
rect -216 82961 -168 82989
rect -478 74175 -168 82961
rect 2086 85890 2114 85895
rect 2086 82026 2114 85862
rect 2086 81993 2114 81998
rect 2709 83175 3019 91961
rect 2709 83147 2757 83175
rect 2785 83147 2819 83175
rect 2847 83147 2881 83175
rect 2909 83147 2943 83175
rect 2971 83147 3019 83175
rect 2709 83113 3019 83147
rect 2709 83085 2757 83113
rect 2785 83085 2819 83113
rect 2847 83085 2881 83113
rect 2909 83085 2943 83113
rect 2971 83085 3019 83113
rect 2709 83051 3019 83085
rect 2709 83023 2757 83051
rect 2785 83023 2819 83051
rect 2847 83023 2881 83051
rect 2909 83023 2943 83051
rect 2971 83023 3019 83051
rect 2709 82989 3019 83023
rect 2709 82961 2757 82989
rect 2785 82961 2819 82989
rect 2847 82961 2881 82989
rect 2909 82961 2943 82989
rect 2971 82961 3019 82989
rect -478 74147 -430 74175
rect -402 74147 -368 74175
rect -340 74147 -306 74175
rect -278 74147 -244 74175
rect -216 74147 -168 74175
rect -478 74113 -168 74147
rect -478 74085 -430 74113
rect -402 74085 -368 74113
rect -340 74085 -306 74113
rect -278 74085 -244 74113
rect -216 74085 -168 74113
rect -478 74051 -168 74085
rect -478 74023 -430 74051
rect -402 74023 -368 74051
rect -340 74023 -306 74051
rect -278 74023 -244 74051
rect -216 74023 -168 74051
rect -478 73989 -168 74023
rect -478 73961 -430 73989
rect -402 73961 -368 73989
rect -340 73961 -306 73989
rect -278 73961 -244 73989
rect -216 73961 -168 73989
rect -478 65175 -168 73961
rect -478 65147 -430 65175
rect -402 65147 -368 65175
rect -340 65147 -306 65175
rect -278 65147 -244 65175
rect -216 65147 -168 65175
rect -478 65113 -168 65147
rect -478 65085 -430 65113
rect -402 65085 -368 65113
rect -340 65085 -306 65113
rect -278 65085 -244 65113
rect -216 65085 -168 65113
rect -478 65051 -168 65085
rect -478 65023 -430 65051
rect -402 65023 -368 65051
rect -340 65023 -306 65051
rect -278 65023 -244 65051
rect -216 65023 -168 65051
rect -478 64989 -168 65023
rect -478 64961 -430 64989
rect -402 64961 -368 64989
rect -340 64961 -306 64989
rect -278 64961 -244 64989
rect -216 64961 -168 64989
rect -478 56175 -168 64961
rect -478 56147 -430 56175
rect -402 56147 -368 56175
rect -340 56147 -306 56175
rect -278 56147 -244 56175
rect -216 56147 -168 56175
rect -478 56113 -168 56147
rect -478 56085 -430 56113
rect -402 56085 -368 56113
rect -340 56085 -306 56113
rect -278 56085 -244 56113
rect -216 56085 -168 56113
rect -478 56051 -168 56085
rect -478 56023 -430 56051
rect -402 56023 -368 56051
rect -340 56023 -306 56051
rect -278 56023 -244 56051
rect -216 56023 -168 56051
rect -478 55989 -168 56023
rect -478 55961 -430 55989
rect -402 55961 -368 55989
rect -340 55961 -306 55989
rect -278 55961 -244 55989
rect -216 55961 -168 55989
rect -478 47175 -168 55961
rect -478 47147 -430 47175
rect -402 47147 -368 47175
rect -340 47147 -306 47175
rect -278 47147 -244 47175
rect -216 47147 -168 47175
rect -478 47113 -168 47147
rect -478 47085 -430 47113
rect -402 47085 -368 47113
rect -340 47085 -306 47113
rect -278 47085 -244 47113
rect -216 47085 -168 47113
rect -478 47051 -168 47085
rect -478 47023 -430 47051
rect -402 47023 -368 47051
rect -340 47023 -306 47051
rect -278 47023 -244 47051
rect -216 47023 -168 47051
rect -478 46989 -168 47023
rect -478 46961 -430 46989
rect -402 46961 -368 46989
rect -340 46961 -306 46989
rect -278 46961 -244 46989
rect -216 46961 -168 46989
rect -478 38175 -168 46961
rect -478 38147 -430 38175
rect -402 38147 -368 38175
rect -340 38147 -306 38175
rect -278 38147 -244 38175
rect -216 38147 -168 38175
rect -478 38113 -168 38147
rect -478 38085 -430 38113
rect -402 38085 -368 38113
rect -340 38085 -306 38113
rect -278 38085 -244 38113
rect -216 38085 -168 38113
rect -478 38051 -168 38085
rect -478 38023 -430 38051
rect -402 38023 -368 38051
rect -340 38023 -306 38051
rect -278 38023 -244 38051
rect -216 38023 -168 38051
rect -478 37989 -168 38023
rect -478 37961 -430 37989
rect -402 37961 -368 37989
rect -340 37961 -306 37989
rect -278 37961 -244 37989
rect -216 37961 -168 37989
rect -478 29175 -168 37961
rect -478 29147 -430 29175
rect -402 29147 -368 29175
rect -340 29147 -306 29175
rect -278 29147 -244 29175
rect -216 29147 -168 29175
rect -478 29113 -168 29147
rect -478 29085 -430 29113
rect -402 29085 -368 29113
rect -340 29085 -306 29113
rect -278 29085 -244 29113
rect -216 29085 -168 29113
rect -478 29051 -168 29085
rect -478 29023 -430 29051
rect -402 29023 -368 29051
rect -340 29023 -306 29051
rect -278 29023 -244 29051
rect -216 29023 -168 29051
rect -478 28989 -168 29023
rect -478 28961 -430 28989
rect -402 28961 -368 28989
rect -340 28961 -306 28989
rect -278 28961 -244 28989
rect -216 28961 -168 28989
rect -478 20175 -168 28961
rect 2709 74175 3019 82961
rect 4569 95175 4879 103961
rect 15904 104175 16064 104192
rect 15904 104147 15939 104175
rect 15967 104147 16001 104175
rect 16029 104147 16064 104175
rect 15904 104113 16064 104147
rect 15904 104085 15939 104113
rect 15967 104085 16001 104113
rect 16029 104085 16064 104113
rect 15904 104051 16064 104085
rect 15904 104023 15939 104051
rect 15967 104023 16001 104051
rect 16029 104023 16064 104051
rect 15904 103989 16064 104023
rect 15904 103961 15939 103989
rect 15967 103961 16001 103989
rect 16029 103961 16064 103989
rect 15904 103944 16064 103961
rect 8224 101175 8384 101192
rect 8224 101147 8259 101175
rect 8287 101147 8321 101175
rect 8349 101147 8384 101175
rect 8224 101113 8384 101147
rect 8224 101085 8259 101113
rect 8287 101085 8321 101113
rect 8349 101085 8384 101113
rect 8224 101051 8384 101085
rect 8224 101023 8259 101051
rect 8287 101023 8321 101051
rect 8349 101023 8384 101051
rect 8224 100989 8384 101023
rect 8224 100961 8259 100989
rect 8287 100961 8321 100989
rect 8349 100961 8384 100989
rect 8224 100944 8384 100961
rect 18069 101175 18379 109961
rect 18069 101147 18117 101175
rect 18145 101147 18179 101175
rect 18207 101147 18241 101175
rect 18269 101147 18303 101175
rect 18331 101147 18379 101175
rect 18069 101113 18379 101147
rect 18069 101085 18117 101113
rect 18145 101085 18179 101113
rect 18207 101085 18241 101113
rect 18269 101085 18303 101113
rect 18331 101085 18379 101113
rect 18069 101051 18379 101085
rect 18069 101023 18117 101051
rect 18145 101023 18179 101051
rect 18207 101023 18241 101051
rect 18269 101023 18303 101051
rect 18331 101023 18379 101051
rect 18069 100989 18379 101023
rect 18069 100961 18117 100989
rect 18145 100961 18179 100989
rect 18207 100961 18241 100989
rect 18269 100961 18303 100989
rect 18331 100961 18379 100989
rect 4569 95147 4617 95175
rect 4645 95147 4679 95175
rect 4707 95147 4741 95175
rect 4769 95147 4803 95175
rect 4831 95147 4879 95175
rect 4569 95113 4879 95147
rect 4569 95085 4617 95113
rect 4645 95085 4679 95113
rect 4707 95085 4741 95113
rect 4769 95085 4803 95113
rect 4831 95085 4879 95113
rect 4569 95051 4879 95085
rect 4569 95023 4617 95051
rect 4645 95023 4679 95051
rect 4707 95023 4741 95051
rect 4769 95023 4803 95051
rect 4831 95023 4879 95051
rect 4569 94989 4879 95023
rect 4569 94961 4617 94989
rect 4645 94961 4679 94989
rect 4707 94961 4741 94989
rect 4769 94961 4803 94989
rect 4831 94961 4879 94989
rect 4569 86175 4879 94961
rect 15904 95175 16064 95192
rect 15904 95147 15939 95175
rect 15967 95147 16001 95175
rect 16029 95147 16064 95175
rect 15904 95113 16064 95147
rect 15904 95085 15939 95113
rect 15967 95085 16001 95113
rect 16029 95085 16064 95113
rect 15904 95051 16064 95085
rect 15904 95023 15939 95051
rect 15967 95023 16001 95051
rect 16029 95023 16064 95051
rect 15904 94989 16064 95023
rect 15904 94961 15939 94989
rect 15967 94961 16001 94989
rect 16029 94961 16064 94989
rect 15904 94944 16064 94961
rect 8224 92175 8384 92192
rect 8224 92147 8259 92175
rect 8287 92147 8321 92175
rect 8349 92147 8384 92175
rect 8224 92113 8384 92147
rect 8224 92085 8259 92113
rect 8287 92085 8321 92113
rect 8349 92085 8384 92113
rect 8224 92051 8384 92085
rect 8224 92023 8259 92051
rect 8287 92023 8321 92051
rect 8349 92023 8384 92051
rect 8224 91989 8384 92023
rect 8224 91961 8259 91989
rect 8287 91961 8321 91989
rect 8349 91961 8384 91989
rect 8224 91944 8384 91961
rect 18069 92175 18379 100961
rect 18069 92147 18117 92175
rect 18145 92147 18179 92175
rect 18207 92147 18241 92175
rect 18269 92147 18303 92175
rect 18331 92147 18379 92175
rect 18069 92113 18379 92147
rect 18069 92085 18117 92113
rect 18145 92085 18179 92113
rect 18207 92085 18241 92113
rect 18269 92085 18303 92113
rect 18331 92085 18379 92113
rect 18069 92051 18379 92085
rect 18069 92023 18117 92051
rect 18145 92023 18179 92051
rect 18207 92023 18241 92051
rect 18269 92023 18303 92051
rect 18331 92023 18379 92051
rect 18069 91989 18379 92023
rect 18069 91961 18117 91989
rect 18145 91961 18179 91989
rect 18207 91961 18241 91989
rect 18269 91961 18303 91989
rect 18331 91961 18379 91989
rect 4569 86147 4617 86175
rect 4645 86147 4679 86175
rect 4707 86147 4741 86175
rect 4769 86147 4803 86175
rect 4831 86147 4879 86175
rect 4569 86113 4879 86147
rect 4569 86085 4617 86113
rect 4645 86085 4679 86113
rect 4707 86085 4741 86113
rect 4769 86085 4803 86113
rect 4831 86085 4879 86113
rect 4569 86051 4879 86085
rect 4569 86023 4617 86051
rect 4645 86023 4679 86051
rect 4707 86023 4741 86051
rect 4769 86023 4803 86051
rect 4831 86023 4879 86051
rect 4569 85989 4879 86023
rect 4569 85961 4617 85989
rect 4645 85961 4679 85989
rect 4707 85961 4741 85989
rect 4769 85961 4803 85989
rect 4831 85961 4879 85989
rect 3766 78610 3794 78615
rect 3766 74970 3794 78582
rect 3766 74937 3794 74942
rect 4569 77175 4879 85961
rect 15904 86175 16064 86192
rect 15904 86147 15939 86175
rect 15967 86147 16001 86175
rect 16029 86147 16064 86175
rect 15904 86113 16064 86147
rect 15904 86085 15939 86113
rect 15967 86085 16001 86113
rect 16029 86085 16064 86113
rect 15904 86051 16064 86085
rect 15904 86023 15939 86051
rect 15967 86023 16001 86051
rect 16029 86023 16064 86051
rect 15904 85989 16064 86023
rect 15904 85961 15939 85989
rect 15967 85961 16001 85989
rect 16029 85961 16064 85989
rect 15904 85944 16064 85961
rect 8224 83175 8384 83192
rect 8224 83147 8259 83175
rect 8287 83147 8321 83175
rect 8349 83147 8384 83175
rect 8224 83113 8384 83147
rect 8224 83085 8259 83113
rect 8287 83085 8321 83113
rect 8349 83085 8384 83113
rect 8224 83051 8384 83085
rect 8224 83023 8259 83051
rect 8287 83023 8321 83051
rect 8349 83023 8384 83051
rect 8224 82989 8384 83023
rect 8224 82961 8259 82989
rect 8287 82961 8321 82989
rect 8349 82961 8384 82989
rect 8224 82944 8384 82961
rect 18069 83175 18379 91961
rect 18069 83147 18117 83175
rect 18145 83147 18179 83175
rect 18207 83147 18241 83175
rect 18269 83147 18303 83175
rect 18331 83147 18379 83175
rect 18069 83113 18379 83147
rect 18069 83085 18117 83113
rect 18145 83085 18179 83113
rect 18207 83085 18241 83113
rect 18269 83085 18303 83113
rect 18331 83085 18379 83113
rect 18069 83051 18379 83085
rect 18069 83023 18117 83051
rect 18145 83023 18179 83051
rect 18207 83023 18241 83051
rect 18269 83023 18303 83051
rect 18331 83023 18379 83051
rect 18069 82989 18379 83023
rect 18069 82961 18117 82989
rect 18145 82961 18179 82989
rect 18207 82961 18241 82989
rect 18269 82961 18303 82989
rect 18331 82961 18379 82989
rect 4569 77147 4617 77175
rect 4645 77147 4679 77175
rect 4707 77147 4741 77175
rect 4769 77147 4803 77175
rect 4831 77147 4879 77175
rect 4569 77113 4879 77147
rect 4569 77085 4617 77113
rect 4645 77085 4679 77113
rect 4707 77085 4741 77113
rect 4769 77085 4803 77113
rect 4831 77085 4879 77113
rect 4569 77051 4879 77085
rect 4569 77023 4617 77051
rect 4645 77023 4679 77051
rect 4707 77023 4741 77051
rect 4769 77023 4803 77051
rect 4831 77023 4879 77051
rect 4569 76989 4879 77023
rect 4569 76961 4617 76989
rect 4645 76961 4679 76989
rect 4707 76961 4741 76989
rect 4769 76961 4803 76989
rect 4831 76961 4879 76989
rect 2709 74147 2757 74175
rect 2785 74147 2819 74175
rect 2847 74147 2881 74175
rect 2909 74147 2943 74175
rect 2971 74147 3019 74175
rect 2709 74113 3019 74147
rect 2709 74085 2757 74113
rect 2785 74085 2819 74113
rect 2847 74085 2881 74113
rect 2909 74085 2943 74113
rect 2971 74085 3019 74113
rect 2709 74051 3019 74085
rect 2709 74023 2757 74051
rect 2785 74023 2819 74051
rect 2847 74023 2881 74051
rect 2909 74023 2943 74051
rect 2971 74023 3019 74051
rect 2709 73989 3019 74023
rect 2709 73961 2757 73989
rect 2785 73961 2819 73989
rect 2847 73961 2881 73989
rect 2909 73961 2943 73989
rect 2971 73961 3019 73989
rect 2709 65175 3019 73961
rect 3766 71330 3794 71335
rect 3766 67914 3794 71302
rect 3766 67881 3794 67886
rect 4569 68175 4879 76961
rect 15904 77175 16064 77192
rect 15904 77147 15939 77175
rect 15967 77147 16001 77175
rect 16029 77147 16064 77175
rect 15904 77113 16064 77147
rect 15904 77085 15939 77113
rect 15967 77085 16001 77113
rect 16029 77085 16064 77113
rect 15904 77051 16064 77085
rect 15904 77023 15939 77051
rect 15967 77023 16001 77051
rect 16029 77023 16064 77051
rect 15904 76989 16064 77023
rect 15904 76961 15939 76989
rect 15967 76961 16001 76989
rect 16029 76961 16064 76989
rect 15904 76944 16064 76961
rect 8224 74175 8384 74192
rect 8224 74147 8259 74175
rect 8287 74147 8321 74175
rect 8349 74147 8384 74175
rect 8224 74113 8384 74147
rect 8224 74085 8259 74113
rect 8287 74085 8321 74113
rect 8349 74085 8384 74113
rect 8224 74051 8384 74085
rect 8224 74023 8259 74051
rect 8287 74023 8321 74051
rect 8349 74023 8384 74051
rect 8224 73989 8384 74023
rect 8224 73961 8259 73989
rect 8287 73961 8321 73989
rect 8349 73961 8384 73989
rect 8224 73944 8384 73961
rect 18069 74175 18379 82961
rect 18069 74147 18117 74175
rect 18145 74147 18179 74175
rect 18207 74147 18241 74175
rect 18269 74147 18303 74175
rect 18331 74147 18379 74175
rect 18069 74113 18379 74147
rect 18069 74085 18117 74113
rect 18145 74085 18179 74113
rect 18207 74085 18241 74113
rect 18269 74085 18303 74113
rect 18331 74085 18379 74113
rect 18069 74051 18379 74085
rect 18069 74023 18117 74051
rect 18145 74023 18179 74051
rect 18207 74023 18241 74051
rect 18269 74023 18303 74051
rect 18331 74023 18379 74051
rect 18069 73989 18379 74023
rect 18069 73961 18117 73989
rect 18145 73961 18179 73989
rect 18207 73961 18241 73989
rect 18269 73961 18303 73989
rect 18331 73961 18379 73989
rect 4569 68147 4617 68175
rect 4645 68147 4679 68175
rect 4707 68147 4741 68175
rect 4769 68147 4803 68175
rect 4831 68147 4879 68175
rect 4569 68113 4879 68147
rect 4569 68085 4617 68113
rect 4645 68085 4679 68113
rect 4707 68085 4741 68113
rect 4769 68085 4803 68113
rect 4831 68085 4879 68113
rect 4569 68051 4879 68085
rect 4569 68023 4617 68051
rect 4645 68023 4679 68051
rect 4707 68023 4741 68051
rect 4769 68023 4803 68051
rect 4831 68023 4879 68051
rect 4569 67989 4879 68023
rect 4569 67961 4617 67989
rect 4645 67961 4679 67989
rect 4707 67961 4741 67989
rect 4769 67961 4803 67989
rect 4831 67961 4879 67989
rect 2709 65147 2757 65175
rect 2785 65147 2819 65175
rect 2847 65147 2881 65175
rect 2909 65147 2943 65175
rect 2971 65147 3019 65175
rect 2709 65113 3019 65147
rect 2709 65085 2757 65113
rect 2785 65085 2819 65113
rect 2847 65085 2881 65113
rect 2909 65085 2943 65113
rect 2971 65085 3019 65113
rect 2709 65051 3019 65085
rect 2709 65023 2757 65051
rect 2785 65023 2819 65051
rect 2847 65023 2881 65051
rect 2909 65023 2943 65051
rect 2971 65023 3019 65051
rect 2709 64989 3019 65023
rect 2709 64961 2757 64989
rect 2785 64961 2819 64989
rect 2847 64961 2881 64989
rect 2909 64961 2943 64989
rect 2971 64961 3019 64989
rect 2709 56175 3019 64961
rect 3374 64050 3402 64055
rect 3374 60858 3402 64022
rect 3374 60825 3402 60830
rect 4569 59175 4879 67961
rect 15904 68175 16064 68192
rect 15904 68147 15939 68175
rect 15967 68147 16001 68175
rect 16029 68147 16064 68175
rect 15904 68113 16064 68147
rect 15904 68085 15939 68113
rect 15967 68085 16001 68113
rect 16029 68085 16064 68113
rect 15904 68051 16064 68085
rect 15904 68023 15939 68051
rect 15967 68023 16001 68051
rect 16029 68023 16064 68051
rect 15904 67989 16064 68023
rect 15904 67961 15939 67989
rect 15967 67961 16001 67989
rect 16029 67961 16064 67989
rect 15904 67944 16064 67961
rect 8224 65175 8384 65192
rect 8224 65147 8259 65175
rect 8287 65147 8321 65175
rect 8349 65147 8384 65175
rect 8224 65113 8384 65147
rect 8224 65085 8259 65113
rect 8287 65085 8321 65113
rect 8349 65085 8384 65113
rect 8224 65051 8384 65085
rect 8224 65023 8259 65051
rect 8287 65023 8321 65051
rect 8349 65023 8384 65051
rect 8224 64989 8384 65023
rect 8224 64961 8259 64989
rect 8287 64961 8321 64989
rect 8349 64961 8384 64989
rect 8224 64944 8384 64961
rect 18069 65175 18379 73961
rect 18069 65147 18117 65175
rect 18145 65147 18179 65175
rect 18207 65147 18241 65175
rect 18269 65147 18303 65175
rect 18331 65147 18379 65175
rect 18069 65113 18379 65147
rect 18069 65085 18117 65113
rect 18145 65085 18179 65113
rect 18207 65085 18241 65113
rect 18269 65085 18303 65113
rect 18331 65085 18379 65113
rect 18069 65051 18379 65085
rect 18069 65023 18117 65051
rect 18145 65023 18179 65051
rect 18207 65023 18241 65051
rect 18269 65023 18303 65051
rect 18331 65023 18379 65051
rect 18069 64989 18379 65023
rect 18069 64961 18117 64989
rect 18145 64961 18179 64989
rect 18207 64961 18241 64989
rect 18269 64961 18303 64989
rect 18331 64961 18379 64989
rect 4569 59147 4617 59175
rect 4645 59147 4679 59175
rect 4707 59147 4741 59175
rect 4769 59147 4803 59175
rect 4831 59147 4879 59175
rect 4569 59113 4879 59147
rect 4569 59085 4617 59113
rect 4645 59085 4679 59113
rect 4707 59085 4741 59113
rect 4769 59085 4803 59113
rect 4831 59085 4879 59113
rect 4569 59051 4879 59085
rect 4569 59023 4617 59051
rect 4645 59023 4679 59051
rect 4707 59023 4741 59051
rect 4769 59023 4803 59051
rect 4831 59023 4879 59051
rect 4569 58989 4879 59023
rect 4569 58961 4617 58989
rect 4645 58961 4679 58989
rect 4707 58961 4741 58989
rect 4769 58961 4803 58989
rect 4831 58961 4879 58989
rect 2709 56147 2757 56175
rect 2785 56147 2819 56175
rect 2847 56147 2881 56175
rect 2909 56147 2943 56175
rect 2971 56147 3019 56175
rect 2709 56113 3019 56147
rect 2709 56085 2757 56113
rect 2785 56085 2819 56113
rect 2847 56085 2881 56113
rect 2909 56085 2943 56113
rect 2971 56085 3019 56113
rect 2709 56051 3019 56085
rect 2709 56023 2757 56051
rect 2785 56023 2819 56051
rect 2847 56023 2881 56051
rect 2909 56023 2943 56051
rect 2971 56023 3019 56051
rect 2709 55989 3019 56023
rect 2709 55961 2757 55989
rect 2785 55961 2819 55989
rect 2847 55961 2881 55989
rect 2909 55961 2943 55989
rect 2971 55961 3019 55989
rect 2709 47175 3019 55961
rect 3374 56770 3402 56775
rect 3374 53746 3402 56742
rect 3374 53713 3402 53718
rect 4569 50175 4879 58961
rect 15904 59175 16064 59192
rect 15904 59147 15939 59175
rect 15967 59147 16001 59175
rect 16029 59147 16064 59175
rect 15904 59113 16064 59147
rect 15904 59085 15939 59113
rect 15967 59085 16001 59113
rect 16029 59085 16064 59113
rect 15904 59051 16064 59085
rect 15904 59023 15939 59051
rect 15967 59023 16001 59051
rect 16029 59023 16064 59051
rect 15904 58989 16064 59023
rect 15904 58961 15939 58989
rect 15967 58961 16001 58989
rect 16029 58961 16064 58989
rect 15904 58944 16064 58961
rect 8224 56175 8384 56192
rect 8224 56147 8259 56175
rect 8287 56147 8321 56175
rect 8349 56147 8384 56175
rect 8224 56113 8384 56147
rect 8224 56085 8259 56113
rect 8287 56085 8321 56113
rect 8349 56085 8384 56113
rect 8224 56051 8384 56085
rect 8224 56023 8259 56051
rect 8287 56023 8321 56051
rect 8349 56023 8384 56051
rect 8224 55989 8384 56023
rect 8224 55961 8259 55989
rect 8287 55961 8321 55989
rect 8349 55961 8384 55989
rect 8224 55944 8384 55961
rect 18069 56175 18379 64961
rect 18069 56147 18117 56175
rect 18145 56147 18179 56175
rect 18207 56147 18241 56175
rect 18269 56147 18303 56175
rect 18331 56147 18379 56175
rect 18069 56113 18379 56147
rect 18069 56085 18117 56113
rect 18145 56085 18179 56113
rect 18207 56085 18241 56113
rect 18269 56085 18303 56113
rect 18331 56085 18379 56113
rect 18069 56051 18379 56085
rect 18069 56023 18117 56051
rect 18145 56023 18179 56051
rect 18207 56023 18241 56051
rect 18269 56023 18303 56051
rect 18331 56023 18379 56051
rect 18069 55989 18379 56023
rect 18069 55961 18117 55989
rect 18145 55961 18179 55989
rect 18207 55961 18241 55989
rect 18269 55961 18303 55989
rect 18331 55961 18379 55989
rect 4569 50147 4617 50175
rect 4645 50147 4679 50175
rect 4707 50147 4741 50175
rect 4769 50147 4803 50175
rect 4831 50147 4879 50175
rect 4569 50113 4879 50147
rect 4569 50085 4617 50113
rect 4645 50085 4679 50113
rect 4707 50085 4741 50113
rect 4769 50085 4803 50113
rect 4831 50085 4879 50113
rect 4569 50051 4879 50085
rect 4569 50023 4617 50051
rect 4645 50023 4679 50051
rect 4707 50023 4741 50051
rect 4769 50023 4803 50051
rect 4831 50023 4879 50051
rect 4569 49989 4879 50023
rect 4569 49961 4617 49989
rect 4645 49961 4679 49989
rect 4707 49961 4741 49989
rect 4769 49961 4803 49989
rect 4831 49961 4879 49989
rect 2709 47147 2757 47175
rect 2785 47147 2819 47175
rect 2847 47147 2881 47175
rect 2909 47147 2943 47175
rect 2971 47147 3019 47175
rect 2709 47113 3019 47147
rect 2709 47085 2757 47113
rect 2785 47085 2819 47113
rect 2847 47085 2881 47113
rect 2909 47085 2943 47113
rect 2971 47085 3019 47113
rect 2709 47051 3019 47085
rect 2709 47023 2757 47051
rect 2785 47023 2819 47051
rect 2847 47023 2881 47051
rect 2909 47023 2943 47051
rect 2971 47023 3019 47051
rect 2709 46989 3019 47023
rect 2709 46961 2757 46989
rect 2785 46961 2819 46989
rect 2847 46961 2881 46989
rect 2909 46961 2943 46989
rect 2971 46961 3019 46989
rect 2709 38175 3019 46961
rect 3766 49490 3794 49495
rect 3766 46746 3794 49462
rect 3766 46713 3794 46718
rect 3766 42210 3794 42215
rect 3766 39690 3794 42182
rect 3766 39657 3794 39662
rect 4569 41175 4879 49961
rect 15904 50175 16064 50192
rect 15904 50147 15939 50175
rect 15967 50147 16001 50175
rect 16029 50147 16064 50175
rect 15904 50113 16064 50147
rect 15904 50085 15939 50113
rect 15967 50085 16001 50113
rect 16029 50085 16064 50113
rect 15904 50051 16064 50085
rect 15904 50023 15939 50051
rect 15967 50023 16001 50051
rect 16029 50023 16064 50051
rect 15904 49989 16064 50023
rect 15904 49961 15939 49989
rect 15967 49961 16001 49989
rect 16029 49961 16064 49989
rect 15904 49944 16064 49961
rect 8224 47175 8384 47192
rect 8224 47147 8259 47175
rect 8287 47147 8321 47175
rect 8349 47147 8384 47175
rect 8224 47113 8384 47147
rect 8224 47085 8259 47113
rect 8287 47085 8321 47113
rect 8349 47085 8384 47113
rect 8224 47051 8384 47085
rect 8224 47023 8259 47051
rect 8287 47023 8321 47051
rect 8349 47023 8384 47051
rect 8224 46989 8384 47023
rect 8224 46961 8259 46989
rect 8287 46961 8321 46989
rect 8349 46961 8384 46989
rect 8224 46944 8384 46961
rect 18069 47175 18379 55961
rect 18069 47147 18117 47175
rect 18145 47147 18179 47175
rect 18207 47147 18241 47175
rect 18269 47147 18303 47175
rect 18331 47147 18379 47175
rect 18069 47113 18379 47147
rect 18069 47085 18117 47113
rect 18145 47085 18179 47113
rect 18207 47085 18241 47113
rect 18269 47085 18303 47113
rect 18331 47085 18379 47113
rect 18069 47051 18379 47085
rect 18069 47023 18117 47051
rect 18145 47023 18179 47051
rect 18207 47023 18241 47051
rect 18269 47023 18303 47051
rect 18331 47023 18379 47051
rect 18069 46989 18379 47023
rect 18069 46961 18117 46989
rect 18145 46961 18179 46989
rect 18207 46961 18241 46989
rect 18269 46961 18303 46989
rect 18331 46961 18379 46989
rect 4569 41147 4617 41175
rect 4645 41147 4679 41175
rect 4707 41147 4741 41175
rect 4769 41147 4803 41175
rect 4831 41147 4879 41175
rect 4569 41113 4879 41147
rect 4569 41085 4617 41113
rect 4645 41085 4679 41113
rect 4707 41085 4741 41113
rect 4769 41085 4803 41113
rect 4831 41085 4879 41113
rect 4569 41051 4879 41085
rect 4569 41023 4617 41051
rect 4645 41023 4679 41051
rect 4707 41023 4741 41051
rect 4769 41023 4803 41051
rect 4831 41023 4879 41051
rect 4569 40989 4879 41023
rect 4569 40961 4617 40989
rect 4645 40961 4679 40989
rect 4707 40961 4741 40989
rect 4769 40961 4803 40989
rect 4831 40961 4879 40989
rect 2709 38147 2757 38175
rect 2785 38147 2819 38175
rect 2847 38147 2881 38175
rect 2909 38147 2943 38175
rect 2971 38147 3019 38175
rect 2709 38113 3019 38147
rect 2709 38085 2757 38113
rect 2785 38085 2819 38113
rect 2847 38085 2881 38113
rect 2909 38085 2943 38113
rect 2971 38085 3019 38113
rect 2709 38051 3019 38085
rect 2709 38023 2757 38051
rect 2785 38023 2819 38051
rect 2847 38023 2881 38051
rect 2909 38023 2943 38051
rect 2971 38023 3019 38051
rect 2709 37989 3019 38023
rect 2709 37961 2757 37989
rect 2785 37961 2819 37989
rect 2847 37961 2881 37989
rect 2909 37961 2943 37989
rect 2971 37961 3019 37989
rect 2709 29175 3019 37961
rect 3374 34930 3402 34935
rect 3374 32634 3402 34902
rect 3374 32601 3402 32606
rect 2709 29147 2757 29175
rect 2785 29147 2819 29175
rect 2847 29147 2881 29175
rect 2909 29147 2943 29175
rect 2971 29147 3019 29175
rect 2709 29113 3019 29147
rect 2709 29085 2757 29113
rect 2785 29085 2819 29113
rect 2847 29085 2881 29113
rect 2909 29085 2943 29113
rect 2971 29085 3019 29113
rect 2709 29051 3019 29085
rect 2709 29023 2757 29051
rect 2785 29023 2819 29051
rect 2847 29023 2881 29051
rect 2909 29023 2943 29051
rect 2971 29023 3019 29051
rect 2709 28989 3019 29023
rect 2709 28961 2757 28989
rect 2785 28961 2819 28989
rect 2847 28961 2881 28989
rect 2909 28961 2943 28989
rect 2971 28961 3019 28989
rect 2478 27650 2506 27655
rect 2478 25578 2506 27622
rect 2478 25545 2506 25550
rect -478 20147 -430 20175
rect -402 20147 -368 20175
rect -340 20147 -306 20175
rect -278 20147 -244 20175
rect -216 20147 -168 20175
rect -478 20113 -168 20147
rect -478 20085 -430 20113
rect -402 20085 -368 20113
rect -340 20085 -306 20113
rect -278 20085 -244 20113
rect -216 20085 -168 20113
rect -478 20051 -168 20085
rect -478 20023 -430 20051
rect -402 20023 -368 20051
rect -340 20023 -306 20051
rect -278 20023 -244 20051
rect -216 20023 -168 20051
rect -478 19989 -168 20023
rect -478 19961 -430 19989
rect -402 19961 -368 19989
rect -340 19961 -306 19989
rect -278 19961 -244 19989
rect -216 19961 -168 19989
rect -478 11175 -168 19961
rect 2709 20175 3019 28961
rect 4569 32175 4879 40961
rect 15904 41175 16064 41192
rect 15904 41147 15939 41175
rect 15967 41147 16001 41175
rect 16029 41147 16064 41175
rect 15904 41113 16064 41147
rect 15904 41085 15939 41113
rect 15967 41085 16001 41113
rect 16029 41085 16064 41113
rect 15904 41051 16064 41085
rect 15904 41023 15939 41051
rect 15967 41023 16001 41051
rect 16029 41023 16064 41051
rect 15904 40989 16064 41023
rect 15904 40961 15939 40989
rect 15967 40961 16001 40989
rect 16029 40961 16064 40989
rect 15904 40944 16064 40961
rect 8224 38175 8384 38192
rect 8224 38147 8259 38175
rect 8287 38147 8321 38175
rect 8349 38147 8384 38175
rect 8224 38113 8384 38147
rect 8224 38085 8259 38113
rect 8287 38085 8321 38113
rect 8349 38085 8384 38113
rect 8224 38051 8384 38085
rect 8224 38023 8259 38051
rect 8287 38023 8321 38051
rect 8349 38023 8384 38051
rect 8224 37989 8384 38023
rect 8224 37961 8259 37989
rect 8287 37961 8321 37989
rect 8349 37961 8384 37989
rect 8224 37944 8384 37961
rect 18069 38175 18379 46961
rect 18069 38147 18117 38175
rect 18145 38147 18179 38175
rect 18207 38147 18241 38175
rect 18269 38147 18303 38175
rect 18331 38147 18379 38175
rect 18069 38113 18379 38147
rect 18069 38085 18117 38113
rect 18145 38085 18179 38113
rect 18207 38085 18241 38113
rect 18269 38085 18303 38113
rect 18331 38085 18379 38113
rect 18069 38051 18379 38085
rect 18069 38023 18117 38051
rect 18145 38023 18179 38051
rect 18207 38023 18241 38051
rect 18269 38023 18303 38051
rect 18331 38023 18379 38051
rect 18069 37989 18379 38023
rect 18069 37961 18117 37989
rect 18145 37961 18179 37989
rect 18207 37961 18241 37989
rect 18269 37961 18303 37989
rect 18331 37961 18379 37989
rect 4569 32147 4617 32175
rect 4645 32147 4679 32175
rect 4707 32147 4741 32175
rect 4769 32147 4803 32175
rect 4831 32147 4879 32175
rect 4569 32113 4879 32147
rect 4569 32085 4617 32113
rect 4645 32085 4679 32113
rect 4707 32085 4741 32113
rect 4769 32085 4803 32113
rect 4831 32085 4879 32113
rect 4569 32051 4879 32085
rect 4569 32023 4617 32051
rect 4645 32023 4679 32051
rect 4707 32023 4741 32051
rect 4769 32023 4803 32051
rect 4831 32023 4879 32051
rect 4569 31989 4879 32023
rect 4569 31961 4617 31989
rect 4645 31961 4679 31989
rect 4707 31961 4741 31989
rect 4769 31961 4803 31989
rect 4831 31961 4879 31989
rect 4569 23175 4879 31961
rect 15904 32175 16064 32192
rect 15904 32147 15939 32175
rect 15967 32147 16001 32175
rect 16029 32147 16064 32175
rect 15904 32113 16064 32147
rect 15904 32085 15939 32113
rect 15967 32085 16001 32113
rect 16029 32085 16064 32113
rect 15904 32051 16064 32085
rect 15904 32023 15939 32051
rect 15967 32023 16001 32051
rect 16029 32023 16064 32051
rect 15904 31989 16064 32023
rect 15904 31961 15939 31989
rect 15967 31961 16001 31989
rect 16029 31961 16064 31989
rect 15904 31944 16064 31961
rect 8224 29175 8384 29192
rect 8224 29147 8259 29175
rect 8287 29147 8321 29175
rect 8349 29147 8384 29175
rect 8224 29113 8384 29147
rect 8224 29085 8259 29113
rect 8287 29085 8321 29113
rect 8349 29085 8384 29113
rect 8224 29051 8384 29085
rect 8224 29023 8259 29051
rect 8287 29023 8321 29051
rect 8349 29023 8384 29051
rect 8224 28989 8384 29023
rect 8224 28961 8259 28989
rect 8287 28961 8321 28989
rect 8349 28961 8384 28989
rect 8224 28944 8384 28961
rect 18069 29175 18379 37961
rect 18069 29147 18117 29175
rect 18145 29147 18179 29175
rect 18207 29147 18241 29175
rect 18269 29147 18303 29175
rect 18331 29147 18379 29175
rect 18069 29113 18379 29147
rect 18069 29085 18117 29113
rect 18145 29085 18179 29113
rect 18207 29085 18241 29113
rect 18269 29085 18303 29113
rect 18331 29085 18379 29113
rect 18069 29051 18379 29085
rect 18069 29023 18117 29051
rect 18145 29023 18179 29051
rect 18207 29023 18241 29051
rect 18269 29023 18303 29051
rect 18331 29023 18379 29051
rect 18069 28989 18379 29023
rect 18069 28961 18117 28989
rect 18145 28961 18179 28989
rect 18207 28961 18241 28989
rect 18269 28961 18303 28989
rect 18331 28961 18379 28989
rect 4569 23147 4617 23175
rect 4645 23147 4679 23175
rect 4707 23147 4741 23175
rect 4769 23147 4803 23175
rect 4831 23147 4879 23175
rect 4569 23113 4879 23147
rect 4569 23085 4617 23113
rect 4645 23085 4679 23113
rect 4707 23085 4741 23113
rect 4769 23085 4803 23113
rect 4831 23085 4879 23113
rect 4569 23051 4879 23085
rect 4569 23023 4617 23051
rect 4645 23023 4679 23051
rect 4707 23023 4741 23051
rect 4769 23023 4803 23051
rect 4831 23023 4879 23051
rect 4569 22989 4879 23023
rect 4569 22961 4617 22989
rect 4645 22961 4679 22989
rect 4707 22961 4741 22989
rect 4769 22961 4803 22989
rect 4831 22961 4879 22989
rect 2709 20147 2757 20175
rect 2785 20147 2819 20175
rect 2847 20147 2881 20175
rect 2909 20147 2943 20175
rect 2971 20147 3019 20175
rect 2709 20113 3019 20147
rect 2709 20085 2757 20113
rect 2785 20085 2819 20113
rect 2847 20085 2881 20113
rect 2909 20085 2943 20113
rect 2971 20085 3019 20113
rect 2709 20051 3019 20085
rect 2709 20023 2757 20051
rect 2785 20023 2819 20051
rect 2847 20023 2881 20051
rect 2909 20023 2943 20051
rect 2971 20023 3019 20051
rect 2709 19989 3019 20023
rect 2709 19961 2757 19989
rect 2785 19961 2819 19989
rect 2847 19961 2881 19989
rect 2909 19961 2943 19989
rect 2971 19961 3019 19989
rect 2086 13090 2114 13095
rect 2086 11466 2114 13062
rect 2086 11433 2114 11438
rect -478 11147 -430 11175
rect -402 11147 -368 11175
rect -340 11147 -306 11175
rect -278 11147 -244 11175
rect -216 11147 -168 11175
rect -478 11113 -168 11147
rect -478 11085 -430 11113
rect -402 11085 -368 11113
rect -340 11085 -306 11113
rect -278 11085 -244 11113
rect -216 11085 -168 11113
rect -478 11051 -168 11085
rect -478 11023 -430 11051
rect -402 11023 -368 11051
rect -340 11023 -306 11051
rect -278 11023 -244 11051
rect -216 11023 -168 11051
rect -478 10989 -168 11023
rect -478 10961 -430 10989
rect -402 10961 -368 10989
rect -340 10961 -306 10989
rect -278 10961 -244 10989
rect -216 10961 -168 10989
rect -478 2175 -168 10961
rect -478 2147 -430 2175
rect -402 2147 -368 2175
rect -340 2147 -306 2175
rect -278 2147 -244 2175
rect -216 2147 -168 2175
rect -478 2113 -168 2147
rect -478 2085 -430 2113
rect -402 2085 -368 2113
rect -340 2085 -306 2113
rect -278 2085 -244 2113
rect -216 2085 -168 2113
rect -478 2051 -168 2085
rect -478 2023 -430 2051
rect -402 2023 -368 2051
rect -340 2023 -306 2051
rect -278 2023 -244 2051
rect -216 2023 -168 2051
rect -478 1989 -168 2023
rect -478 1961 -430 1989
rect -402 1961 -368 1989
rect -340 1961 -306 1989
rect -278 1961 -244 1989
rect -216 1961 -168 1989
rect -478 -80 -168 1961
rect -478 -108 -430 -80
rect -402 -108 -368 -80
rect -340 -108 -306 -80
rect -278 -108 -244 -80
rect -216 -108 -168 -80
rect -478 -142 -168 -108
rect -478 -170 -430 -142
rect -402 -170 -368 -142
rect -340 -170 -306 -142
rect -278 -170 -244 -142
rect -216 -170 -168 -142
rect -478 -204 -168 -170
rect -478 -232 -430 -204
rect -402 -232 -368 -204
rect -340 -232 -306 -204
rect -278 -232 -244 -204
rect -216 -232 -168 -204
rect -478 -266 -168 -232
rect -478 -294 -430 -266
rect -402 -294 -368 -266
rect -340 -294 -306 -266
rect -278 -294 -244 -266
rect -216 -294 -168 -266
rect -478 -342 -168 -294
rect 2709 11175 3019 19961
rect 3374 20370 3402 20375
rect 3374 18466 3402 20342
rect 3374 18433 3402 18438
rect 2709 11147 2757 11175
rect 2785 11147 2819 11175
rect 2847 11147 2881 11175
rect 2909 11147 2943 11175
rect 2971 11147 3019 11175
rect 2709 11113 3019 11147
rect 2709 11085 2757 11113
rect 2785 11085 2819 11113
rect 2847 11085 2881 11113
rect 2909 11085 2943 11113
rect 2971 11085 3019 11113
rect 2709 11051 3019 11085
rect 2709 11023 2757 11051
rect 2785 11023 2819 11051
rect 2847 11023 2881 11051
rect 2909 11023 2943 11051
rect 2971 11023 3019 11051
rect 2709 10989 3019 11023
rect 2709 10961 2757 10989
rect 2785 10961 2819 10989
rect 2847 10961 2881 10989
rect 2909 10961 2943 10989
rect 2971 10961 3019 10989
rect 2709 2175 3019 10961
rect 4569 14175 4879 22961
rect 15904 23175 16064 23192
rect 15904 23147 15939 23175
rect 15967 23147 16001 23175
rect 16029 23147 16064 23175
rect 15904 23113 16064 23147
rect 15904 23085 15939 23113
rect 15967 23085 16001 23113
rect 16029 23085 16064 23113
rect 15904 23051 16064 23085
rect 15904 23023 15939 23051
rect 15967 23023 16001 23051
rect 16029 23023 16064 23051
rect 15904 22989 16064 23023
rect 15904 22961 15939 22989
rect 15967 22961 16001 22989
rect 16029 22961 16064 22989
rect 15904 22944 16064 22961
rect 8224 20175 8384 20192
rect 8224 20147 8259 20175
rect 8287 20147 8321 20175
rect 8349 20147 8384 20175
rect 8224 20113 8384 20147
rect 8224 20085 8259 20113
rect 8287 20085 8321 20113
rect 8349 20085 8384 20113
rect 8224 20051 8384 20085
rect 8224 20023 8259 20051
rect 8287 20023 8321 20051
rect 8349 20023 8384 20051
rect 8224 19989 8384 20023
rect 8224 19961 8259 19989
rect 8287 19961 8321 19989
rect 8349 19961 8384 19989
rect 8224 19944 8384 19961
rect 18069 20175 18379 28961
rect 18069 20147 18117 20175
rect 18145 20147 18179 20175
rect 18207 20147 18241 20175
rect 18269 20147 18303 20175
rect 18331 20147 18379 20175
rect 18069 20113 18379 20147
rect 18069 20085 18117 20113
rect 18145 20085 18179 20113
rect 18207 20085 18241 20113
rect 18269 20085 18303 20113
rect 18331 20085 18379 20113
rect 18069 20051 18379 20085
rect 18069 20023 18117 20051
rect 18145 20023 18179 20051
rect 18207 20023 18241 20051
rect 18269 20023 18303 20051
rect 18331 20023 18379 20051
rect 18069 19989 18379 20023
rect 18069 19961 18117 19989
rect 18145 19961 18179 19989
rect 18207 19961 18241 19989
rect 18269 19961 18303 19989
rect 18331 19961 18379 19989
rect 4569 14147 4617 14175
rect 4645 14147 4679 14175
rect 4707 14147 4741 14175
rect 4769 14147 4803 14175
rect 4831 14147 4879 14175
rect 4569 14113 4879 14147
rect 4569 14085 4617 14113
rect 4645 14085 4679 14113
rect 4707 14085 4741 14113
rect 4769 14085 4803 14113
rect 4831 14085 4879 14113
rect 4569 14051 4879 14085
rect 4569 14023 4617 14051
rect 4645 14023 4679 14051
rect 4707 14023 4741 14051
rect 4769 14023 4803 14051
rect 4831 14023 4879 14051
rect 4569 13989 4879 14023
rect 4569 13961 4617 13989
rect 4645 13961 4679 13989
rect 4707 13961 4741 13989
rect 4769 13961 4803 13989
rect 4831 13961 4879 13989
rect 3374 5810 3402 5815
rect 3374 4410 3402 5782
rect 3374 4377 3402 4382
rect 4569 5175 4879 13961
rect 15904 14175 16064 14192
rect 15904 14147 15939 14175
rect 15967 14147 16001 14175
rect 16029 14147 16064 14175
rect 15904 14113 16064 14147
rect 15904 14085 15939 14113
rect 15967 14085 16001 14113
rect 16029 14085 16064 14113
rect 15904 14051 16064 14085
rect 15904 14023 15939 14051
rect 15967 14023 16001 14051
rect 16029 14023 16064 14051
rect 15904 13989 16064 14023
rect 15904 13961 15939 13989
rect 15967 13961 16001 13989
rect 16029 13961 16064 13989
rect 15904 13944 16064 13961
rect 8224 11175 8384 11192
rect 8224 11147 8259 11175
rect 8287 11147 8321 11175
rect 8349 11147 8384 11175
rect 8224 11113 8384 11147
rect 8224 11085 8259 11113
rect 8287 11085 8321 11113
rect 8349 11085 8384 11113
rect 8224 11051 8384 11085
rect 8224 11023 8259 11051
rect 8287 11023 8321 11051
rect 8349 11023 8384 11051
rect 8224 10989 8384 11023
rect 8224 10961 8259 10989
rect 8287 10961 8321 10989
rect 8349 10961 8384 10989
rect 8224 10944 8384 10961
rect 18069 11175 18379 19961
rect 18069 11147 18117 11175
rect 18145 11147 18179 11175
rect 18207 11147 18241 11175
rect 18269 11147 18303 11175
rect 18331 11147 18379 11175
rect 18069 11113 18379 11147
rect 18069 11085 18117 11113
rect 18145 11085 18179 11113
rect 18207 11085 18241 11113
rect 18269 11085 18303 11113
rect 18331 11085 18379 11113
rect 18069 11051 18379 11085
rect 18069 11023 18117 11051
rect 18145 11023 18179 11051
rect 18207 11023 18241 11051
rect 18269 11023 18303 11051
rect 18331 11023 18379 11051
rect 18069 10989 18379 11023
rect 18069 10961 18117 10989
rect 18145 10961 18179 10989
rect 18207 10961 18241 10989
rect 18269 10961 18303 10989
rect 18331 10961 18379 10989
rect 4569 5147 4617 5175
rect 4645 5147 4679 5175
rect 4707 5147 4741 5175
rect 4769 5147 4803 5175
rect 4831 5147 4879 5175
rect 4569 5113 4879 5147
rect 4569 5085 4617 5113
rect 4645 5085 4679 5113
rect 4707 5085 4741 5113
rect 4769 5085 4803 5113
rect 4831 5085 4879 5113
rect 4569 5051 4879 5085
rect 4569 5023 4617 5051
rect 4645 5023 4679 5051
rect 4707 5023 4741 5051
rect 4769 5023 4803 5051
rect 4831 5023 4879 5051
rect 4569 4989 4879 5023
rect 4569 4961 4617 4989
rect 4645 4961 4679 4989
rect 4707 4961 4741 4989
rect 4769 4961 4803 4989
rect 4831 4961 4879 4989
rect 2709 2147 2757 2175
rect 2785 2147 2819 2175
rect 2847 2147 2881 2175
rect 2909 2147 2943 2175
rect 2971 2147 3019 2175
rect 2709 2113 3019 2147
rect 2709 2085 2757 2113
rect 2785 2085 2819 2113
rect 2847 2085 2881 2113
rect 2909 2085 2943 2113
rect 2971 2085 3019 2113
rect 2709 2051 3019 2085
rect 2709 2023 2757 2051
rect 2785 2023 2819 2051
rect 2847 2023 2881 2051
rect 2909 2023 2943 2051
rect 2971 2023 3019 2051
rect 2709 1989 3019 2023
rect 2709 1961 2757 1989
rect 2785 1961 2819 1989
rect 2847 1961 2881 1989
rect 2909 1961 2943 1989
rect 2971 1961 3019 1989
rect 2709 -80 3019 1961
rect 2709 -108 2757 -80
rect 2785 -108 2819 -80
rect 2847 -108 2881 -80
rect 2909 -108 2943 -80
rect 2971 -108 3019 -80
rect 2709 -142 3019 -108
rect 2709 -170 2757 -142
rect 2785 -170 2819 -142
rect 2847 -170 2881 -142
rect 2909 -170 2943 -142
rect 2971 -170 3019 -142
rect 2709 -204 3019 -170
rect 2709 -232 2757 -204
rect 2785 -232 2819 -204
rect 2847 -232 2881 -204
rect 2909 -232 2943 -204
rect 2971 -232 3019 -204
rect 2709 -266 3019 -232
rect 2709 -294 2757 -266
rect 2785 -294 2819 -266
rect 2847 -294 2881 -266
rect 2909 -294 2943 -266
rect 2971 -294 3019 -266
rect -958 -588 -910 -560
rect -882 -588 -848 -560
rect -820 -588 -786 -560
rect -758 -588 -724 -560
rect -696 -588 -648 -560
rect -958 -622 -648 -588
rect -958 -650 -910 -622
rect -882 -650 -848 -622
rect -820 -650 -786 -622
rect -758 -650 -724 -622
rect -696 -650 -648 -622
rect -958 -684 -648 -650
rect -958 -712 -910 -684
rect -882 -712 -848 -684
rect -820 -712 -786 -684
rect -758 -712 -724 -684
rect -696 -712 -648 -684
rect -958 -746 -648 -712
rect -958 -774 -910 -746
rect -882 -774 -848 -746
rect -820 -774 -786 -746
rect -758 -774 -724 -746
rect -696 -774 -648 -746
rect -958 -822 -648 -774
rect 2709 -822 3019 -294
rect 4569 -560 4879 4961
rect 15904 5175 16064 5192
rect 15904 5147 15939 5175
rect 15967 5147 16001 5175
rect 16029 5147 16064 5175
rect 15904 5113 16064 5147
rect 15904 5085 15939 5113
rect 15967 5085 16001 5113
rect 16029 5085 16064 5113
rect 15904 5051 16064 5085
rect 15904 5023 15939 5051
rect 15967 5023 16001 5051
rect 16029 5023 16064 5051
rect 15904 4989 16064 5023
rect 15904 4961 15939 4989
rect 15967 4961 16001 4989
rect 16029 4961 16064 4989
rect 15904 4944 16064 4961
rect 4569 -588 4617 -560
rect 4645 -588 4679 -560
rect 4707 -588 4741 -560
rect 4769 -588 4803 -560
rect 4831 -588 4879 -560
rect 4569 -622 4879 -588
rect 4569 -650 4617 -622
rect 4645 -650 4679 -622
rect 4707 -650 4741 -622
rect 4769 -650 4803 -622
rect 4831 -650 4879 -622
rect 4569 -684 4879 -650
rect 4569 -712 4617 -684
rect 4645 -712 4679 -684
rect 4707 -712 4741 -684
rect 4769 -712 4803 -684
rect 4831 -712 4879 -684
rect 4569 -746 4879 -712
rect 4569 -774 4617 -746
rect 4645 -774 4679 -746
rect 4707 -774 4741 -746
rect 4769 -774 4803 -746
rect 4831 -774 4879 -746
rect 4569 -822 4879 -774
rect 18069 2175 18379 10961
rect 18069 2147 18117 2175
rect 18145 2147 18179 2175
rect 18207 2147 18241 2175
rect 18269 2147 18303 2175
rect 18331 2147 18379 2175
rect 18069 2113 18379 2147
rect 18069 2085 18117 2113
rect 18145 2085 18179 2113
rect 18207 2085 18241 2113
rect 18269 2085 18303 2113
rect 18331 2085 18379 2113
rect 18069 2051 18379 2085
rect 18069 2023 18117 2051
rect 18145 2023 18179 2051
rect 18207 2023 18241 2051
rect 18269 2023 18303 2051
rect 18331 2023 18379 2051
rect 18069 1989 18379 2023
rect 18069 1961 18117 1989
rect 18145 1961 18179 1989
rect 18207 1961 18241 1989
rect 18269 1961 18303 1989
rect 18331 1961 18379 1989
rect 18069 -80 18379 1961
rect 18069 -108 18117 -80
rect 18145 -108 18179 -80
rect 18207 -108 18241 -80
rect 18269 -108 18303 -80
rect 18331 -108 18379 -80
rect 18069 -142 18379 -108
rect 18069 -170 18117 -142
rect 18145 -170 18179 -142
rect 18207 -170 18241 -142
rect 18269 -170 18303 -142
rect 18331 -170 18379 -142
rect 18069 -204 18379 -170
rect 18069 -232 18117 -204
rect 18145 -232 18179 -204
rect 18207 -232 18241 -204
rect 18269 -232 18303 -204
rect 18331 -232 18379 -204
rect 18069 -266 18379 -232
rect 18069 -294 18117 -266
rect 18145 -294 18179 -266
rect 18207 -294 18241 -266
rect 18269 -294 18303 -266
rect 18331 -294 18379 -266
rect 18069 -822 18379 -294
rect 19929 299086 20239 299134
rect 19929 299058 19977 299086
rect 20005 299058 20039 299086
rect 20067 299058 20101 299086
rect 20129 299058 20163 299086
rect 20191 299058 20239 299086
rect 19929 299024 20239 299058
rect 19929 298996 19977 299024
rect 20005 298996 20039 299024
rect 20067 298996 20101 299024
rect 20129 298996 20163 299024
rect 20191 298996 20239 299024
rect 19929 298962 20239 298996
rect 19929 298934 19977 298962
rect 20005 298934 20039 298962
rect 20067 298934 20101 298962
rect 20129 298934 20163 298962
rect 20191 298934 20239 298962
rect 19929 298900 20239 298934
rect 19929 298872 19977 298900
rect 20005 298872 20039 298900
rect 20067 298872 20101 298900
rect 20129 298872 20163 298900
rect 20191 298872 20239 298900
rect 19929 293175 20239 298872
rect 19929 293147 19977 293175
rect 20005 293147 20039 293175
rect 20067 293147 20101 293175
rect 20129 293147 20163 293175
rect 20191 293147 20239 293175
rect 19929 293113 20239 293147
rect 19929 293085 19977 293113
rect 20005 293085 20039 293113
rect 20067 293085 20101 293113
rect 20129 293085 20163 293113
rect 20191 293085 20239 293113
rect 19929 293051 20239 293085
rect 19929 293023 19977 293051
rect 20005 293023 20039 293051
rect 20067 293023 20101 293051
rect 20129 293023 20163 293051
rect 20191 293023 20239 293051
rect 19929 292989 20239 293023
rect 19929 292961 19977 292989
rect 20005 292961 20039 292989
rect 20067 292961 20101 292989
rect 20129 292961 20163 292989
rect 20191 292961 20239 292989
rect 19929 284175 20239 292961
rect 19929 284147 19977 284175
rect 20005 284147 20039 284175
rect 20067 284147 20101 284175
rect 20129 284147 20163 284175
rect 20191 284147 20239 284175
rect 19929 284113 20239 284147
rect 19929 284085 19977 284113
rect 20005 284085 20039 284113
rect 20067 284085 20101 284113
rect 20129 284085 20163 284113
rect 20191 284085 20239 284113
rect 19929 284051 20239 284085
rect 19929 284023 19977 284051
rect 20005 284023 20039 284051
rect 20067 284023 20101 284051
rect 20129 284023 20163 284051
rect 20191 284023 20239 284051
rect 19929 283989 20239 284023
rect 19929 283961 19977 283989
rect 20005 283961 20039 283989
rect 20067 283961 20101 283989
rect 20129 283961 20163 283989
rect 20191 283961 20239 283989
rect 19929 275175 20239 283961
rect 19929 275147 19977 275175
rect 20005 275147 20039 275175
rect 20067 275147 20101 275175
rect 20129 275147 20163 275175
rect 20191 275147 20239 275175
rect 19929 275113 20239 275147
rect 19929 275085 19977 275113
rect 20005 275085 20039 275113
rect 20067 275085 20101 275113
rect 20129 275085 20163 275113
rect 20191 275085 20239 275113
rect 19929 275051 20239 275085
rect 19929 275023 19977 275051
rect 20005 275023 20039 275051
rect 20067 275023 20101 275051
rect 20129 275023 20163 275051
rect 20191 275023 20239 275051
rect 19929 274989 20239 275023
rect 19929 274961 19977 274989
rect 20005 274961 20039 274989
rect 20067 274961 20101 274989
rect 20129 274961 20163 274989
rect 20191 274961 20239 274989
rect 19929 266175 20239 274961
rect 19929 266147 19977 266175
rect 20005 266147 20039 266175
rect 20067 266147 20101 266175
rect 20129 266147 20163 266175
rect 20191 266147 20239 266175
rect 19929 266113 20239 266147
rect 19929 266085 19977 266113
rect 20005 266085 20039 266113
rect 20067 266085 20101 266113
rect 20129 266085 20163 266113
rect 20191 266085 20239 266113
rect 19929 266051 20239 266085
rect 19929 266023 19977 266051
rect 20005 266023 20039 266051
rect 20067 266023 20101 266051
rect 20129 266023 20163 266051
rect 20191 266023 20239 266051
rect 19929 265989 20239 266023
rect 19929 265961 19977 265989
rect 20005 265961 20039 265989
rect 20067 265961 20101 265989
rect 20129 265961 20163 265989
rect 20191 265961 20239 265989
rect 19929 257175 20239 265961
rect 19929 257147 19977 257175
rect 20005 257147 20039 257175
rect 20067 257147 20101 257175
rect 20129 257147 20163 257175
rect 20191 257147 20239 257175
rect 19929 257113 20239 257147
rect 19929 257085 19977 257113
rect 20005 257085 20039 257113
rect 20067 257085 20101 257113
rect 20129 257085 20163 257113
rect 20191 257085 20239 257113
rect 19929 257051 20239 257085
rect 19929 257023 19977 257051
rect 20005 257023 20039 257051
rect 20067 257023 20101 257051
rect 20129 257023 20163 257051
rect 20191 257023 20239 257051
rect 19929 256989 20239 257023
rect 19929 256961 19977 256989
rect 20005 256961 20039 256989
rect 20067 256961 20101 256989
rect 20129 256961 20163 256989
rect 20191 256961 20239 256989
rect 19929 248175 20239 256961
rect 19929 248147 19977 248175
rect 20005 248147 20039 248175
rect 20067 248147 20101 248175
rect 20129 248147 20163 248175
rect 20191 248147 20239 248175
rect 19929 248113 20239 248147
rect 19929 248085 19977 248113
rect 20005 248085 20039 248113
rect 20067 248085 20101 248113
rect 20129 248085 20163 248113
rect 20191 248085 20239 248113
rect 19929 248051 20239 248085
rect 19929 248023 19977 248051
rect 20005 248023 20039 248051
rect 20067 248023 20101 248051
rect 20129 248023 20163 248051
rect 20191 248023 20239 248051
rect 19929 247989 20239 248023
rect 19929 247961 19977 247989
rect 20005 247961 20039 247989
rect 20067 247961 20101 247989
rect 20129 247961 20163 247989
rect 20191 247961 20239 247989
rect 19929 239175 20239 247961
rect 19929 239147 19977 239175
rect 20005 239147 20039 239175
rect 20067 239147 20101 239175
rect 20129 239147 20163 239175
rect 20191 239147 20239 239175
rect 19929 239113 20239 239147
rect 19929 239085 19977 239113
rect 20005 239085 20039 239113
rect 20067 239085 20101 239113
rect 20129 239085 20163 239113
rect 20191 239085 20239 239113
rect 19929 239051 20239 239085
rect 19929 239023 19977 239051
rect 20005 239023 20039 239051
rect 20067 239023 20101 239051
rect 20129 239023 20163 239051
rect 20191 239023 20239 239051
rect 19929 238989 20239 239023
rect 19929 238961 19977 238989
rect 20005 238961 20039 238989
rect 20067 238961 20101 238989
rect 20129 238961 20163 238989
rect 20191 238961 20239 238989
rect 19929 230175 20239 238961
rect 19929 230147 19977 230175
rect 20005 230147 20039 230175
rect 20067 230147 20101 230175
rect 20129 230147 20163 230175
rect 20191 230147 20239 230175
rect 19929 230113 20239 230147
rect 19929 230085 19977 230113
rect 20005 230085 20039 230113
rect 20067 230085 20101 230113
rect 20129 230085 20163 230113
rect 20191 230085 20239 230113
rect 19929 230051 20239 230085
rect 19929 230023 19977 230051
rect 20005 230023 20039 230051
rect 20067 230023 20101 230051
rect 20129 230023 20163 230051
rect 20191 230023 20239 230051
rect 19929 229989 20239 230023
rect 19929 229961 19977 229989
rect 20005 229961 20039 229989
rect 20067 229961 20101 229989
rect 20129 229961 20163 229989
rect 20191 229961 20239 229989
rect 19929 221175 20239 229961
rect 19929 221147 19977 221175
rect 20005 221147 20039 221175
rect 20067 221147 20101 221175
rect 20129 221147 20163 221175
rect 20191 221147 20239 221175
rect 19929 221113 20239 221147
rect 19929 221085 19977 221113
rect 20005 221085 20039 221113
rect 20067 221085 20101 221113
rect 20129 221085 20163 221113
rect 20191 221085 20239 221113
rect 19929 221051 20239 221085
rect 19929 221023 19977 221051
rect 20005 221023 20039 221051
rect 20067 221023 20101 221051
rect 20129 221023 20163 221051
rect 20191 221023 20239 221051
rect 19929 220989 20239 221023
rect 19929 220961 19977 220989
rect 20005 220961 20039 220989
rect 20067 220961 20101 220989
rect 20129 220961 20163 220989
rect 20191 220961 20239 220989
rect 19929 212175 20239 220961
rect 19929 212147 19977 212175
rect 20005 212147 20039 212175
rect 20067 212147 20101 212175
rect 20129 212147 20163 212175
rect 20191 212147 20239 212175
rect 19929 212113 20239 212147
rect 19929 212085 19977 212113
rect 20005 212085 20039 212113
rect 20067 212085 20101 212113
rect 20129 212085 20163 212113
rect 20191 212085 20239 212113
rect 19929 212051 20239 212085
rect 19929 212023 19977 212051
rect 20005 212023 20039 212051
rect 20067 212023 20101 212051
rect 20129 212023 20163 212051
rect 20191 212023 20239 212051
rect 19929 211989 20239 212023
rect 19929 211961 19977 211989
rect 20005 211961 20039 211989
rect 20067 211961 20101 211989
rect 20129 211961 20163 211989
rect 20191 211961 20239 211989
rect 19929 203175 20239 211961
rect 19929 203147 19977 203175
rect 20005 203147 20039 203175
rect 20067 203147 20101 203175
rect 20129 203147 20163 203175
rect 20191 203147 20239 203175
rect 19929 203113 20239 203147
rect 19929 203085 19977 203113
rect 20005 203085 20039 203113
rect 20067 203085 20101 203113
rect 20129 203085 20163 203113
rect 20191 203085 20239 203113
rect 19929 203051 20239 203085
rect 19929 203023 19977 203051
rect 20005 203023 20039 203051
rect 20067 203023 20101 203051
rect 20129 203023 20163 203051
rect 20191 203023 20239 203051
rect 19929 202989 20239 203023
rect 19929 202961 19977 202989
rect 20005 202961 20039 202989
rect 20067 202961 20101 202989
rect 20129 202961 20163 202989
rect 20191 202961 20239 202989
rect 19929 194175 20239 202961
rect 19929 194147 19977 194175
rect 20005 194147 20039 194175
rect 20067 194147 20101 194175
rect 20129 194147 20163 194175
rect 20191 194147 20239 194175
rect 19929 194113 20239 194147
rect 19929 194085 19977 194113
rect 20005 194085 20039 194113
rect 20067 194085 20101 194113
rect 20129 194085 20163 194113
rect 20191 194085 20239 194113
rect 19929 194051 20239 194085
rect 19929 194023 19977 194051
rect 20005 194023 20039 194051
rect 20067 194023 20101 194051
rect 20129 194023 20163 194051
rect 20191 194023 20239 194051
rect 19929 193989 20239 194023
rect 19929 193961 19977 193989
rect 20005 193961 20039 193989
rect 20067 193961 20101 193989
rect 20129 193961 20163 193989
rect 20191 193961 20239 193989
rect 19929 185175 20239 193961
rect 19929 185147 19977 185175
rect 20005 185147 20039 185175
rect 20067 185147 20101 185175
rect 20129 185147 20163 185175
rect 20191 185147 20239 185175
rect 19929 185113 20239 185147
rect 19929 185085 19977 185113
rect 20005 185085 20039 185113
rect 20067 185085 20101 185113
rect 20129 185085 20163 185113
rect 20191 185085 20239 185113
rect 19929 185051 20239 185085
rect 19929 185023 19977 185051
rect 20005 185023 20039 185051
rect 20067 185023 20101 185051
rect 20129 185023 20163 185051
rect 20191 185023 20239 185051
rect 19929 184989 20239 185023
rect 19929 184961 19977 184989
rect 20005 184961 20039 184989
rect 20067 184961 20101 184989
rect 20129 184961 20163 184989
rect 20191 184961 20239 184989
rect 19929 176175 20239 184961
rect 19929 176147 19977 176175
rect 20005 176147 20039 176175
rect 20067 176147 20101 176175
rect 20129 176147 20163 176175
rect 20191 176147 20239 176175
rect 19929 176113 20239 176147
rect 19929 176085 19977 176113
rect 20005 176085 20039 176113
rect 20067 176085 20101 176113
rect 20129 176085 20163 176113
rect 20191 176085 20239 176113
rect 19929 176051 20239 176085
rect 19929 176023 19977 176051
rect 20005 176023 20039 176051
rect 20067 176023 20101 176051
rect 20129 176023 20163 176051
rect 20191 176023 20239 176051
rect 19929 175989 20239 176023
rect 19929 175961 19977 175989
rect 20005 175961 20039 175989
rect 20067 175961 20101 175989
rect 20129 175961 20163 175989
rect 20191 175961 20239 175989
rect 19929 167175 20239 175961
rect 33429 298606 33739 299134
rect 33429 298578 33477 298606
rect 33505 298578 33539 298606
rect 33567 298578 33601 298606
rect 33629 298578 33663 298606
rect 33691 298578 33739 298606
rect 33429 298544 33739 298578
rect 33429 298516 33477 298544
rect 33505 298516 33539 298544
rect 33567 298516 33601 298544
rect 33629 298516 33663 298544
rect 33691 298516 33739 298544
rect 33429 298482 33739 298516
rect 33429 298454 33477 298482
rect 33505 298454 33539 298482
rect 33567 298454 33601 298482
rect 33629 298454 33663 298482
rect 33691 298454 33739 298482
rect 33429 298420 33739 298454
rect 33429 298392 33477 298420
rect 33505 298392 33539 298420
rect 33567 298392 33601 298420
rect 33629 298392 33663 298420
rect 33691 298392 33739 298420
rect 33429 290175 33739 298392
rect 33429 290147 33477 290175
rect 33505 290147 33539 290175
rect 33567 290147 33601 290175
rect 33629 290147 33663 290175
rect 33691 290147 33739 290175
rect 33429 290113 33739 290147
rect 33429 290085 33477 290113
rect 33505 290085 33539 290113
rect 33567 290085 33601 290113
rect 33629 290085 33663 290113
rect 33691 290085 33739 290113
rect 33429 290051 33739 290085
rect 33429 290023 33477 290051
rect 33505 290023 33539 290051
rect 33567 290023 33601 290051
rect 33629 290023 33663 290051
rect 33691 290023 33739 290051
rect 33429 289989 33739 290023
rect 33429 289961 33477 289989
rect 33505 289961 33539 289989
rect 33567 289961 33601 289989
rect 33629 289961 33663 289989
rect 33691 289961 33739 289989
rect 33429 281175 33739 289961
rect 33429 281147 33477 281175
rect 33505 281147 33539 281175
rect 33567 281147 33601 281175
rect 33629 281147 33663 281175
rect 33691 281147 33739 281175
rect 33429 281113 33739 281147
rect 33429 281085 33477 281113
rect 33505 281085 33539 281113
rect 33567 281085 33601 281113
rect 33629 281085 33663 281113
rect 33691 281085 33739 281113
rect 33429 281051 33739 281085
rect 33429 281023 33477 281051
rect 33505 281023 33539 281051
rect 33567 281023 33601 281051
rect 33629 281023 33663 281051
rect 33691 281023 33739 281051
rect 33429 280989 33739 281023
rect 33429 280961 33477 280989
rect 33505 280961 33539 280989
rect 33567 280961 33601 280989
rect 33629 280961 33663 280989
rect 33691 280961 33739 280989
rect 33429 272175 33739 280961
rect 33429 272147 33477 272175
rect 33505 272147 33539 272175
rect 33567 272147 33601 272175
rect 33629 272147 33663 272175
rect 33691 272147 33739 272175
rect 33429 272113 33739 272147
rect 33429 272085 33477 272113
rect 33505 272085 33539 272113
rect 33567 272085 33601 272113
rect 33629 272085 33663 272113
rect 33691 272085 33739 272113
rect 33429 272051 33739 272085
rect 33429 272023 33477 272051
rect 33505 272023 33539 272051
rect 33567 272023 33601 272051
rect 33629 272023 33663 272051
rect 33691 272023 33739 272051
rect 33429 271989 33739 272023
rect 33429 271961 33477 271989
rect 33505 271961 33539 271989
rect 33567 271961 33601 271989
rect 33629 271961 33663 271989
rect 33691 271961 33739 271989
rect 33429 263175 33739 271961
rect 33429 263147 33477 263175
rect 33505 263147 33539 263175
rect 33567 263147 33601 263175
rect 33629 263147 33663 263175
rect 33691 263147 33739 263175
rect 33429 263113 33739 263147
rect 33429 263085 33477 263113
rect 33505 263085 33539 263113
rect 33567 263085 33601 263113
rect 33629 263085 33663 263113
rect 33691 263085 33739 263113
rect 33429 263051 33739 263085
rect 33429 263023 33477 263051
rect 33505 263023 33539 263051
rect 33567 263023 33601 263051
rect 33629 263023 33663 263051
rect 33691 263023 33739 263051
rect 33429 262989 33739 263023
rect 33429 262961 33477 262989
rect 33505 262961 33539 262989
rect 33567 262961 33601 262989
rect 33629 262961 33663 262989
rect 33691 262961 33739 262989
rect 33429 254175 33739 262961
rect 33429 254147 33477 254175
rect 33505 254147 33539 254175
rect 33567 254147 33601 254175
rect 33629 254147 33663 254175
rect 33691 254147 33739 254175
rect 33429 254113 33739 254147
rect 33429 254085 33477 254113
rect 33505 254085 33539 254113
rect 33567 254085 33601 254113
rect 33629 254085 33663 254113
rect 33691 254085 33739 254113
rect 33429 254051 33739 254085
rect 33429 254023 33477 254051
rect 33505 254023 33539 254051
rect 33567 254023 33601 254051
rect 33629 254023 33663 254051
rect 33691 254023 33739 254051
rect 33429 253989 33739 254023
rect 33429 253961 33477 253989
rect 33505 253961 33539 253989
rect 33567 253961 33601 253989
rect 33629 253961 33663 253989
rect 33691 253961 33739 253989
rect 33429 245175 33739 253961
rect 33429 245147 33477 245175
rect 33505 245147 33539 245175
rect 33567 245147 33601 245175
rect 33629 245147 33663 245175
rect 33691 245147 33739 245175
rect 33429 245113 33739 245147
rect 33429 245085 33477 245113
rect 33505 245085 33539 245113
rect 33567 245085 33601 245113
rect 33629 245085 33663 245113
rect 33691 245085 33739 245113
rect 33429 245051 33739 245085
rect 33429 245023 33477 245051
rect 33505 245023 33539 245051
rect 33567 245023 33601 245051
rect 33629 245023 33663 245051
rect 33691 245023 33739 245051
rect 33429 244989 33739 245023
rect 33429 244961 33477 244989
rect 33505 244961 33539 244989
rect 33567 244961 33601 244989
rect 33629 244961 33663 244989
rect 33691 244961 33739 244989
rect 33429 236175 33739 244961
rect 33429 236147 33477 236175
rect 33505 236147 33539 236175
rect 33567 236147 33601 236175
rect 33629 236147 33663 236175
rect 33691 236147 33739 236175
rect 33429 236113 33739 236147
rect 33429 236085 33477 236113
rect 33505 236085 33539 236113
rect 33567 236085 33601 236113
rect 33629 236085 33663 236113
rect 33691 236085 33739 236113
rect 33429 236051 33739 236085
rect 33429 236023 33477 236051
rect 33505 236023 33539 236051
rect 33567 236023 33601 236051
rect 33629 236023 33663 236051
rect 33691 236023 33739 236051
rect 33429 235989 33739 236023
rect 33429 235961 33477 235989
rect 33505 235961 33539 235989
rect 33567 235961 33601 235989
rect 33629 235961 33663 235989
rect 33691 235961 33739 235989
rect 33429 227175 33739 235961
rect 33429 227147 33477 227175
rect 33505 227147 33539 227175
rect 33567 227147 33601 227175
rect 33629 227147 33663 227175
rect 33691 227147 33739 227175
rect 33429 227113 33739 227147
rect 33429 227085 33477 227113
rect 33505 227085 33539 227113
rect 33567 227085 33601 227113
rect 33629 227085 33663 227113
rect 33691 227085 33739 227113
rect 33429 227051 33739 227085
rect 33429 227023 33477 227051
rect 33505 227023 33539 227051
rect 33567 227023 33601 227051
rect 33629 227023 33663 227051
rect 33691 227023 33739 227051
rect 33429 226989 33739 227023
rect 33429 226961 33477 226989
rect 33505 226961 33539 226989
rect 33567 226961 33601 226989
rect 33629 226961 33663 226989
rect 33691 226961 33739 226989
rect 33429 218175 33739 226961
rect 33429 218147 33477 218175
rect 33505 218147 33539 218175
rect 33567 218147 33601 218175
rect 33629 218147 33663 218175
rect 33691 218147 33739 218175
rect 33429 218113 33739 218147
rect 33429 218085 33477 218113
rect 33505 218085 33539 218113
rect 33567 218085 33601 218113
rect 33629 218085 33663 218113
rect 33691 218085 33739 218113
rect 33429 218051 33739 218085
rect 33429 218023 33477 218051
rect 33505 218023 33539 218051
rect 33567 218023 33601 218051
rect 33629 218023 33663 218051
rect 33691 218023 33739 218051
rect 33429 217989 33739 218023
rect 33429 217961 33477 217989
rect 33505 217961 33539 217989
rect 33567 217961 33601 217989
rect 33629 217961 33663 217989
rect 33691 217961 33739 217989
rect 33429 209175 33739 217961
rect 33429 209147 33477 209175
rect 33505 209147 33539 209175
rect 33567 209147 33601 209175
rect 33629 209147 33663 209175
rect 33691 209147 33739 209175
rect 33429 209113 33739 209147
rect 33429 209085 33477 209113
rect 33505 209085 33539 209113
rect 33567 209085 33601 209113
rect 33629 209085 33663 209113
rect 33691 209085 33739 209113
rect 33429 209051 33739 209085
rect 33429 209023 33477 209051
rect 33505 209023 33539 209051
rect 33567 209023 33601 209051
rect 33629 209023 33663 209051
rect 33691 209023 33739 209051
rect 33429 208989 33739 209023
rect 33429 208961 33477 208989
rect 33505 208961 33539 208989
rect 33567 208961 33601 208989
rect 33629 208961 33663 208989
rect 33691 208961 33739 208989
rect 33429 200175 33739 208961
rect 33429 200147 33477 200175
rect 33505 200147 33539 200175
rect 33567 200147 33601 200175
rect 33629 200147 33663 200175
rect 33691 200147 33739 200175
rect 33429 200113 33739 200147
rect 33429 200085 33477 200113
rect 33505 200085 33539 200113
rect 33567 200085 33601 200113
rect 33629 200085 33663 200113
rect 33691 200085 33739 200113
rect 33429 200051 33739 200085
rect 33429 200023 33477 200051
rect 33505 200023 33539 200051
rect 33567 200023 33601 200051
rect 33629 200023 33663 200051
rect 33691 200023 33739 200051
rect 33429 199989 33739 200023
rect 33429 199961 33477 199989
rect 33505 199961 33539 199989
rect 33567 199961 33601 199989
rect 33629 199961 33663 199989
rect 33691 199961 33739 199989
rect 33429 191175 33739 199961
rect 33429 191147 33477 191175
rect 33505 191147 33539 191175
rect 33567 191147 33601 191175
rect 33629 191147 33663 191175
rect 33691 191147 33739 191175
rect 33429 191113 33739 191147
rect 33429 191085 33477 191113
rect 33505 191085 33539 191113
rect 33567 191085 33601 191113
rect 33629 191085 33663 191113
rect 33691 191085 33739 191113
rect 33429 191051 33739 191085
rect 33429 191023 33477 191051
rect 33505 191023 33539 191051
rect 33567 191023 33601 191051
rect 33629 191023 33663 191051
rect 33691 191023 33739 191051
rect 33429 190989 33739 191023
rect 33429 190961 33477 190989
rect 33505 190961 33539 190989
rect 33567 190961 33601 190989
rect 33629 190961 33663 190989
rect 33691 190961 33739 190989
rect 33429 182175 33739 190961
rect 33429 182147 33477 182175
rect 33505 182147 33539 182175
rect 33567 182147 33601 182175
rect 33629 182147 33663 182175
rect 33691 182147 33739 182175
rect 33429 182113 33739 182147
rect 33429 182085 33477 182113
rect 33505 182085 33539 182113
rect 33567 182085 33601 182113
rect 33629 182085 33663 182113
rect 33691 182085 33739 182113
rect 33429 182051 33739 182085
rect 33429 182023 33477 182051
rect 33505 182023 33539 182051
rect 33567 182023 33601 182051
rect 33629 182023 33663 182051
rect 33691 182023 33739 182051
rect 33429 181989 33739 182023
rect 33429 181961 33477 181989
rect 33505 181961 33539 181989
rect 33567 181961 33601 181989
rect 33629 181961 33663 181989
rect 33691 181961 33739 181989
rect 23584 173175 23744 173192
rect 23584 173147 23619 173175
rect 23647 173147 23681 173175
rect 23709 173147 23744 173175
rect 23584 173113 23744 173147
rect 23584 173085 23619 173113
rect 23647 173085 23681 173113
rect 23709 173085 23744 173113
rect 23584 173051 23744 173085
rect 23584 173023 23619 173051
rect 23647 173023 23681 173051
rect 23709 173023 23744 173051
rect 23584 172989 23744 173023
rect 23584 172961 23619 172989
rect 23647 172961 23681 172989
rect 23709 172961 23744 172989
rect 23584 172944 23744 172961
rect 33429 173175 33739 181961
rect 33429 173147 33477 173175
rect 33505 173147 33539 173175
rect 33567 173147 33601 173175
rect 33629 173147 33663 173175
rect 33691 173147 33739 173175
rect 33429 173113 33739 173147
rect 33429 173085 33477 173113
rect 33505 173085 33539 173113
rect 33567 173085 33601 173113
rect 33629 173085 33663 173113
rect 33691 173085 33739 173113
rect 33429 173051 33739 173085
rect 33429 173023 33477 173051
rect 33505 173023 33539 173051
rect 33567 173023 33601 173051
rect 33629 173023 33663 173051
rect 33691 173023 33739 173051
rect 33429 172989 33739 173023
rect 33429 172961 33477 172989
rect 33505 172961 33539 172989
rect 33567 172961 33601 172989
rect 33629 172961 33663 172989
rect 33691 172961 33739 172989
rect 19929 167147 19977 167175
rect 20005 167147 20039 167175
rect 20067 167147 20101 167175
rect 20129 167147 20163 167175
rect 20191 167147 20239 167175
rect 19929 167113 20239 167147
rect 19929 167085 19977 167113
rect 20005 167085 20039 167113
rect 20067 167085 20101 167113
rect 20129 167085 20163 167113
rect 20191 167085 20239 167113
rect 19929 167051 20239 167085
rect 19929 167023 19977 167051
rect 20005 167023 20039 167051
rect 20067 167023 20101 167051
rect 20129 167023 20163 167051
rect 20191 167023 20239 167051
rect 19929 166989 20239 167023
rect 19929 166961 19977 166989
rect 20005 166961 20039 166989
rect 20067 166961 20101 166989
rect 20129 166961 20163 166989
rect 20191 166961 20239 166989
rect 19929 158175 20239 166961
rect 31264 167175 31424 167192
rect 31264 167147 31299 167175
rect 31327 167147 31361 167175
rect 31389 167147 31424 167175
rect 31264 167113 31424 167147
rect 31264 167085 31299 167113
rect 31327 167085 31361 167113
rect 31389 167085 31424 167113
rect 31264 167051 31424 167085
rect 31264 167023 31299 167051
rect 31327 167023 31361 167051
rect 31389 167023 31424 167051
rect 31264 166989 31424 167023
rect 31264 166961 31299 166989
rect 31327 166961 31361 166989
rect 31389 166961 31424 166989
rect 31264 166944 31424 166961
rect 23584 164175 23744 164192
rect 23584 164147 23619 164175
rect 23647 164147 23681 164175
rect 23709 164147 23744 164175
rect 23584 164113 23744 164147
rect 23584 164085 23619 164113
rect 23647 164085 23681 164113
rect 23709 164085 23744 164113
rect 23584 164051 23744 164085
rect 23584 164023 23619 164051
rect 23647 164023 23681 164051
rect 23709 164023 23744 164051
rect 23584 163989 23744 164023
rect 23584 163961 23619 163989
rect 23647 163961 23681 163989
rect 23709 163961 23744 163989
rect 23584 163944 23744 163961
rect 33429 164175 33739 172961
rect 33429 164147 33477 164175
rect 33505 164147 33539 164175
rect 33567 164147 33601 164175
rect 33629 164147 33663 164175
rect 33691 164147 33739 164175
rect 33429 164113 33739 164147
rect 33429 164085 33477 164113
rect 33505 164085 33539 164113
rect 33567 164085 33601 164113
rect 33629 164085 33663 164113
rect 33691 164085 33739 164113
rect 33429 164051 33739 164085
rect 33429 164023 33477 164051
rect 33505 164023 33539 164051
rect 33567 164023 33601 164051
rect 33629 164023 33663 164051
rect 33691 164023 33739 164051
rect 33429 163989 33739 164023
rect 33429 163961 33477 163989
rect 33505 163961 33539 163989
rect 33567 163961 33601 163989
rect 33629 163961 33663 163989
rect 33691 163961 33739 163989
rect 19929 158147 19977 158175
rect 20005 158147 20039 158175
rect 20067 158147 20101 158175
rect 20129 158147 20163 158175
rect 20191 158147 20239 158175
rect 19929 158113 20239 158147
rect 19929 158085 19977 158113
rect 20005 158085 20039 158113
rect 20067 158085 20101 158113
rect 20129 158085 20163 158113
rect 20191 158085 20239 158113
rect 19929 158051 20239 158085
rect 19929 158023 19977 158051
rect 20005 158023 20039 158051
rect 20067 158023 20101 158051
rect 20129 158023 20163 158051
rect 20191 158023 20239 158051
rect 19929 157989 20239 158023
rect 19929 157961 19977 157989
rect 20005 157961 20039 157989
rect 20067 157961 20101 157989
rect 20129 157961 20163 157989
rect 20191 157961 20239 157989
rect 19929 149175 20239 157961
rect 31264 158175 31424 158192
rect 31264 158147 31299 158175
rect 31327 158147 31361 158175
rect 31389 158147 31424 158175
rect 31264 158113 31424 158147
rect 31264 158085 31299 158113
rect 31327 158085 31361 158113
rect 31389 158085 31424 158113
rect 31264 158051 31424 158085
rect 31264 158023 31299 158051
rect 31327 158023 31361 158051
rect 31389 158023 31424 158051
rect 31264 157989 31424 158023
rect 31264 157961 31299 157989
rect 31327 157961 31361 157989
rect 31389 157961 31424 157989
rect 31264 157944 31424 157961
rect 23584 155175 23744 155192
rect 23584 155147 23619 155175
rect 23647 155147 23681 155175
rect 23709 155147 23744 155175
rect 23584 155113 23744 155147
rect 23584 155085 23619 155113
rect 23647 155085 23681 155113
rect 23709 155085 23744 155113
rect 23584 155051 23744 155085
rect 23584 155023 23619 155051
rect 23647 155023 23681 155051
rect 23709 155023 23744 155051
rect 23584 154989 23744 155023
rect 23584 154961 23619 154989
rect 23647 154961 23681 154989
rect 23709 154961 23744 154989
rect 23584 154944 23744 154961
rect 33429 155175 33739 163961
rect 33429 155147 33477 155175
rect 33505 155147 33539 155175
rect 33567 155147 33601 155175
rect 33629 155147 33663 155175
rect 33691 155147 33739 155175
rect 33429 155113 33739 155147
rect 33429 155085 33477 155113
rect 33505 155085 33539 155113
rect 33567 155085 33601 155113
rect 33629 155085 33663 155113
rect 33691 155085 33739 155113
rect 33429 155051 33739 155085
rect 33429 155023 33477 155051
rect 33505 155023 33539 155051
rect 33567 155023 33601 155051
rect 33629 155023 33663 155051
rect 33691 155023 33739 155051
rect 33429 154989 33739 155023
rect 33429 154961 33477 154989
rect 33505 154961 33539 154989
rect 33567 154961 33601 154989
rect 33629 154961 33663 154989
rect 33691 154961 33739 154989
rect 19929 149147 19977 149175
rect 20005 149147 20039 149175
rect 20067 149147 20101 149175
rect 20129 149147 20163 149175
rect 20191 149147 20239 149175
rect 19929 149113 20239 149147
rect 19929 149085 19977 149113
rect 20005 149085 20039 149113
rect 20067 149085 20101 149113
rect 20129 149085 20163 149113
rect 20191 149085 20239 149113
rect 19929 149051 20239 149085
rect 19929 149023 19977 149051
rect 20005 149023 20039 149051
rect 20067 149023 20101 149051
rect 20129 149023 20163 149051
rect 20191 149023 20239 149051
rect 19929 148989 20239 149023
rect 19929 148961 19977 148989
rect 20005 148961 20039 148989
rect 20067 148961 20101 148989
rect 20129 148961 20163 148989
rect 20191 148961 20239 148989
rect 19929 140175 20239 148961
rect 31264 149175 31424 149192
rect 31264 149147 31299 149175
rect 31327 149147 31361 149175
rect 31389 149147 31424 149175
rect 31264 149113 31424 149147
rect 31264 149085 31299 149113
rect 31327 149085 31361 149113
rect 31389 149085 31424 149113
rect 31264 149051 31424 149085
rect 31264 149023 31299 149051
rect 31327 149023 31361 149051
rect 31389 149023 31424 149051
rect 31264 148989 31424 149023
rect 31264 148961 31299 148989
rect 31327 148961 31361 148989
rect 31389 148961 31424 148989
rect 31264 148944 31424 148961
rect 23584 146175 23744 146192
rect 23584 146147 23619 146175
rect 23647 146147 23681 146175
rect 23709 146147 23744 146175
rect 23584 146113 23744 146147
rect 23584 146085 23619 146113
rect 23647 146085 23681 146113
rect 23709 146085 23744 146113
rect 23584 146051 23744 146085
rect 23584 146023 23619 146051
rect 23647 146023 23681 146051
rect 23709 146023 23744 146051
rect 23584 145989 23744 146023
rect 23584 145961 23619 145989
rect 23647 145961 23681 145989
rect 23709 145961 23744 145989
rect 23584 145944 23744 145961
rect 33429 146175 33739 154961
rect 33429 146147 33477 146175
rect 33505 146147 33539 146175
rect 33567 146147 33601 146175
rect 33629 146147 33663 146175
rect 33691 146147 33739 146175
rect 33429 146113 33739 146147
rect 33429 146085 33477 146113
rect 33505 146085 33539 146113
rect 33567 146085 33601 146113
rect 33629 146085 33663 146113
rect 33691 146085 33739 146113
rect 33429 146051 33739 146085
rect 33429 146023 33477 146051
rect 33505 146023 33539 146051
rect 33567 146023 33601 146051
rect 33629 146023 33663 146051
rect 33691 146023 33739 146051
rect 33429 145989 33739 146023
rect 33429 145961 33477 145989
rect 33505 145961 33539 145989
rect 33567 145961 33601 145989
rect 33629 145961 33663 145989
rect 33691 145961 33739 145989
rect 19929 140147 19977 140175
rect 20005 140147 20039 140175
rect 20067 140147 20101 140175
rect 20129 140147 20163 140175
rect 20191 140147 20239 140175
rect 19929 140113 20239 140147
rect 19929 140085 19977 140113
rect 20005 140085 20039 140113
rect 20067 140085 20101 140113
rect 20129 140085 20163 140113
rect 20191 140085 20239 140113
rect 19929 140051 20239 140085
rect 19929 140023 19977 140051
rect 20005 140023 20039 140051
rect 20067 140023 20101 140051
rect 20129 140023 20163 140051
rect 20191 140023 20239 140051
rect 19929 139989 20239 140023
rect 19929 139961 19977 139989
rect 20005 139961 20039 139989
rect 20067 139961 20101 139989
rect 20129 139961 20163 139989
rect 20191 139961 20239 139989
rect 19929 131175 20239 139961
rect 31264 140175 31424 140192
rect 31264 140147 31299 140175
rect 31327 140147 31361 140175
rect 31389 140147 31424 140175
rect 31264 140113 31424 140147
rect 31264 140085 31299 140113
rect 31327 140085 31361 140113
rect 31389 140085 31424 140113
rect 31264 140051 31424 140085
rect 31264 140023 31299 140051
rect 31327 140023 31361 140051
rect 31389 140023 31424 140051
rect 31264 139989 31424 140023
rect 31264 139961 31299 139989
rect 31327 139961 31361 139989
rect 31389 139961 31424 139989
rect 31264 139944 31424 139961
rect 23584 137175 23744 137192
rect 23584 137147 23619 137175
rect 23647 137147 23681 137175
rect 23709 137147 23744 137175
rect 23584 137113 23744 137147
rect 23584 137085 23619 137113
rect 23647 137085 23681 137113
rect 23709 137085 23744 137113
rect 23584 137051 23744 137085
rect 23584 137023 23619 137051
rect 23647 137023 23681 137051
rect 23709 137023 23744 137051
rect 23584 136989 23744 137023
rect 23584 136961 23619 136989
rect 23647 136961 23681 136989
rect 23709 136961 23744 136989
rect 23584 136944 23744 136961
rect 33429 137175 33739 145961
rect 33429 137147 33477 137175
rect 33505 137147 33539 137175
rect 33567 137147 33601 137175
rect 33629 137147 33663 137175
rect 33691 137147 33739 137175
rect 33429 137113 33739 137147
rect 33429 137085 33477 137113
rect 33505 137085 33539 137113
rect 33567 137085 33601 137113
rect 33629 137085 33663 137113
rect 33691 137085 33739 137113
rect 33429 137051 33739 137085
rect 33429 137023 33477 137051
rect 33505 137023 33539 137051
rect 33567 137023 33601 137051
rect 33629 137023 33663 137051
rect 33691 137023 33739 137051
rect 33429 136989 33739 137023
rect 33429 136961 33477 136989
rect 33505 136961 33539 136989
rect 33567 136961 33601 136989
rect 33629 136961 33663 136989
rect 33691 136961 33739 136989
rect 19929 131147 19977 131175
rect 20005 131147 20039 131175
rect 20067 131147 20101 131175
rect 20129 131147 20163 131175
rect 20191 131147 20239 131175
rect 19929 131113 20239 131147
rect 19929 131085 19977 131113
rect 20005 131085 20039 131113
rect 20067 131085 20101 131113
rect 20129 131085 20163 131113
rect 20191 131085 20239 131113
rect 19929 131051 20239 131085
rect 19929 131023 19977 131051
rect 20005 131023 20039 131051
rect 20067 131023 20101 131051
rect 20129 131023 20163 131051
rect 20191 131023 20239 131051
rect 19929 130989 20239 131023
rect 19929 130961 19977 130989
rect 20005 130961 20039 130989
rect 20067 130961 20101 130989
rect 20129 130961 20163 130989
rect 20191 130961 20239 130989
rect 19929 122175 20239 130961
rect 31264 131175 31424 131192
rect 31264 131147 31299 131175
rect 31327 131147 31361 131175
rect 31389 131147 31424 131175
rect 31264 131113 31424 131147
rect 31264 131085 31299 131113
rect 31327 131085 31361 131113
rect 31389 131085 31424 131113
rect 31264 131051 31424 131085
rect 31264 131023 31299 131051
rect 31327 131023 31361 131051
rect 31389 131023 31424 131051
rect 31264 130989 31424 131023
rect 31264 130961 31299 130989
rect 31327 130961 31361 130989
rect 31389 130961 31424 130989
rect 31264 130944 31424 130961
rect 23584 128175 23744 128192
rect 23584 128147 23619 128175
rect 23647 128147 23681 128175
rect 23709 128147 23744 128175
rect 23584 128113 23744 128147
rect 23584 128085 23619 128113
rect 23647 128085 23681 128113
rect 23709 128085 23744 128113
rect 23584 128051 23744 128085
rect 23584 128023 23619 128051
rect 23647 128023 23681 128051
rect 23709 128023 23744 128051
rect 23584 127989 23744 128023
rect 23584 127961 23619 127989
rect 23647 127961 23681 127989
rect 23709 127961 23744 127989
rect 23584 127944 23744 127961
rect 33429 128175 33739 136961
rect 33429 128147 33477 128175
rect 33505 128147 33539 128175
rect 33567 128147 33601 128175
rect 33629 128147 33663 128175
rect 33691 128147 33739 128175
rect 33429 128113 33739 128147
rect 33429 128085 33477 128113
rect 33505 128085 33539 128113
rect 33567 128085 33601 128113
rect 33629 128085 33663 128113
rect 33691 128085 33739 128113
rect 33429 128051 33739 128085
rect 33429 128023 33477 128051
rect 33505 128023 33539 128051
rect 33567 128023 33601 128051
rect 33629 128023 33663 128051
rect 33691 128023 33739 128051
rect 33429 127989 33739 128023
rect 33429 127961 33477 127989
rect 33505 127961 33539 127989
rect 33567 127961 33601 127989
rect 33629 127961 33663 127989
rect 33691 127961 33739 127989
rect 19929 122147 19977 122175
rect 20005 122147 20039 122175
rect 20067 122147 20101 122175
rect 20129 122147 20163 122175
rect 20191 122147 20239 122175
rect 19929 122113 20239 122147
rect 19929 122085 19977 122113
rect 20005 122085 20039 122113
rect 20067 122085 20101 122113
rect 20129 122085 20163 122113
rect 20191 122085 20239 122113
rect 19929 122051 20239 122085
rect 19929 122023 19977 122051
rect 20005 122023 20039 122051
rect 20067 122023 20101 122051
rect 20129 122023 20163 122051
rect 20191 122023 20239 122051
rect 19929 121989 20239 122023
rect 19929 121961 19977 121989
rect 20005 121961 20039 121989
rect 20067 121961 20101 121989
rect 20129 121961 20163 121989
rect 20191 121961 20239 121989
rect 19929 113175 20239 121961
rect 31264 122175 31424 122192
rect 31264 122147 31299 122175
rect 31327 122147 31361 122175
rect 31389 122147 31424 122175
rect 31264 122113 31424 122147
rect 31264 122085 31299 122113
rect 31327 122085 31361 122113
rect 31389 122085 31424 122113
rect 31264 122051 31424 122085
rect 31264 122023 31299 122051
rect 31327 122023 31361 122051
rect 31389 122023 31424 122051
rect 31264 121989 31424 122023
rect 31264 121961 31299 121989
rect 31327 121961 31361 121989
rect 31389 121961 31424 121989
rect 31264 121944 31424 121961
rect 23584 119175 23744 119192
rect 23584 119147 23619 119175
rect 23647 119147 23681 119175
rect 23709 119147 23744 119175
rect 23584 119113 23744 119147
rect 23584 119085 23619 119113
rect 23647 119085 23681 119113
rect 23709 119085 23744 119113
rect 23584 119051 23744 119085
rect 23584 119023 23619 119051
rect 23647 119023 23681 119051
rect 23709 119023 23744 119051
rect 23584 118989 23744 119023
rect 23584 118961 23619 118989
rect 23647 118961 23681 118989
rect 23709 118961 23744 118989
rect 23584 118944 23744 118961
rect 33429 119175 33739 127961
rect 33429 119147 33477 119175
rect 33505 119147 33539 119175
rect 33567 119147 33601 119175
rect 33629 119147 33663 119175
rect 33691 119147 33739 119175
rect 33429 119113 33739 119147
rect 33429 119085 33477 119113
rect 33505 119085 33539 119113
rect 33567 119085 33601 119113
rect 33629 119085 33663 119113
rect 33691 119085 33739 119113
rect 33429 119051 33739 119085
rect 33429 119023 33477 119051
rect 33505 119023 33539 119051
rect 33567 119023 33601 119051
rect 33629 119023 33663 119051
rect 33691 119023 33739 119051
rect 33429 118989 33739 119023
rect 33429 118961 33477 118989
rect 33505 118961 33539 118989
rect 33567 118961 33601 118989
rect 33629 118961 33663 118989
rect 33691 118961 33739 118989
rect 19929 113147 19977 113175
rect 20005 113147 20039 113175
rect 20067 113147 20101 113175
rect 20129 113147 20163 113175
rect 20191 113147 20239 113175
rect 19929 113113 20239 113147
rect 19929 113085 19977 113113
rect 20005 113085 20039 113113
rect 20067 113085 20101 113113
rect 20129 113085 20163 113113
rect 20191 113085 20239 113113
rect 19929 113051 20239 113085
rect 19929 113023 19977 113051
rect 20005 113023 20039 113051
rect 20067 113023 20101 113051
rect 20129 113023 20163 113051
rect 20191 113023 20239 113051
rect 19929 112989 20239 113023
rect 19929 112961 19977 112989
rect 20005 112961 20039 112989
rect 20067 112961 20101 112989
rect 20129 112961 20163 112989
rect 20191 112961 20239 112989
rect 19929 104175 20239 112961
rect 31264 113175 31424 113192
rect 31264 113147 31299 113175
rect 31327 113147 31361 113175
rect 31389 113147 31424 113175
rect 31264 113113 31424 113147
rect 31264 113085 31299 113113
rect 31327 113085 31361 113113
rect 31389 113085 31424 113113
rect 31264 113051 31424 113085
rect 31264 113023 31299 113051
rect 31327 113023 31361 113051
rect 31389 113023 31424 113051
rect 31264 112989 31424 113023
rect 31264 112961 31299 112989
rect 31327 112961 31361 112989
rect 31389 112961 31424 112989
rect 31264 112944 31424 112961
rect 23584 110175 23744 110192
rect 23584 110147 23619 110175
rect 23647 110147 23681 110175
rect 23709 110147 23744 110175
rect 23584 110113 23744 110147
rect 23584 110085 23619 110113
rect 23647 110085 23681 110113
rect 23709 110085 23744 110113
rect 23584 110051 23744 110085
rect 23584 110023 23619 110051
rect 23647 110023 23681 110051
rect 23709 110023 23744 110051
rect 23584 109989 23744 110023
rect 23584 109961 23619 109989
rect 23647 109961 23681 109989
rect 23709 109961 23744 109989
rect 23584 109944 23744 109961
rect 33429 110175 33739 118961
rect 33429 110147 33477 110175
rect 33505 110147 33539 110175
rect 33567 110147 33601 110175
rect 33629 110147 33663 110175
rect 33691 110147 33739 110175
rect 33429 110113 33739 110147
rect 33429 110085 33477 110113
rect 33505 110085 33539 110113
rect 33567 110085 33601 110113
rect 33629 110085 33663 110113
rect 33691 110085 33739 110113
rect 33429 110051 33739 110085
rect 33429 110023 33477 110051
rect 33505 110023 33539 110051
rect 33567 110023 33601 110051
rect 33629 110023 33663 110051
rect 33691 110023 33739 110051
rect 33429 109989 33739 110023
rect 33429 109961 33477 109989
rect 33505 109961 33539 109989
rect 33567 109961 33601 109989
rect 33629 109961 33663 109989
rect 33691 109961 33739 109989
rect 19929 104147 19977 104175
rect 20005 104147 20039 104175
rect 20067 104147 20101 104175
rect 20129 104147 20163 104175
rect 20191 104147 20239 104175
rect 19929 104113 20239 104147
rect 19929 104085 19977 104113
rect 20005 104085 20039 104113
rect 20067 104085 20101 104113
rect 20129 104085 20163 104113
rect 20191 104085 20239 104113
rect 19929 104051 20239 104085
rect 19929 104023 19977 104051
rect 20005 104023 20039 104051
rect 20067 104023 20101 104051
rect 20129 104023 20163 104051
rect 20191 104023 20239 104051
rect 19929 103989 20239 104023
rect 19929 103961 19977 103989
rect 20005 103961 20039 103989
rect 20067 103961 20101 103989
rect 20129 103961 20163 103989
rect 20191 103961 20239 103989
rect 19929 95175 20239 103961
rect 31264 104175 31424 104192
rect 31264 104147 31299 104175
rect 31327 104147 31361 104175
rect 31389 104147 31424 104175
rect 31264 104113 31424 104147
rect 31264 104085 31299 104113
rect 31327 104085 31361 104113
rect 31389 104085 31424 104113
rect 31264 104051 31424 104085
rect 31264 104023 31299 104051
rect 31327 104023 31361 104051
rect 31389 104023 31424 104051
rect 31264 103989 31424 104023
rect 31264 103961 31299 103989
rect 31327 103961 31361 103989
rect 31389 103961 31424 103989
rect 31264 103944 31424 103961
rect 23584 101175 23744 101192
rect 23584 101147 23619 101175
rect 23647 101147 23681 101175
rect 23709 101147 23744 101175
rect 23584 101113 23744 101147
rect 23584 101085 23619 101113
rect 23647 101085 23681 101113
rect 23709 101085 23744 101113
rect 23584 101051 23744 101085
rect 23584 101023 23619 101051
rect 23647 101023 23681 101051
rect 23709 101023 23744 101051
rect 23584 100989 23744 101023
rect 23584 100961 23619 100989
rect 23647 100961 23681 100989
rect 23709 100961 23744 100989
rect 23584 100944 23744 100961
rect 33429 101175 33739 109961
rect 33429 101147 33477 101175
rect 33505 101147 33539 101175
rect 33567 101147 33601 101175
rect 33629 101147 33663 101175
rect 33691 101147 33739 101175
rect 33429 101113 33739 101147
rect 33429 101085 33477 101113
rect 33505 101085 33539 101113
rect 33567 101085 33601 101113
rect 33629 101085 33663 101113
rect 33691 101085 33739 101113
rect 33429 101051 33739 101085
rect 33429 101023 33477 101051
rect 33505 101023 33539 101051
rect 33567 101023 33601 101051
rect 33629 101023 33663 101051
rect 33691 101023 33739 101051
rect 33429 100989 33739 101023
rect 33429 100961 33477 100989
rect 33505 100961 33539 100989
rect 33567 100961 33601 100989
rect 33629 100961 33663 100989
rect 33691 100961 33739 100989
rect 19929 95147 19977 95175
rect 20005 95147 20039 95175
rect 20067 95147 20101 95175
rect 20129 95147 20163 95175
rect 20191 95147 20239 95175
rect 19929 95113 20239 95147
rect 19929 95085 19977 95113
rect 20005 95085 20039 95113
rect 20067 95085 20101 95113
rect 20129 95085 20163 95113
rect 20191 95085 20239 95113
rect 19929 95051 20239 95085
rect 19929 95023 19977 95051
rect 20005 95023 20039 95051
rect 20067 95023 20101 95051
rect 20129 95023 20163 95051
rect 20191 95023 20239 95051
rect 19929 94989 20239 95023
rect 19929 94961 19977 94989
rect 20005 94961 20039 94989
rect 20067 94961 20101 94989
rect 20129 94961 20163 94989
rect 20191 94961 20239 94989
rect 19929 86175 20239 94961
rect 31264 95175 31424 95192
rect 31264 95147 31299 95175
rect 31327 95147 31361 95175
rect 31389 95147 31424 95175
rect 31264 95113 31424 95147
rect 31264 95085 31299 95113
rect 31327 95085 31361 95113
rect 31389 95085 31424 95113
rect 31264 95051 31424 95085
rect 31264 95023 31299 95051
rect 31327 95023 31361 95051
rect 31389 95023 31424 95051
rect 31264 94989 31424 95023
rect 31264 94961 31299 94989
rect 31327 94961 31361 94989
rect 31389 94961 31424 94989
rect 31264 94944 31424 94961
rect 23584 92175 23744 92192
rect 23584 92147 23619 92175
rect 23647 92147 23681 92175
rect 23709 92147 23744 92175
rect 23584 92113 23744 92147
rect 23584 92085 23619 92113
rect 23647 92085 23681 92113
rect 23709 92085 23744 92113
rect 23584 92051 23744 92085
rect 23584 92023 23619 92051
rect 23647 92023 23681 92051
rect 23709 92023 23744 92051
rect 23584 91989 23744 92023
rect 23584 91961 23619 91989
rect 23647 91961 23681 91989
rect 23709 91961 23744 91989
rect 23584 91944 23744 91961
rect 33429 92175 33739 100961
rect 33429 92147 33477 92175
rect 33505 92147 33539 92175
rect 33567 92147 33601 92175
rect 33629 92147 33663 92175
rect 33691 92147 33739 92175
rect 33429 92113 33739 92147
rect 33429 92085 33477 92113
rect 33505 92085 33539 92113
rect 33567 92085 33601 92113
rect 33629 92085 33663 92113
rect 33691 92085 33739 92113
rect 33429 92051 33739 92085
rect 33429 92023 33477 92051
rect 33505 92023 33539 92051
rect 33567 92023 33601 92051
rect 33629 92023 33663 92051
rect 33691 92023 33739 92051
rect 33429 91989 33739 92023
rect 33429 91961 33477 91989
rect 33505 91961 33539 91989
rect 33567 91961 33601 91989
rect 33629 91961 33663 91989
rect 33691 91961 33739 91989
rect 19929 86147 19977 86175
rect 20005 86147 20039 86175
rect 20067 86147 20101 86175
rect 20129 86147 20163 86175
rect 20191 86147 20239 86175
rect 19929 86113 20239 86147
rect 19929 86085 19977 86113
rect 20005 86085 20039 86113
rect 20067 86085 20101 86113
rect 20129 86085 20163 86113
rect 20191 86085 20239 86113
rect 19929 86051 20239 86085
rect 19929 86023 19977 86051
rect 20005 86023 20039 86051
rect 20067 86023 20101 86051
rect 20129 86023 20163 86051
rect 20191 86023 20239 86051
rect 19929 85989 20239 86023
rect 19929 85961 19977 85989
rect 20005 85961 20039 85989
rect 20067 85961 20101 85989
rect 20129 85961 20163 85989
rect 20191 85961 20239 85989
rect 19929 77175 20239 85961
rect 31264 86175 31424 86192
rect 31264 86147 31299 86175
rect 31327 86147 31361 86175
rect 31389 86147 31424 86175
rect 31264 86113 31424 86147
rect 31264 86085 31299 86113
rect 31327 86085 31361 86113
rect 31389 86085 31424 86113
rect 31264 86051 31424 86085
rect 31264 86023 31299 86051
rect 31327 86023 31361 86051
rect 31389 86023 31424 86051
rect 31264 85989 31424 86023
rect 31264 85961 31299 85989
rect 31327 85961 31361 85989
rect 31389 85961 31424 85989
rect 31264 85944 31424 85961
rect 23584 83175 23744 83192
rect 23584 83147 23619 83175
rect 23647 83147 23681 83175
rect 23709 83147 23744 83175
rect 23584 83113 23744 83147
rect 23584 83085 23619 83113
rect 23647 83085 23681 83113
rect 23709 83085 23744 83113
rect 23584 83051 23744 83085
rect 23584 83023 23619 83051
rect 23647 83023 23681 83051
rect 23709 83023 23744 83051
rect 23584 82989 23744 83023
rect 23584 82961 23619 82989
rect 23647 82961 23681 82989
rect 23709 82961 23744 82989
rect 23584 82944 23744 82961
rect 33429 83175 33739 91961
rect 33429 83147 33477 83175
rect 33505 83147 33539 83175
rect 33567 83147 33601 83175
rect 33629 83147 33663 83175
rect 33691 83147 33739 83175
rect 33429 83113 33739 83147
rect 33429 83085 33477 83113
rect 33505 83085 33539 83113
rect 33567 83085 33601 83113
rect 33629 83085 33663 83113
rect 33691 83085 33739 83113
rect 33429 83051 33739 83085
rect 33429 83023 33477 83051
rect 33505 83023 33539 83051
rect 33567 83023 33601 83051
rect 33629 83023 33663 83051
rect 33691 83023 33739 83051
rect 33429 82989 33739 83023
rect 33429 82961 33477 82989
rect 33505 82961 33539 82989
rect 33567 82961 33601 82989
rect 33629 82961 33663 82989
rect 33691 82961 33739 82989
rect 19929 77147 19977 77175
rect 20005 77147 20039 77175
rect 20067 77147 20101 77175
rect 20129 77147 20163 77175
rect 20191 77147 20239 77175
rect 19929 77113 20239 77147
rect 19929 77085 19977 77113
rect 20005 77085 20039 77113
rect 20067 77085 20101 77113
rect 20129 77085 20163 77113
rect 20191 77085 20239 77113
rect 19929 77051 20239 77085
rect 19929 77023 19977 77051
rect 20005 77023 20039 77051
rect 20067 77023 20101 77051
rect 20129 77023 20163 77051
rect 20191 77023 20239 77051
rect 19929 76989 20239 77023
rect 19929 76961 19977 76989
rect 20005 76961 20039 76989
rect 20067 76961 20101 76989
rect 20129 76961 20163 76989
rect 20191 76961 20239 76989
rect 19929 68175 20239 76961
rect 31264 77175 31424 77192
rect 31264 77147 31299 77175
rect 31327 77147 31361 77175
rect 31389 77147 31424 77175
rect 31264 77113 31424 77147
rect 31264 77085 31299 77113
rect 31327 77085 31361 77113
rect 31389 77085 31424 77113
rect 31264 77051 31424 77085
rect 31264 77023 31299 77051
rect 31327 77023 31361 77051
rect 31389 77023 31424 77051
rect 31264 76989 31424 77023
rect 31264 76961 31299 76989
rect 31327 76961 31361 76989
rect 31389 76961 31424 76989
rect 31264 76944 31424 76961
rect 23584 74175 23744 74192
rect 23584 74147 23619 74175
rect 23647 74147 23681 74175
rect 23709 74147 23744 74175
rect 23584 74113 23744 74147
rect 23584 74085 23619 74113
rect 23647 74085 23681 74113
rect 23709 74085 23744 74113
rect 23584 74051 23744 74085
rect 23584 74023 23619 74051
rect 23647 74023 23681 74051
rect 23709 74023 23744 74051
rect 23584 73989 23744 74023
rect 23584 73961 23619 73989
rect 23647 73961 23681 73989
rect 23709 73961 23744 73989
rect 23584 73944 23744 73961
rect 33429 74175 33739 82961
rect 33429 74147 33477 74175
rect 33505 74147 33539 74175
rect 33567 74147 33601 74175
rect 33629 74147 33663 74175
rect 33691 74147 33739 74175
rect 33429 74113 33739 74147
rect 33429 74085 33477 74113
rect 33505 74085 33539 74113
rect 33567 74085 33601 74113
rect 33629 74085 33663 74113
rect 33691 74085 33739 74113
rect 33429 74051 33739 74085
rect 33429 74023 33477 74051
rect 33505 74023 33539 74051
rect 33567 74023 33601 74051
rect 33629 74023 33663 74051
rect 33691 74023 33739 74051
rect 33429 73989 33739 74023
rect 33429 73961 33477 73989
rect 33505 73961 33539 73989
rect 33567 73961 33601 73989
rect 33629 73961 33663 73989
rect 33691 73961 33739 73989
rect 19929 68147 19977 68175
rect 20005 68147 20039 68175
rect 20067 68147 20101 68175
rect 20129 68147 20163 68175
rect 20191 68147 20239 68175
rect 19929 68113 20239 68147
rect 19929 68085 19977 68113
rect 20005 68085 20039 68113
rect 20067 68085 20101 68113
rect 20129 68085 20163 68113
rect 20191 68085 20239 68113
rect 19929 68051 20239 68085
rect 19929 68023 19977 68051
rect 20005 68023 20039 68051
rect 20067 68023 20101 68051
rect 20129 68023 20163 68051
rect 20191 68023 20239 68051
rect 19929 67989 20239 68023
rect 19929 67961 19977 67989
rect 20005 67961 20039 67989
rect 20067 67961 20101 67989
rect 20129 67961 20163 67989
rect 20191 67961 20239 67989
rect 19929 59175 20239 67961
rect 31264 68175 31424 68192
rect 31264 68147 31299 68175
rect 31327 68147 31361 68175
rect 31389 68147 31424 68175
rect 31264 68113 31424 68147
rect 31264 68085 31299 68113
rect 31327 68085 31361 68113
rect 31389 68085 31424 68113
rect 31264 68051 31424 68085
rect 31264 68023 31299 68051
rect 31327 68023 31361 68051
rect 31389 68023 31424 68051
rect 31264 67989 31424 68023
rect 31264 67961 31299 67989
rect 31327 67961 31361 67989
rect 31389 67961 31424 67989
rect 31264 67944 31424 67961
rect 23584 65175 23744 65192
rect 23584 65147 23619 65175
rect 23647 65147 23681 65175
rect 23709 65147 23744 65175
rect 23584 65113 23744 65147
rect 23584 65085 23619 65113
rect 23647 65085 23681 65113
rect 23709 65085 23744 65113
rect 23584 65051 23744 65085
rect 23584 65023 23619 65051
rect 23647 65023 23681 65051
rect 23709 65023 23744 65051
rect 23584 64989 23744 65023
rect 23584 64961 23619 64989
rect 23647 64961 23681 64989
rect 23709 64961 23744 64989
rect 23584 64944 23744 64961
rect 33429 65175 33739 73961
rect 33429 65147 33477 65175
rect 33505 65147 33539 65175
rect 33567 65147 33601 65175
rect 33629 65147 33663 65175
rect 33691 65147 33739 65175
rect 33429 65113 33739 65147
rect 33429 65085 33477 65113
rect 33505 65085 33539 65113
rect 33567 65085 33601 65113
rect 33629 65085 33663 65113
rect 33691 65085 33739 65113
rect 33429 65051 33739 65085
rect 33429 65023 33477 65051
rect 33505 65023 33539 65051
rect 33567 65023 33601 65051
rect 33629 65023 33663 65051
rect 33691 65023 33739 65051
rect 33429 64989 33739 65023
rect 33429 64961 33477 64989
rect 33505 64961 33539 64989
rect 33567 64961 33601 64989
rect 33629 64961 33663 64989
rect 33691 64961 33739 64989
rect 19929 59147 19977 59175
rect 20005 59147 20039 59175
rect 20067 59147 20101 59175
rect 20129 59147 20163 59175
rect 20191 59147 20239 59175
rect 19929 59113 20239 59147
rect 19929 59085 19977 59113
rect 20005 59085 20039 59113
rect 20067 59085 20101 59113
rect 20129 59085 20163 59113
rect 20191 59085 20239 59113
rect 19929 59051 20239 59085
rect 19929 59023 19977 59051
rect 20005 59023 20039 59051
rect 20067 59023 20101 59051
rect 20129 59023 20163 59051
rect 20191 59023 20239 59051
rect 19929 58989 20239 59023
rect 19929 58961 19977 58989
rect 20005 58961 20039 58989
rect 20067 58961 20101 58989
rect 20129 58961 20163 58989
rect 20191 58961 20239 58989
rect 19929 50175 20239 58961
rect 31264 59175 31424 59192
rect 31264 59147 31299 59175
rect 31327 59147 31361 59175
rect 31389 59147 31424 59175
rect 31264 59113 31424 59147
rect 31264 59085 31299 59113
rect 31327 59085 31361 59113
rect 31389 59085 31424 59113
rect 31264 59051 31424 59085
rect 31264 59023 31299 59051
rect 31327 59023 31361 59051
rect 31389 59023 31424 59051
rect 31264 58989 31424 59023
rect 31264 58961 31299 58989
rect 31327 58961 31361 58989
rect 31389 58961 31424 58989
rect 31264 58944 31424 58961
rect 23584 56175 23744 56192
rect 23584 56147 23619 56175
rect 23647 56147 23681 56175
rect 23709 56147 23744 56175
rect 23584 56113 23744 56147
rect 23584 56085 23619 56113
rect 23647 56085 23681 56113
rect 23709 56085 23744 56113
rect 23584 56051 23744 56085
rect 23584 56023 23619 56051
rect 23647 56023 23681 56051
rect 23709 56023 23744 56051
rect 23584 55989 23744 56023
rect 23584 55961 23619 55989
rect 23647 55961 23681 55989
rect 23709 55961 23744 55989
rect 23584 55944 23744 55961
rect 33429 56175 33739 64961
rect 33429 56147 33477 56175
rect 33505 56147 33539 56175
rect 33567 56147 33601 56175
rect 33629 56147 33663 56175
rect 33691 56147 33739 56175
rect 33429 56113 33739 56147
rect 33429 56085 33477 56113
rect 33505 56085 33539 56113
rect 33567 56085 33601 56113
rect 33629 56085 33663 56113
rect 33691 56085 33739 56113
rect 33429 56051 33739 56085
rect 33429 56023 33477 56051
rect 33505 56023 33539 56051
rect 33567 56023 33601 56051
rect 33629 56023 33663 56051
rect 33691 56023 33739 56051
rect 33429 55989 33739 56023
rect 33429 55961 33477 55989
rect 33505 55961 33539 55989
rect 33567 55961 33601 55989
rect 33629 55961 33663 55989
rect 33691 55961 33739 55989
rect 19929 50147 19977 50175
rect 20005 50147 20039 50175
rect 20067 50147 20101 50175
rect 20129 50147 20163 50175
rect 20191 50147 20239 50175
rect 19929 50113 20239 50147
rect 19929 50085 19977 50113
rect 20005 50085 20039 50113
rect 20067 50085 20101 50113
rect 20129 50085 20163 50113
rect 20191 50085 20239 50113
rect 19929 50051 20239 50085
rect 19929 50023 19977 50051
rect 20005 50023 20039 50051
rect 20067 50023 20101 50051
rect 20129 50023 20163 50051
rect 20191 50023 20239 50051
rect 19929 49989 20239 50023
rect 19929 49961 19977 49989
rect 20005 49961 20039 49989
rect 20067 49961 20101 49989
rect 20129 49961 20163 49989
rect 20191 49961 20239 49989
rect 19929 41175 20239 49961
rect 31264 50175 31424 50192
rect 31264 50147 31299 50175
rect 31327 50147 31361 50175
rect 31389 50147 31424 50175
rect 31264 50113 31424 50147
rect 31264 50085 31299 50113
rect 31327 50085 31361 50113
rect 31389 50085 31424 50113
rect 31264 50051 31424 50085
rect 31264 50023 31299 50051
rect 31327 50023 31361 50051
rect 31389 50023 31424 50051
rect 31264 49989 31424 50023
rect 31264 49961 31299 49989
rect 31327 49961 31361 49989
rect 31389 49961 31424 49989
rect 31264 49944 31424 49961
rect 23584 47175 23744 47192
rect 23584 47147 23619 47175
rect 23647 47147 23681 47175
rect 23709 47147 23744 47175
rect 23584 47113 23744 47147
rect 23584 47085 23619 47113
rect 23647 47085 23681 47113
rect 23709 47085 23744 47113
rect 23584 47051 23744 47085
rect 23584 47023 23619 47051
rect 23647 47023 23681 47051
rect 23709 47023 23744 47051
rect 23584 46989 23744 47023
rect 23584 46961 23619 46989
rect 23647 46961 23681 46989
rect 23709 46961 23744 46989
rect 23584 46944 23744 46961
rect 33429 47175 33739 55961
rect 33429 47147 33477 47175
rect 33505 47147 33539 47175
rect 33567 47147 33601 47175
rect 33629 47147 33663 47175
rect 33691 47147 33739 47175
rect 33429 47113 33739 47147
rect 33429 47085 33477 47113
rect 33505 47085 33539 47113
rect 33567 47085 33601 47113
rect 33629 47085 33663 47113
rect 33691 47085 33739 47113
rect 33429 47051 33739 47085
rect 33429 47023 33477 47051
rect 33505 47023 33539 47051
rect 33567 47023 33601 47051
rect 33629 47023 33663 47051
rect 33691 47023 33739 47051
rect 33429 46989 33739 47023
rect 33429 46961 33477 46989
rect 33505 46961 33539 46989
rect 33567 46961 33601 46989
rect 33629 46961 33663 46989
rect 33691 46961 33739 46989
rect 19929 41147 19977 41175
rect 20005 41147 20039 41175
rect 20067 41147 20101 41175
rect 20129 41147 20163 41175
rect 20191 41147 20239 41175
rect 19929 41113 20239 41147
rect 19929 41085 19977 41113
rect 20005 41085 20039 41113
rect 20067 41085 20101 41113
rect 20129 41085 20163 41113
rect 20191 41085 20239 41113
rect 19929 41051 20239 41085
rect 19929 41023 19977 41051
rect 20005 41023 20039 41051
rect 20067 41023 20101 41051
rect 20129 41023 20163 41051
rect 20191 41023 20239 41051
rect 19929 40989 20239 41023
rect 19929 40961 19977 40989
rect 20005 40961 20039 40989
rect 20067 40961 20101 40989
rect 20129 40961 20163 40989
rect 20191 40961 20239 40989
rect 19929 32175 20239 40961
rect 31264 41175 31424 41192
rect 31264 41147 31299 41175
rect 31327 41147 31361 41175
rect 31389 41147 31424 41175
rect 31264 41113 31424 41147
rect 31264 41085 31299 41113
rect 31327 41085 31361 41113
rect 31389 41085 31424 41113
rect 31264 41051 31424 41085
rect 31264 41023 31299 41051
rect 31327 41023 31361 41051
rect 31389 41023 31424 41051
rect 31264 40989 31424 41023
rect 31264 40961 31299 40989
rect 31327 40961 31361 40989
rect 31389 40961 31424 40989
rect 31264 40944 31424 40961
rect 23584 38175 23744 38192
rect 23584 38147 23619 38175
rect 23647 38147 23681 38175
rect 23709 38147 23744 38175
rect 23584 38113 23744 38147
rect 23584 38085 23619 38113
rect 23647 38085 23681 38113
rect 23709 38085 23744 38113
rect 23584 38051 23744 38085
rect 23584 38023 23619 38051
rect 23647 38023 23681 38051
rect 23709 38023 23744 38051
rect 23584 37989 23744 38023
rect 23584 37961 23619 37989
rect 23647 37961 23681 37989
rect 23709 37961 23744 37989
rect 23584 37944 23744 37961
rect 33429 38175 33739 46961
rect 33429 38147 33477 38175
rect 33505 38147 33539 38175
rect 33567 38147 33601 38175
rect 33629 38147 33663 38175
rect 33691 38147 33739 38175
rect 33429 38113 33739 38147
rect 33429 38085 33477 38113
rect 33505 38085 33539 38113
rect 33567 38085 33601 38113
rect 33629 38085 33663 38113
rect 33691 38085 33739 38113
rect 33429 38051 33739 38085
rect 33429 38023 33477 38051
rect 33505 38023 33539 38051
rect 33567 38023 33601 38051
rect 33629 38023 33663 38051
rect 33691 38023 33739 38051
rect 33429 37989 33739 38023
rect 33429 37961 33477 37989
rect 33505 37961 33539 37989
rect 33567 37961 33601 37989
rect 33629 37961 33663 37989
rect 33691 37961 33739 37989
rect 19929 32147 19977 32175
rect 20005 32147 20039 32175
rect 20067 32147 20101 32175
rect 20129 32147 20163 32175
rect 20191 32147 20239 32175
rect 19929 32113 20239 32147
rect 19929 32085 19977 32113
rect 20005 32085 20039 32113
rect 20067 32085 20101 32113
rect 20129 32085 20163 32113
rect 20191 32085 20239 32113
rect 19929 32051 20239 32085
rect 19929 32023 19977 32051
rect 20005 32023 20039 32051
rect 20067 32023 20101 32051
rect 20129 32023 20163 32051
rect 20191 32023 20239 32051
rect 19929 31989 20239 32023
rect 19929 31961 19977 31989
rect 20005 31961 20039 31989
rect 20067 31961 20101 31989
rect 20129 31961 20163 31989
rect 20191 31961 20239 31989
rect 19929 23175 20239 31961
rect 31264 32175 31424 32192
rect 31264 32147 31299 32175
rect 31327 32147 31361 32175
rect 31389 32147 31424 32175
rect 31264 32113 31424 32147
rect 31264 32085 31299 32113
rect 31327 32085 31361 32113
rect 31389 32085 31424 32113
rect 31264 32051 31424 32085
rect 31264 32023 31299 32051
rect 31327 32023 31361 32051
rect 31389 32023 31424 32051
rect 31264 31989 31424 32023
rect 31264 31961 31299 31989
rect 31327 31961 31361 31989
rect 31389 31961 31424 31989
rect 31264 31944 31424 31961
rect 23584 29175 23744 29192
rect 23584 29147 23619 29175
rect 23647 29147 23681 29175
rect 23709 29147 23744 29175
rect 23584 29113 23744 29147
rect 23584 29085 23619 29113
rect 23647 29085 23681 29113
rect 23709 29085 23744 29113
rect 23584 29051 23744 29085
rect 23584 29023 23619 29051
rect 23647 29023 23681 29051
rect 23709 29023 23744 29051
rect 23584 28989 23744 29023
rect 23584 28961 23619 28989
rect 23647 28961 23681 28989
rect 23709 28961 23744 28989
rect 23584 28944 23744 28961
rect 33429 29175 33739 37961
rect 33429 29147 33477 29175
rect 33505 29147 33539 29175
rect 33567 29147 33601 29175
rect 33629 29147 33663 29175
rect 33691 29147 33739 29175
rect 33429 29113 33739 29147
rect 33429 29085 33477 29113
rect 33505 29085 33539 29113
rect 33567 29085 33601 29113
rect 33629 29085 33663 29113
rect 33691 29085 33739 29113
rect 33429 29051 33739 29085
rect 33429 29023 33477 29051
rect 33505 29023 33539 29051
rect 33567 29023 33601 29051
rect 33629 29023 33663 29051
rect 33691 29023 33739 29051
rect 33429 28989 33739 29023
rect 33429 28961 33477 28989
rect 33505 28961 33539 28989
rect 33567 28961 33601 28989
rect 33629 28961 33663 28989
rect 33691 28961 33739 28989
rect 19929 23147 19977 23175
rect 20005 23147 20039 23175
rect 20067 23147 20101 23175
rect 20129 23147 20163 23175
rect 20191 23147 20239 23175
rect 19929 23113 20239 23147
rect 19929 23085 19977 23113
rect 20005 23085 20039 23113
rect 20067 23085 20101 23113
rect 20129 23085 20163 23113
rect 20191 23085 20239 23113
rect 19929 23051 20239 23085
rect 19929 23023 19977 23051
rect 20005 23023 20039 23051
rect 20067 23023 20101 23051
rect 20129 23023 20163 23051
rect 20191 23023 20239 23051
rect 19929 22989 20239 23023
rect 19929 22961 19977 22989
rect 20005 22961 20039 22989
rect 20067 22961 20101 22989
rect 20129 22961 20163 22989
rect 20191 22961 20239 22989
rect 19929 14175 20239 22961
rect 31264 23175 31424 23192
rect 31264 23147 31299 23175
rect 31327 23147 31361 23175
rect 31389 23147 31424 23175
rect 31264 23113 31424 23147
rect 31264 23085 31299 23113
rect 31327 23085 31361 23113
rect 31389 23085 31424 23113
rect 31264 23051 31424 23085
rect 31264 23023 31299 23051
rect 31327 23023 31361 23051
rect 31389 23023 31424 23051
rect 31264 22989 31424 23023
rect 31264 22961 31299 22989
rect 31327 22961 31361 22989
rect 31389 22961 31424 22989
rect 31264 22944 31424 22961
rect 23584 20175 23744 20192
rect 23584 20147 23619 20175
rect 23647 20147 23681 20175
rect 23709 20147 23744 20175
rect 23584 20113 23744 20147
rect 23584 20085 23619 20113
rect 23647 20085 23681 20113
rect 23709 20085 23744 20113
rect 23584 20051 23744 20085
rect 23584 20023 23619 20051
rect 23647 20023 23681 20051
rect 23709 20023 23744 20051
rect 23584 19989 23744 20023
rect 23584 19961 23619 19989
rect 23647 19961 23681 19989
rect 23709 19961 23744 19989
rect 23584 19944 23744 19961
rect 33429 20175 33739 28961
rect 33429 20147 33477 20175
rect 33505 20147 33539 20175
rect 33567 20147 33601 20175
rect 33629 20147 33663 20175
rect 33691 20147 33739 20175
rect 33429 20113 33739 20147
rect 33429 20085 33477 20113
rect 33505 20085 33539 20113
rect 33567 20085 33601 20113
rect 33629 20085 33663 20113
rect 33691 20085 33739 20113
rect 33429 20051 33739 20085
rect 33429 20023 33477 20051
rect 33505 20023 33539 20051
rect 33567 20023 33601 20051
rect 33629 20023 33663 20051
rect 33691 20023 33739 20051
rect 33429 19989 33739 20023
rect 33429 19961 33477 19989
rect 33505 19961 33539 19989
rect 33567 19961 33601 19989
rect 33629 19961 33663 19989
rect 33691 19961 33739 19989
rect 19929 14147 19977 14175
rect 20005 14147 20039 14175
rect 20067 14147 20101 14175
rect 20129 14147 20163 14175
rect 20191 14147 20239 14175
rect 19929 14113 20239 14147
rect 19929 14085 19977 14113
rect 20005 14085 20039 14113
rect 20067 14085 20101 14113
rect 20129 14085 20163 14113
rect 20191 14085 20239 14113
rect 19929 14051 20239 14085
rect 19929 14023 19977 14051
rect 20005 14023 20039 14051
rect 20067 14023 20101 14051
rect 20129 14023 20163 14051
rect 20191 14023 20239 14051
rect 19929 13989 20239 14023
rect 19929 13961 19977 13989
rect 20005 13961 20039 13989
rect 20067 13961 20101 13989
rect 20129 13961 20163 13989
rect 20191 13961 20239 13989
rect 19929 5175 20239 13961
rect 31264 14175 31424 14192
rect 31264 14147 31299 14175
rect 31327 14147 31361 14175
rect 31389 14147 31424 14175
rect 31264 14113 31424 14147
rect 31264 14085 31299 14113
rect 31327 14085 31361 14113
rect 31389 14085 31424 14113
rect 31264 14051 31424 14085
rect 31264 14023 31299 14051
rect 31327 14023 31361 14051
rect 31389 14023 31424 14051
rect 31264 13989 31424 14023
rect 31264 13961 31299 13989
rect 31327 13961 31361 13989
rect 31389 13961 31424 13989
rect 31264 13944 31424 13961
rect 23584 11175 23744 11192
rect 23584 11147 23619 11175
rect 23647 11147 23681 11175
rect 23709 11147 23744 11175
rect 23584 11113 23744 11147
rect 23584 11085 23619 11113
rect 23647 11085 23681 11113
rect 23709 11085 23744 11113
rect 23584 11051 23744 11085
rect 23584 11023 23619 11051
rect 23647 11023 23681 11051
rect 23709 11023 23744 11051
rect 23584 10989 23744 11023
rect 23584 10961 23619 10989
rect 23647 10961 23681 10989
rect 23709 10961 23744 10989
rect 23584 10944 23744 10961
rect 33429 11175 33739 19961
rect 33429 11147 33477 11175
rect 33505 11147 33539 11175
rect 33567 11147 33601 11175
rect 33629 11147 33663 11175
rect 33691 11147 33739 11175
rect 33429 11113 33739 11147
rect 33429 11085 33477 11113
rect 33505 11085 33539 11113
rect 33567 11085 33601 11113
rect 33629 11085 33663 11113
rect 33691 11085 33739 11113
rect 33429 11051 33739 11085
rect 33429 11023 33477 11051
rect 33505 11023 33539 11051
rect 33567 11023 33601 11051
rect 33629 11023 33663 11051
rect 33691 11023 33739 11051
rect 33429 10989 33739 11023
rect 33429 10961 33477 10989
rect 33505 10961 33539 10989
rect 33567 10961 33601 10989
rect 33629 10961 33663 10989
rect 33691 10961 33739 10989
rect 19929 5147 19977 5175
rect 20005 5147 20039 5175
rect 20067 5147 20101 5175
rect 20129 5147 20163 5175
rect 20191 5147 20239 5175
rect 19929 5113 20239 5147
rect 19929 5085 19977 5113
rect 20005 5085 20039 5113
rect 20067 5085 20101 5113
rect 20129 5085 20163 5113
rect 20191 5085 20239 5113
rect 19929 5051 20239 5085
rect 19929 5023 19977 5051
rect 20005 5023 20039 5051
rect 20067 5023 20101 5051
rect 20129 5023 20163 5051
rect 20191 5023 20239 5051
rect 19929 4989 20239 5023
rect 19929 4961 19977 4989
rect 20005 4961 20039 4989
rect 20067 4961 20101 4989
rect 20129 4961 20163 4989
rect 20191 4961 20239 4989
rect 19929 -560 20239 4961
rect 31264 5175 31424 5192
rect 31264 5147 31299 5175
rect 31327 5147 31361 5175
rect 31389 5147 31424 5175
rect 31264 5113 31424 5147
rect 31264 5085 31299 5113
rect 31327 5085 31361 5113
rect 31389 5085 31424 5113
rect 31264 5051 31424 5085
rect 31264 5023 31299 5051
rect 31327 5023 31361 5051
rect 31389 5023 31424 5051
rect 31264 4989 31424 5023
rect 31264 4961 31299 4989
rect 31327 4961 31361 4989
rect 31389 4961 31424 4989
rect 31264 4944 31424 4961
rect 19929 -588 19977 -560
rect 20005 -588 20039 -560
rect 20067 -588 20101 -560
rect 20129 -588 20163 -560
rect 20191 -588 20239 -560
rect 19929 -622 20239 -588
rect 19929 -650 19977 -622
rect 20005 -650 20039 -622
rect 20067 -650 20101 -622
rect 20129 -650 20163 -622
rect 20191 -650 20239 -622
rect 19929 -684 20239 -650
rect 19929 -712 19977 -684
rect 20005 -712 20039 -684
rect 20067 -712 20101 -684
rect 20129 -712 20163 -684
rect 20191 -712 20239 -684
rect 19929 -746 20239 -712
rect 19929 -774 19977 -746
rect 20005 -774 20039 -746
rect 20067 -774 20101 -746
rect 20129 -774 20163 -746
rect 20191 -774 20239 -746
rect 19929 -822 20239 -774
rect 33429 2175 33739 10961
rect 33429 2147 33477 2175
rect 33505 2147 33539 2175
rect 33567 2147 33601 2175
rect 33629 2147 33663 2175
rect 33691 2147 33739 2175
rect 33429 2113 33739 2147
rect 33429 2085 33477 2113
rect 33505 2085 33539 2113
rect 33567 2085 33601 2113
rect 33629 2085 33663 2113
rect 33691 2085 33739 2113
rect 33429 2051 33739 2085
rect 33429 2023 33477 2051
rect 33505 2023 33539 2051
rect 33567 2023 33601 2051
rect 33629 2023 33663 2051
rect 33691 2023 33739 2051
rect 33429 1989 33739 2023
rect 33429 1961 33477 1989
rect 33505 1961 33539 1989
rect 33567 1961 33601 1989
rect 33629 1961 33663 1989
rect 33691 1961 33739 1989
rect 33429 -80 33739 1961
rect 33429 -108 33477 -80
rect 33505 -108 33539 -80
rect 33567 -108 33601 -80
rect 33629 -108 33663 -80
rect 33691 -108 33739 -80
rect 33429 -142 33739 -108
rect 33429 -170 33477 -142
rect 33505 -170 33539 -142
rect 33567 -170 33601 -142
rect 33629 -170 33663 -142
rect 33691 -170 33739 -142
rect 33429 -204 33739 -170
rect 33429 -232 33477 -204
rect 33505 -232 33539 -204
rect 33567 -232 33601 -204
rect 33629 -232 33663 -204
rect 33691 -232 33739 -204
rect 33429 -266 33739 -232
rect 33429 -294 33477 -266
rect 33505 -294 33539 -266
rect 33567 -294 33601 -266
rect 33629 -294 33663 -266
rect 33691 -294 33739 -266
rect 33429 -822 33739 -294
rect 35289 299086 35599 299134
rect 35289 299058 35337 299086
rect 35365 299058 35399 299086
rect 35427 299058 35461 299086
rect 35489 299058 35523 299086
rect 35551 299058 35599 299086
rect 35289 299024 35599 299058
rect 35289 298996 35337 299024
rect 35365 298996 35399 299024
rect 35427 298996 35461 299024
rect 35489 298996 35523 299024
rect 35551 298996 35599 299024
rect 35289 298962 35599 298996
rect 35289 298934 35337 298962
rect 35365 298934 35399 298962
rect 35427 298934 35461 298962
rect 35489 298934 35523 298962
rect 35551 298934 35599 298962
rect 35289 298900 35599 298934
rect 35289 298872 35337 298900
rect 35365 298872 35399 298900
rect 35427 298872 35461 298900
rect 35489 298872 35523 298900
rect 35551 298872 35599 298900
rect 35289 293175 35599 298872
rect 35289 293147 35337 293175
rect 35365 293147 35399 293175
rect 35427 293147 35461 293175
rect 35489 293147 35523 293175
rect 35551 293147 35599 293175
rect 35289 293113 35599 293147
rect 35289 293085 35337 293113
rect 35365 293085 35399 293113
rect 35427 293085 35461 293113
rect 35489 293085 35523 293113
rect 35551 293085 35599 293113
rect 35289 293051 35599 293085
rect 35289 293023 35337 293051
rect 35365 293023 35399 293051
rect 35427 293023 35461 293051
rect 35489 293023 35523 293051
rect 35551 293023 35599 293051
rect 35289 292989 35599 293023
rect 35289 292961 35337 292989
rect 35365 292961 35399 292989
rect 35427 292961 35461 292989
rect 35489 292961 35523 292989
rect 35551 292961 35599 292989
rect 35289 284175 35599 292961
rect 35289 284147 35337 284175
rect 35365 284147 35399 284175
rect 35427 284147 35461 284175
rect 35489 284147 35523 284175
rect 35551 284147 35599 284175
rect 35289 284113 35599 284147
rect 35289 284085 35337 284113
rect 35365 284085 35399 284113
rect 35427 284085 35461 284113
rect 35489 284085 35523 284113
rect 35551 284085 35599 284113
rect 35289 284051 35599 284085
rect 35289 284023 35337 284051
rect 35365 284023 35399 284051
rect 35427 284023 35461 284051
rect 35489 284023 35523 284051
rect 35551 284023 35599 284051
rect 35289 283989 35599 284023
rect 35289 283961 35337 283989
rect 35365 283961 35399 283989
rect 35427 283961 35461 283989
rect 35489 283961 35523 283989
rect 35551 283961 35599 283989
rect 35289 275175 35599 283961
rect 35289 275147 35337 275175
rect 35365 275147 35399 275175
rect 35427 275147 35461 275175
rect 35489 275147 35523 275175
rect 35551 275147 35599 275175
rect 35289 275113 35599 275147
rect 35289 275085 35337 275113
rect 35365 275085 35399 275113
rect 35427 275085 35461 275113
rect 35489 275085 35523 275113
rect 35551 275085 35599 275113
rect 35289 275051 35599 275085
rect 35289 275023 35337 275051
rect 35365 275023 35399 275051
rect 35427 275023 35461 275051
rect 35489 275023 35523 275051
rect 35551 275023 35599 275051
rect 35289 274989 35599 275023
rect 35289 274961 35337 274989
rect 35365 274961 35399 274989
rect 35427 274961 35461 274989
rect 35489 274961 35523 274989
rect 35551 274961 35599 274989
rect 35289 266175 35599 274961
rect 35289 266147 35337 266175
rect 35365 266147 35399 266175
rect 35427 266147 35461 266175
rect 35489 266147 35523 266175
rect 35551 266147 35599 266175
rect 35289 266113 35599 266147
rect 35289 266085 35337 266113
rect 35365 266085 35399 266113
rect 35427 266085 35461 266113
rect 35489 266085 35523 266113
rect 35551 266085 35599 266113
rect 35289 266051 35599 266085
rect 35289 266023 35337 266051
rect 35365 266023 35399 266051
rect 35427 266023 35461 266051
rect 35489 266023 35523 266051
rect 35551 266023 35599 266051
rect 35289 265989 35599 266023
rect 35289 265961 35337 265989
rect 35365 265961 35399 265989
rect 35427 265961 35461 265989
rect 35489 265961 35523 265989
rect 35551 265961 35599 265989
rect 35289 257175 35599 265961
rect 35289 257147 35337 257175
rect 35365 257147 35399 257175
rect 35427 257147 35461 257175
rect 35489 257147 35523 257175
rect 35551 257147 35599 257175
rect 35289 257113 35599 257147
rect 35289 257085 35337 257113
rect 35365 257085 35399 257113
rect 35427 257085 35461 257113
rect 35489 257085 35523 257113
rect 35551 257085 35599 257113
rect 35289 257051 35599 257085
rect 35289 257023 35337 257051
rect 35365 257023 35399 257051
rect 35427 257023 35461 257051
rect 35489 257023 35523 257051
rect 35551 257023 35599 257051
rect 35289 256989 35599 257023
rect 35289 256961 35337 256989
rect 35365 256961 35399 256989
rect 35427 256961 35461 256989
rect 35489 256961 35523 256989
rect 35551 256961 35599 256989
rect 35289 248175 35599 256961
rect 35289 248147 35337 248175
rect 35365 248147 35399 248175
rect 35427 248147 35461 248175
rect 35489 248147 35523 248175
rect 35551 248147 35599 248175
rect 35289 248113 35599 248147
rect 35289 248085 35337 248113
rect 35365 248085 35399 248113
rect 35427 248085 35461 248113
rect 35489 248085 35523 248113
rect 35551 248085 35599 248113
rect 35289 248051 35599 248085
rect 35289 248023 35337 248051
rect 35365 248023 35399 248051
rect 35427 248023 35461 248051
rect 35489 248023 35523 248051
rect 35551 248023 35599 248051
rect 35289 247989 35599 248023
rect 35289 247961 35337 247989
rect 35365 247961 35399 247989
rect 35427 247961 35461 247989
rect 35489 247961 35523 247989
rect 35551 247961 35599 247989
rect 35289 239175 35599 247961
rect 35289 239147 35337 239175
rect 35365 239147 35399 239175
rect 35427 239147 35461 239175
rect 35489 239147 35523 239175
rect 35551 239147 35599 239175
rect 35289 239113 35599 239147
rect 35289 239085 35337 239113
rect 35365 239085 35399 239113
rect 35427 239085 35461 239113
rect 35489 239085 35523 239113
rect 35551 239085 35599 239113
rect 35289 239051 35599 239085
rect 35289 239023 35337 239051
rect 35365 239023 35399 239051
rect 35427 239023 35461 239051
rect 35489 239023 35523 239051
rect 35551 239023 35599 239051
rect 35289 238989 35599 239023
rect 35289 238961 35337 238989
rect 35365 238961 35399 238989
rect 35427 238961 35461 238989
rect 35489 238961 35523 238989
rect 35551 238961 35599 238989
rect 35289 230175 35599 238961
rect 35289 230147 35337 230175
rect 35365 230147 35399 230175
rect 35427 230147 35461 230175
rect 35489 230147 35523 230175
rect 35551 230147 35599 230175
rect 35289 230113 35599 230147
rect 35289 230085 35337 230113
rect 35365 230085 35399 230113
rect 35427 230085 35461 230113
rect 35489 230085 35523 230113
rect 35551 230085 35599 230113
rect 35289 230051 35599 230085
rect 35289 230023 35337 230051
rect 35365 230023 35399 230051
rect 35427 230023 35461 230051
rect 35489 230023 35523 230051
rect 35551 230023 35599 230051
rect 35289 229989 35599 230023
rect 35289 229961 35337 229989
rect 35365 229961 35399 229989
rect 35427 229961 35461 229989
rect 35489 229961 35523 229989
rect 35551 229961 35599 229989
rect 35289 221175 35599 229961
rect 35289 221147 35337 221175
rect 35365 221147 35399 221175
rect 35427 221147 35461 221175
rect 35489 221147 35523 221175
rect 35551 221147 35599 221175
rect 35289 221113 35599 221147
rect 35289 221085 35337 221113
rect 35365 221085 35399 221113
rect 35427 221085 35461 221113
rect 35489 221085 35523 221113
rect 35551 221085 35599 221113
rect 35289 221051 35599 221085
rect 35289 221023 35337 221051
rect 35365 221023 35399 221051
rect 35427 221023 35461 221051
rect 35489 221023 35523 221051
rect 35551 221023 35599 221051
rect 35289 220989 35599 221023
rect 35289 220961 35337 220989
rect 35365 220961 35399 220989
rect 35427 220961 35461 220989
rect 35489 220961 35523 220989
rect 35551 220961 35599 220989
rect 35289 212175 35599 220961
rect 35289 212147 35337 212175
rect 35365 212147 35399 212175
rect 35427 212147 35461 212175
rect 35489 212147 35523 212175
rect 35551 212147 35599 212175
rect 35289 212113 35599 212147
rect 35289 212085 35337 212113
rect 35365 212085 35399 212113
rect 35427 212085 35461 212113
rect 35489 212085 35523 212113
rect 35551 212085 35599 212113
rect 35289 212051 35599 212085
rect 35289 212023 35337 212051
rect 35365 212023 35399 212051
rect 35427 212023 35461 212051
rect 35489 212023 35523 212051
rect 35551 212023 35599 212051
rect 35289 211989 35599 212023
rect 35289 211961 35337 211989
rect 35365 211961 35399 211989
rect 35427 211961 35461 211989
rect 35489 211961 35523 211989
rect 35551 211961 35599 211989
rect 35289 203175 35599 211961
rect 35289 203147 35337 203175
rect 35365 203147 35399 203175
rect 35427 203147 35461 203175
rect 35489 203147 35523 203175
rect 35551 203147 35599 203175
rect 35289 203113 35599 203147
rect 35289 203085 35337 203113
rect 35365 203085 35399 203113
rect 35427 203085 35461 203113
rect 35489 203085 35523 203113
rect 35551 203085 35599 203113
rect 35289 203051 35599 203085
rect 35289 203023 35337 203051
rect 35365 203023 35399 203051
rect 35427 203023 35461 203051
rect 35489 203023 35523 203051
rect 35551 203023 35599 203051
rect 35289 202989 35599 203023
rect 35289 202961 35337 202989
rect 35365 202961 35399 202989
rect 35427 202961 35461 202989
rect 35489 202961 35523 202989
rect 35551 202961 35599 202989
rect 35289 194175 35599 202961
rect 35289 194147 35337 194175
rect 35365 194147 35399 194175
rect 35427 194147 35461 194175
rect 35489 194147 35523 194175
rect 35551 194147 35599 194175
rect 35289 194113 35599 194147
rect 35289 194085 35337 194113
rect 35365 194085 35399 194113
rect 35427 194085 35461 194113
rect 35489 194085 35523 194113
rect 35551 194085 35599 194113
rect 35289 194051 35599 194085
rect 35289 194023 35337 194051
rect 35365 194023 35399 194051
rect 35427 194023 35461 194051
rect 35489 194023 35523 194051
rect 35551 194023 35599 194051
rect 35289 193989 35599 194023
rect 35289 193961 35337 193989
rect 35365 193961 35399 193989
rect 35427 193961 35461 193989
rect 35489 193961 35523 193989
rect 35551 193961 35599 193989
rect 35289 185175 35599 193961
rect 35289 185147 35337 185175
rect 35365 185147 35399 185175
rect 35427 185147 35461 185175
rect 35489 185147 35523 185175
rect 35551 185147 35599 185175
rect 35289 185113 35599 185147
rect 35289 185085 35337 185113
rect 35365 185085 35399 185113
rect 35427 185085 35461 185113
rect 35489 185085 35523 185113
rect 35551 185085 35599 185113
rect 35289 185051 35599 185085
rect 35289 185023 35337 185051
rect 35365 185023 35399 185051
rect 35427 185023 35461 185051
rect 35489 185023 35523 185051
rect 35551 185023 35599 185051
rect 35289 184989 35599 185023
rect 35289 184961 35337 184989
rect 35365 184961 35399 184989
rect 35427 184961 35461 184989
rect 35489 184961 35523 184989
rect 35551 184961 35599 184989
rect 35289 176175 35599 184961
rect 35289 176147 35337 176175
rect 35365 176147 35399 176175
rect 35427 176147 35461 176175
rect 35489 176147 35523 176175
rect 35551 176147 35599 176175
rect 35289 176113 35599 176147
rect 35289 176085 35337 176113
rect 35365 176085 35399 176113
rect 35427 176085 35461 176113
rect 35489 176085 35523 176113
rect 35551 176085 35599 176113
rect 35289 176051 35599 176085
rect 35289 176023 35337 176051
rect 35365 176023 35399 176051
rect 35427 176023 35461 176051
rect 35489 176023 35523 176051
rect 35551 176023 35599 176051
rect 35289 175989 35599 176023
rect 35289 175961 35337 175989
rect 35365 175961 35399 175989
rect 35427 175961 35461 175989
rect 35489 175961 35523 175989
rect 35551 175961 35599 175989
rect 35289 167175 35599 175961
rect 48789 298606 49099 299134
rect 48789 298578 48837 298606
rect 48865 298578 48899 298606
rect 48927 298578 48961 298606
rect 48989 298578 49023 298606
rect 49051 298578 49099 298606
rect 48789 298544 49099 298578
rect 48789 298516 48837 298544
rect 48865 298516 48899 298544
rect 48927 298516 48961 298544
rect 48989 298516 49023 298544
rect 49051 298516 49099 298544
rect 48789 298482 49099 298516
rect 48789 298454 48837 298482
rect 48865 298454 48899 298482
rect 48927 298454 48961 298482
rect 48989 298454 49023 298482
rect 49051 298454 49099 298482
rect 48789 298420 49099 298454
rect 48789 298392 48837 298420
rect 48865 298392 48899 298420
rect 48927 298392 48961 298420
rect 48989 298392 49023 298420
rect 49051 298392 49099 298420
rect 48789 290175 49099 298392
rect 48789 290147 48837 290175
rect 48865 290147 48899 290175
rect 48927 290147 48961 290175
rect 48989 290147 49023 290175
rect 49051 290147 49099 290175
rect 48789 290113 49099 290147
rect 48789 290085 48837 290113
rect 48865 290085 48899 290113
rect 48927 290085 48961 290113
rect 48989 290085 49023 290113
rect 49051 290085 49099 290113
rect 48789 290051 49099 290085
rect 48789 290023 48837 290051
rect 48865 290023 48899 290051
rect 48927 290023 48961 290051
rect 48989 290023 49023 290051
rect 49051 290023 49099 290051
rect 48789 289989 49099 290023
rect 48789 289961 48837 289989
rect 48865 289961 48899 289989
rect 48927 289961 48961 289989
rect 48989 289961 49023 289989
rect 49051 289961 49099 289989
rect 48789 281175 49099 289961
rect 48789 281147 48837 281175
rect 48865 281147 48899 281175
rect 48927 281147 48961 281175
rect 48989 281147 49023 281175
rect 49051 281147 49099 281175
rect 48789 281113 49099 281147
rect 48789 281085 48837 281113
rect 48865 281085 48899 281113
rect 48927 281085 48961 281113
rect 48989 281085 49023 281113
rect 49051 281085 49099 281113
rect 48789 281051 49099 281085
rect 48789 281023 48837 281051
rect 48865 281023 48899 281051
rect 48927 281023 48961 281051
rect 48989 281023 49023 281051
rect 49051 281023 49099 281051
rect 48789 280989 49099 281023
rect 48789 280961 48837 280989
rect 48865 280961 48899 280989
rect 48927 280961 48961 280989
rect 48989 280961 49023 280989
rect 49051 280961 49099 280989
rect 48789 272175 49099 280961
rect 48789 272147 48837 272175
rect 48865 272147 48899 272175
rect 48927 272147 48961 272175
rect 48989 272147 49023 272175
rect 49051 272147 49099 272175
rect 48789 272113 49099 272147
rect 48789 272085 48837 272113
rect 48865 272085 48899 272113
rect 48927 272085 48961 272113
rect 48989 272085 49023 272113
rect 49051 272085 49099 272113
rect 48789 272051 49099 272085
rect 48789 272023 48837 272051
rect 48865 272023 48899 272051
rect 48927 272023 48961 272051
rect 48989 272023 49023 272051
rect 49051 272023 49099 272051
rect 48789 271989 49099 272023
rect 48789 271961 48837 271989
rect 48865 271961 48899 271989
rect 48927 271961 48961 271989
rect 48989 271961 49023 271989
rect 49051 271961 49099 271989
rect 48789 263175 49099 271961
rect 48789 263147 48837 263175
rect 48865 263147 48899 263175
rect 48927 263147 48961 263175
rect 48989 263147 49023 263175
rect 49051 263147 49099 263175
rect 48789 263113 49099 263147
rect 48789 263085 48837 263113
rect 48865 263085 48899 263113
rect 48927 263085 48961 263113
rect 48989 263085 49023 263113
rect 49051 263085 49099 263113
rect 48789 263051 49099 263085
rect 48789 263023 48837 263051
rect 48865 263023 48899 263051
rect 48927 263023 48961 263051
rect 48989 263023 49023 263051
rect 49051 263023 49099 263051
rect 48789 262989 49099 263023
rect 48789 262961 48837 262989
rect 48865 262961 48899 262989
rect 48927 262961 48961 262989
rect 48989 262961 49023 262989
rect 49051 262961 49099 262989
rect 48789 254175 49099 262961
rect 48789 254147 48837 254175
rect 48865 254147 48899 254175
rect 48927 254147 48961 254175
rect 48989 254147 49023 254175
rect 49051 254147 49099 254175
rect 48789 254113 49099 254147
rect 48789 254085 48837 254113
rect 48865 254085 48899 254113
rect 48927 254085 48961 254113
rect 48989 254085 49023 254113
rect 49051 254085 49099 254113
rect 48789 254051 49099 254085
rect 48789 254023 48837 254051
rect 48865 254023 48899 254051
rect 48927 254023 48961 254051
rect 48989 254023 49023 254051
rect 49051 254023 49099 254051
rect 48789 253989 49099 254023
rect 48789 253961 48837 253989
rect 48865 253961 48899 253989
rect 48927 253961 48961 253989
rect 48989 253961 49023 253989
rect 49051 253961 49099 253989
rect 48789 245175 49099 253961
rect 48789 245147 48837 245175
rect 48865 245147 48899 245175
rect 48927 245147 48961 245175
rect 48989 245147 49023 245175
rect 49051 245147 49099 245175
rect 48789 245113 49099 245147
rect 48789 245085 48837 245113
rect 48865 245085 48899 245113
rect 48927 245085 48961 245113
rect 48989 245085 49023 245113
rect 49051 245085 49099 245113
rect 48789 245051 49099 245085
rect 48789 245023 48837 245051
rect 48865 245023 48899 245051
rect 48927 245023 48961 245051
rect 48989 245023 49023 245051
rect 49051 245023 49099 245051
rect 48789 244989 49099 245023
rect 48789 244961 48837 244989
rect 48865 244961 48899 244989
rect 48927 244961 48961 244989
rect 48989 244961 49023 244989
rect 49051 244961 49099 244989
rect 48789 236175 49099 244961
rect 48789 236147 48837 236175
rect 48865 236147 48899 236175
rect 48927 236147 48961 236175
rect 48989 236147 49023 236175
rect 49051 236147 49099 236175
rect 48789 236113 49099 236147
rect 48789 236085 48837 236113
rect 48865 236085 48899 236113
rect 48927 236085 48961 236113
rect 48989 236085 49023 236113
rect 49051 236085 49099 236113
rect 48789 236051 49099 236085
rect 48789 236023 48837 236051
rect 48865 236023 48899 236051
rect 48927 236023 48961 236051
rect 48989 236023 49023 236051
rect 49051 236023 49099 236051
rect 48789 235989 49099 236023
rect 48789 235961 48837 235989
rect 48865 235961 48899 235989
rect 48927 235961 48961 235989
rect 48989 235961 49023 235989
rect 49051 235961 49099 235989
rect 48789 227175 49099 235961
rect 48789 227147 48837 227175
rect 48865 227147 48899 227175
rect 48927 227147 48961 227175
rect 48989 227147 49023 227175
rect 49051 227147 49099 227175
rect 48789 227113 49099 227147
rect 48789 227085 48837 227113
rect 48865 227085 48899 227113
rect 48927 227085 48961 227113
rect 48989 227085 49023 227113
rect 49051 227085 49099 227113
rect 48789 227051 49099 227085
rect 48789 227023 48837 227051
rect 48865 227023 48899 227051
rect 48927 227023 48961 227051
rect 48989 227023 49023 227051
rect 49051 227023 49099 227051
rect 48789 226989 49099 227023
rect 48789 226961 48837 226989
rect 48865 226961 48899 226989
rect 48927 226961 48961 226989
rect 48989 226961 49023 226989
rect 49051 226961 49099 226989
rect 48789 218175 49099 226961
rect 48789 218147 48837 218175
rect 48865 218147 48899 218175
rect 48927 218147 48961 218175
rect 48989 218147 49023 218175
rect 49051 218147 49099 218175
rect 48789 218113 49099 218147
rect 48789 218085 48837 218113
rect 48865 218085 48899 218113
rect 48927 218085 48961 218113
rect 48989 218085 49023 218113
rect 49051 218085 49099 218113
rect 48789 218051 49099 218085
rect 48789 218023 48837 218051
rect 48865 218023 48899 218051
rect 48927 218023 48961 218051
rect 48989 218023 49023 218051
rect 49051 218023 49099 218051
rect 48789 217989 49099 218023
rect 48789 217961 48837 217989
rect 48865 217961 48899 217989
rect 48927 217961 48961 217989
rect 48989 217961 49023 217989
rect 49051 217961 49099 217989
rect 48789 209175 49099 217961
rect 48789 209147 48837 209175
rect 48865 209147 48899 209175
rect 48927 209147 48961 209175
rect 48989 209147 49023 209175
rect 49051 209147 49099 209175
rect 48789 209113 49099 209147
rect 48789 209085 48837 209113
rect 48865 209085 48899 209113
rect 48927 209085 48961 209113
rect 48989 209085 49023 209113
rect 49051 209085 49099 209113
rect 48789 209051 49099 209085
rect 48789 209023 48837 209051
rect 48865 209023 48899 209051
rect 48927 209023 48961 209051
rect 48989 209023 49023 209051
rect 49051 209023 49099 209051
rect 48789 208989 49099 209023
rect 48789 208961 48837 208989
rect 48865 208961 48899 208989
rect 48927 208961 48961 208989
rect 48989 208961 49023 208989
rect 49051 208961 49099 208989
rect 48789 200175 49099 208961
rect 48789 200147 48837 200175
rect 48865 200147 48899 200175
rect 48927 200147 48961 200175
rect 48989 200147 49023 200175
rect 49051 200147 49099 200175
rect 48789 200113 49099 200147
rect 48789 200085 48837 200113
rect 48865 200085 48899 200113
rect 48927 200085 48961 200113
rect 48989 200085 49023 200113
rect 49051 200085 49099 200113
rect 48789 200051 49099 200085
rect 48789 200023 48837 200051
rect 48865 200023 48899 200051
rect 48927 200023 48961 200051
rect 48989 200023 49023 200051
rect 49051 200023 49099 200051
rect 48789 199989 49099 200023
rect 48789 199961 48837 199989
rect 48865 199961 48899 199989
rect 48927 199961 48961 199989
rect 48989 199961 49023 199989
rect 49051 199961 49099 199989
rect 48789 191175 49099 199961
rect 48789 191147 48837 191175
rect 48865 191147 48899 191175
rect 48927 191147 48961 191175
rect 48989 191147 49023 191175
rect 49051 191147 49099 191175
rect 48789 191113 49099 191147
rect 48789 191085 48837 191113
rect 48865 191085 48899 191113
rect 48927 191085 48961 191113
rect 48989 191085 49023 191113
rect 49051 191085 49099 191113
rect 48789 191051 49099 191085
rect 48789 191023 48837 191051
rect 48865 191023 48899 191051
rect 48927 191023 48961 191051
rect 48989 191023 49023 191051
rect 49051 191023 49099 191051
rect 48789 190989 49099 191023
rect 48789 190961 48837 190989
rect 48865 190961 48899 190989
rect 48927 190961 48961 190989
rect 48989 190961 49023 190989
rect 49051 190961 49099 190989
rect 48789 182175 49099 190961
rect 48789 182147 48837 182175
rect 48865 182147 48899 182175
rect 48927 182147 48961 182175
rect 48989 182147 49023 182175
rect 49051 182147 49099 182175
rect 48789 182113 49099 182147
rect 48789 182085 48837 182113
rect 48865 182085 48899 182113
rect 48927 182085 48961 182113
rect 48989 182085 49023 182113
rect 49051 182085 49099 182113
rect 48789 182051 49099 182085
rect 48789 182023 48837 182051
rect 48865 182023 48899 182051
rect 48927 182023 48961 182051
rect 48989 182023 49023 182051
rect 49051 182023 49099 182051
rect 48789 181989 49099 182023
rect 48789 181961 48837 181989
rect 48865 181961 48899 181989
rect 48927 181961 48961 181989
rect 48989 181961 49023 181989
rect 49051 181961 49099 181989
rect 38944 173175 39104 173192
rect 38944 173147 38979 173175
rect 39007 173147 39041 173175
rect 39069 173147 39104 173175
rect 38944 173113 39104 173147
rect 38944 173085 38979 173113
rect 39007 173085 39041 173113
rect 39069 173085 39104 173113
rect 38944 173051 39104 173085
rect 38944 173023 38979 173051
rect 39007 173023 39041 173051
rect 39069 173023 39104 173051
rect 38944 172989 39104 173023
rect 38944 172961 38979 172989
rect 39007 172961 39041 172989
rect 39069 172961 39104 172989
rect 38944 172944 39104 172961
rect 48789 173175 49099 181961
rect 48789 173147 48837 173175
rect 48865 173147 48899 173175
rect 48927 173147 48961 173175
rect 48989 173147 49023 173175
rect 49051 173147 49099 173175
rect 48789 173113 49099 173147
rect 48789 173085 48837 173113
rect 48865 173085 48899 173113
rect 48927 173085 48961 173113
rect 48989 173085 49023 173113
rect 49051 173085 49099 173113
rect 48789 173051 49099 173085
rect 48789 173023 48837 173051
rect 48865 173023 48899 173051
rect 48927 173023 48961 173051
rect 48989 173023 49023 173051
rect 49051 173023 49099 173051
rect 48789 172989 49099 173023
rect 48789 172961 48837 172989
rect 48865 172961 48899 172989
rect 48927 172961 48961 172989
rect 48989 172961 49023 172989
rect 49051 172961 49099 172989
rect 35289 167147 35337 167175
rect 35365 167147 35399 167175
rect 35427 167147 35461 167175
rect 35489 167147 35523 167175
rect 35551 167147 35599 167175
rect 35289 167113 35599 167147
rect 35289 167085 35337 167113
rect 35365 167085 35399 167113
rect 35427 167085 35461 167113
rect 35489 167085 35523 167113
rect 35551 167085 35599 167113
rect 35289 167051 35599 167085
rect 35289 167023 35337 167051
rect 35365 167023 35399 167051
rect 35427 167023 35461 167051
rect 35489 167023 35523 167051
rect 35551 167023 35599 167051
rect 35289 166989 35599 167023
rect 35289 166961 35337 166989
rect 35365 166961 35399 166989
rect 35427 166961 35461 166989
rect 35489 166961 35523 166989
rect 35551 166961 35599 166989
rect 35289 158175 35599 166961
rect 46624 167175 46784 167192
rect 46624 167147 46659 167175
rect 46687 167147 46721 167175
rect 46749 167147 46784 167175
rect 46624 167113 46784 167147
rect 46624 167085 46659 167113
rect 46687 167085 46721 167113
rect 46749 167085 46784 167113
rect 46624 167051 46784 167085
rect 46624 167023 46659 167051
rect 46687 167023 46721 167051
rect 46749 167023 46784 167051
rect 46624 166989 46784 167023
rect 46624 166961 46659 166989
rect 46687 166961 46721 166989
rect 46749 166961 46784 166989
rect 46624 166944 46784 166961
rect 38944 164175 39104 164192
rect 38944 164147 38979 164175
rect 39007 164147 39041 164175
rect 39069 164147 39104 164175
rect 38944 164113 39104 164147
rect 38944 164085 38979 164113
rect 39007 164085 39041 164113
rect 39069 164085 39104 164113
rect 38944 164051 39104 164085
rect 38944 164023 38979 164051
rect 39007 164023 39041 164051
rect 39069 164023 39104 164051
rect 38944 163989 39104 164023
rect 38944 163961 38979 163989
rect 39007 163961 39041 163989
rect 39069 163961 39104 163989
rect 38944 163944 39104 163961
rect 48789 164175 49099 172961
rect 48789 164147 48837 164175
rect 48865 164147 48899 164175
rect 48927 164147 48961 164175
rect 48989 164147 49023 164175
rect 49051 164147 49099 164175
rect 48789 164113 49099 164147
rect 48789 164085 48837 164113
rect 48865 164085 48899 164113
rect 48927 164085 48961 164113
rect 48989 164085 49023 164113
rect 49051 164085 49099 164113
rect 48789 164051 49099 164085
rect 48789 164023 48837 164051
rect 48865 164023 48899 164051
rect 48927 164023 48961 164051
rect 48989 164023 49023 164051
rect 49051 164023 49099 164051
rect 48789 163989 49099 164023
rect 48789 163961 48837 163989
rect 48865 163961 48899 163989
rect 48927 163961 48961 163989
rect 48989 163961 49023 163989
rect 49051 163961 49099 163989
rect 35289 158147 35337 158175
rect 35365 158147 35399 158175
rect 35427 158147 35461 158175
rect 35489 158147 35523 158175
rect 35551 158147 35599 158175
rect 35289 158113 35599 158147
rect 35289 158085 35337 158113
rect 35365 158085 35399 158113
rect 35427 158085 35461 158113
rect 35489 158085 35523 158113
rect 35551 158085 35599 158113
rect 35289 158051 35599 158085
rect 35289 158023 35337 158051
rect 35365 158023 35399 158051
rect 35427 158023 35461 158051
rect 35489 158023 35523 158051
rect 35551 158023 35599 158051
rect 35289 157989 35599 158023
rect 35289 157961 35337 157989
rect 35365 157961 35399 157989
rect 35427 157961 35461 157989
rect 35489 157961 35523 157989
rect 35551 157961 35599 157989
rect 35289 149175 35599 157961
rect 46624 158175 46784 158192
rect 46624 158147 46659 158175
rect 46687 158147 46721 158175
rect 46749 158147 46784 158175
rect 46624 158113 46784 158147
rect 46624 158085 46659 158113
rect 46687 158085 46721 158113
rect 46749 158085 46784 158113
rect 46624 158051 46784 158085
rect 46624 158023 46659 158051
rect 46687 158023 46721 158051
rect 46749 158023 46784 158051
rect 46624 157989 46784 158023
rect 46624 157961 46659 157989
rect 46687 157961 46721 157989
rect 46749 157961 46784 157989
rect 46624 157944 46784 157961
rect 38944 155175 39104 155192
rect 38944 155147 38979 155175
rect 39007 155147 39041 155175
rect 39069 155147 39104 155175
rect 38944 155113 39104 155147
rect 38944 155085 38979 155113
rect 39007 155085 39041 155113
rect 39069 155085 39104 155113
rect 38944 155051 39104 155085
rect 38944 155023 38979 155051
rect 39007 155023 39041 155051
rect 39069 155023 39104 155051
rect 38944 154989 39104 155023
rect 38944 154961 38979 154989
rect 39007 154961 39041 154989
rect 39069 154961 39104 154989
rect 38944 154944 39104 154961
rect 48789 155175 49099 163961
rect 48789 155147 48837 155175
rect 48865 155147 48899 155175
rect 48927 155147 48961 155175
rect 48989 155147 49023 155175
rect 49051 155147 49099 155175
rect 48789 155113 49099 155147
rect 48789 155085 48837 155113
rect 48865 155085 48899 155113
rect 48927 155085 48961 155113
rect 48989 155085 49023 155113
rect 49051 155085 49099 155113
rect 48789 155051 49099 155085
rect 48789 155023 48837 155051
rect 48865 155023 48899 155051
rect 48927 155023 48961 155051
rect 48989 155023 49023 155051
rect 49051 155023 49099 155051
rect 48789 154989 49099 155023
rect 48789 154961 48837 154989
rect 48865 154961 48899 154989
rect 48927 154961 48961 154989
rect 48989 154961 49023 154989
rect 49051 154961 49099 154989
rect 35289 149147 35337 149175
rect 35365 149147 35399 149175
rect 35427 149147 35461 149175
rect 35489 149147 35523 149175
rect 35551 149147 35599 149175
rect 35289 149113 35599 149147
rect 35289 149085 35337 149113
rect 35365 149085 35399 149113
rect 35427 149085 35461 149113
rect 35489 149085 35523 149113
rect 35551 149085 35599 149113
rect 35289 149051 35599 149085
rect 35289 149023 35337 149051
rect 35365 149023 35399 149051
rect 35427 149023 35461 149051
rect 35489 149023 35523 149051
rect 35551 149023 35599 149051
rect 35289 148989 35599 149023
rect 35289 148961 35337 148989
rect 35365 148961 35399 148989
rect 35427 148961 35461 148989
rect 35489 148961 35523 148989
rect 35551 148961 35599 148989
rect 35289 140175 35599 148961
rect 46624 149175 46784 149192
rect 46624 149147 46659 149175
rect 46687 149147 46721 149175
rect 46749 149147 46784 149175
rect 46624 149113 46784 149147
rect 46624 149085 46659 149113
rect 46687 149085 46721 149113
rect 46749 149085 46784 149113
rect 46624 149051 46784 149085
rect 46624 149023 46659 149051
rect 46687 149023 46721 149051
rect 46749 149023 46784 149051
rect 46624 148989 46784 149023
rect 46624 148961 46659 148989
rect 46687 148961 46721 148989
rect 46749 148961 46784 148989
rect 46624 148944 46784 148961
rect 38944 146175 39104 146192
rect 38944 146147 38979 146175
rect 39007 146147 39041 146175
rect 39069 146147 39104 146175
rect 38944 146113 39104 146147
rect 38944 146085 38979 146113
rect 39007 146085 39041 146113
rect 39069 146085 39104 146113
rect 38944 146051 39104 146085
rect 38944 146023 38979 146051
rect 39007 146023 39041 146051
rect 39069 146023 39104 146051
rect 38944 145989 39104 146023
rect 38944 145961 38979 145989
rect 39007 145961 39041 145989
rect 39069 145961 39104 145989
rect 38944 145944 39104 145961
rect 48789 146175 49099 154961
rect 48789 146147 48837 146175
rect 48865 146147 48899 146175
rect 48927 146147 48961 146175
rect 48989 146147 49023 146175
rect 49051 146147 49099 146175
rect 48789 146113 49099 146147
rect 48789 146085 48837 146113
rect 48865 146085 48899 146113
rect 48927 146085 48961 146113
rect 48989 146085 49023 146113
rect 49051 146085 49099 146113
rect 48789 146051 49099 146085
rect 48789 146023 48837 146051
rect 48865 146023 48899 146051
rect 48927 146023 48961 146051
rect 48989 146023 49023 146051
rect 49051 146023 49099 146051
rect 48789 145989 49099 146023
rect 48789 145961 48837 145989
rect 48865 145961 48899 145989
rect 48927 145961 48961 145989
rect 48989 145961 49023 145989
rect 49051 145961 49099 145989
rect 35289 140147 35337 140175
rect 35365 140147 35399 140175
rect 35427 140147 35461 140175
rect 35489 140147 35523 140175
rect 35551 140147 35599 140175
rect 35289 140113 35599 140147
rect 35289 140085 35337 140113
rect 35365 140085 35399 140113
rect 35427 140085 35461 140113
rect 35489 140085 35523 140113
rect 35551 140085 35599 140113
rect 35289 140051 35599 140085
rect 35289 140023 35337 140051
rect 35365 140023 35399 140051
rect 35427 140023 35461 140051
rect 35489 140023 35523 140051
rect 35551 140023 35599 140051
rect 35289 139989 35599 140023
rect 35289 139961 35337 139989
rect 35365 139961 35399 139989
rect 35427 139961 35461 139989
rect 35489 139961 35523 139989
rect 35551 139961 35599 139989
rect 35289 131175 35599 139961
rect 46624 140175 46784 140192
rect 46624 140147 46659 140175
rect 46687 140147 46721 140175
rect 46749 140147 46784 140175
rect 46624 140113 46784 140147
rect 46624 140085 46659 140113
rect 46687 140085 46721 140113
rect 46749 140085 46784 140113
rect 46624 140051 46784 140085
rect 46624 140023 46659 140051
rect 46687 140023 46721 140051
rect 46749 140023 46784 140051
rect 46624 139989 46784 140023
rect 46624 139961 46659 139989
rect 46687 139961 46721 139989
rect 46749 139961 46784 139989
rect 46624 139944 46784 139961
rect 38944 137175 39104 137192
rect 38944 137147 38979 137175
rect 39007 137147 39041 137175
rect 39069 137147 39104 137175
rect 38944 137113 39104 137147
rect 38944 137085 38979 137113
rect 39007 137085 39041 137113
rect 39069 137085 39104 137113
rect 38944 137051 39104 137085
rect 38944 137023 38979 137051
rect 39007 137023 39041 137051
rect 39069 137023 39104 137051
rect 38944 136989 39104 137023
rect 38944 136961 38979 136989
rect 39007 136961 39041 136989
rect 39069 136961 39104 136989
rect 38944 136944 39104 136961
rect 48789 137175 49099 145961
rect 48789 137147 48837 137175
rect 48865 137147 48899 137175
rect 48927 137147 48961 137175
rect 48989 137147 49023 137175
rect 49051 137147 49099 137175
rect 48789 137113 49099 137147
rect 48789 137085 48837 137113
rect 48865 137085 48899 137113
rect 48927 137085 48961 137113
rect 48989 137085 49023 137113
rect 49051 137085 49099 137113
rect 48789 137051 49099 137085
rect 48789 137023 48837 137051
rect 48865 137023 48899 137051
rect 48927 137023 48961 137051
rect 48989 137023 49023 137051
rect 49051 137023 49099 137051
rect 48789 136989 49099 137023
rect 48789 136961 48837 136989
rect 48865 136961 48899 136989
rect 48927 136961 48961 136989
rect 48989 136961 49023 136989
rect 49051 136961 49099 136989
rect 35289 131147 35337 131175
rect 35365 131147 35399 131175
rect 35427 131147 35461 131175
rect 35489 131147 35523 131175
rect 35551 131147 35599 131175
rect 35289 131113 35599 131147
rect 35289 131085 35337 131113
rect 35365 131085 35399 131113
rect 35427 131085 35461 131113
rect 35489 131085 35523 131113
rect 35551 131085 35599 131113
rect 35289 131051 35599 131085
rect 35289 131023 35337 131051
rect 35365 131023 35399 131051
rect 35427 131023 35461 131051
rect 35489 131023 35523 131051
rect 35551 131023 35599 131051
rect 35289 130989 35599 131023
rect 35289 130961 35337 130989
rect 35365 130961 35399 130989
rect 35427 130961 35461 130989
rect 35489 130961 35523 130989
rect 35551 130961 35599 130989
rect 35289 122175 35599 130961
rect 46624 131175 46784 131192
rect 46624 131147 46659 131175
rect 46687 131147 46721 131175
rect 46749 131147 46784 131175
rect 46624 131113 46784 131147
rect 46624 131085 46659 131113
rect 46687 131085 46721 131113
rect 46749 131085 46784 131113
rect 46624 131051 46784 131085
rect 46624 131023 46659 131051
rect 46687 131023 46721 131051
rect 46749 131023 46784 131051
rect 46624 130989 46784 131023
rect 46624 130961 46659 130989
rect 46687 130961 46721 130989
rect 46749 130961 46784 130989
rect 46624 130944 46784 130961
rect 38944 128175 39104 128192
rect 38944 128147 38979 128175
rect 39007 128147 39041 128175
rect 39069 128147 39104 128175
rect 38944 128113 39104 128147
rect 38944 128085 38979 128113
rect 39007 128085 39041 128113
rect 39069 128085 39104 128113
rect 38944 128051 39104 128085
rect 38944 128023 38979 128051
rect 39007 128023 39041 128051
rect 39069 128023 39104 128051
rect 38944 127989 39104 128023
rect 38944 127961 38979 127989
rect 39007 127961 39041 127989
rect 39069 127961 39104 127989
rect 38944 127944 39104 127961
rect 48789 128175 49099 136961
rect 48789 128147 48837 128175
rect 48865 128147 48899 128175
rect 48927 128147 48961 128175
rect 48989 128147 49023 128175
rect 49051 128147 49099 128175
rect 48789 128113 49099 128147
rect 48789 128085 48837 128113
rect 48865 128085 48899 128113
rect 48927 128085 48961 128113
rect 48989 128085 49023 128113
rect 49051 128085 49099 128113
rect 48789 128051 49099 128085
rect 48789 128023 48837 128051
rect 48865 128023 48899 128051
rect 48927 128023 48961 128051
rect 48989 128023 49023 128051
rect 49051 128023 49099 128051
rect 48789 127989 49099 128023
rect 48789 127961 48837 127989
rect 48865 127961 48899 127989
rect 48927 127961 48961 127989
rect 48989 127961 49023 127989
rect 49051 127961 49099 127989
rect 35289 122147 35337 122175
rect 35365 122147 35399 122175
rect 35427 122147 35461 122175
rect 35489 122147 35523 122175
rect 35551 122147 35599 122175
rect 35289 122113 35599 122147
rect 35289 122085 35337 122113
rect 35365 122085 35399 122113
rect 35427 122085 35461 122113
rect 35489 122085 35523 122113
rect 35551 122085 35599 122113
rect 35289 122051 35599 122085
rect 35289 122023 35337 122051
rect 35365 122023 35399 122051
rect 35427 122023 35461 122051
rect 35489 122023 35523 122051
rect 35551 122023 35599 122051
rect 35289 121989 35599 122023
rect 35289 121961 35337 121989
rect 35365 121961 35399 121989
rect 35427 121961 35461 121989
rect 35489 121961 35523 121989
rect 35551 121961 35599 121989
rect 35289 113175 35599 121961
rect 46624 122175 46784 122192
rect 46624 122147 46659 122175
rect 46687 122147 46721 122175
rect 46749 122147 46784 122175
rect 46624 122113 46784 122147
rect 46624 122085 46659 122113
rect 46687 122085 46721 122113
rect 46749 122085 46784 122113
rect 46624 122051 46784 122085
rect 46624 122023 46659 122051
rect 46687 122023 46721 122051
rect 46749 122023 46784 122051
rect 46624 121989 46784 122023
rect 46624 121961 46659 121989
rect 46687 121961 46721 121989
rect 46749 121961 46784 121989
rect 46624 121944 46784 121961
rect 38944 119175 39104 119192
rect 38944 119147 38979 119175
rect 39007 119147 39041 119175
rect 39069 119147 39104 119175
rect 38944 119113 39104 119147
rect 38944 119085 38979 119113
rect 39007 119085 39041 119113
rect 39069 119085 39104 119113
rect 38944 119051 39104 119085
rect 38944 119023 38979 119051
rect 39007 119023 39041 119051
rect 39069 119023 39104 119051
rect 38944 118989 39104 119023
rect 38944 118961 38979 118989
rect 39007 118961 39041 118989
rect 39069 118961 39104 118989
rect 38944 118944 39104 118961
rect 48789 119175 49099 127961
rect 48789 119147 48837 119175
rect 48865 119147 48899 119175
rect 48927 119147 48961 119175
rect 48989 119147 49023 119175
rect 49051 119147 49099 119175
rect 48789 119113 49099 119147
rect 48789 119085 48837 119113
rect 48865 119085 48899 119113
rect 48927 119085 48961 119113
rect 48989 119085 49023 119113
rect 49051 119085 49099 119113
rect 48789 119051 49099 119085
rect 48789 119023 48837 119051
rect 48865 119023 48899 119051
rect 48927 119023 48961 119051
rect 48989 119023 49023 119051
rect 49051 119023 49099 119051
rect 48789 118989 49099 119023
rect 48789 118961 48837 118989
rect 48865 118961 48899 118989
rect 48927 118961 48961 118989
rect 48989 118961 49023 118989
rect 49051 118961 49099 118989
rect 35289 113147 35337 113175
rect 35365 113147 35399 113175
rect 35427 113147 35461 113175
rect 35489 113147 35523 113175
rect 35551 113147 35599 113175
rect 35289 113113 35599 113147
rect 35289 113085 35337 113113
rect 35365 113085 35399 113113
rect 35427 113085 35461 113113
rect 35489 113085 35523 113113
rect 35551 113085 35599 113113
rect 35289 113051 35599 113085
rect 35289 113023 35337 113051
rect 35365 113023 35399 113051
rect 35427 113023 35461 113051
rect 35489 113023 35523 113051
rect 35551 113023 35599 113051
rect 35289 112989 35599 113023
rect 35289 112961 35337 112989
rect 35365 112961 35399 112989
rect 35427 112961 35461 112989
rect 35489 112961 35523 112989
rect 35551 112961 35599 112989
rect 35289 104175 35599 112961
rect 46624 113175 46784 113192
rect 46624 113147 46659 113175
rect 46687 113147 46721 113175
rect 46749 113147 46784 113175
rect 46624 113113 46784 113147
rect 46624 113085 46659 113113
rect 46687 113085 46721 113113
rect 46749 113085 46784 113113
rect 46624 113051 46784 113085
rect 46624 113023 46659 113051
rect 46687 113023 46721 113051
rect 46749 113023 46784 113051
rect 46624 112989 46784 113023
rect 46624 112961 46659 112989
rect 46687 112961 46721 112989
rect 46749 112961 46784 112989
rect 46624 112944 46784 112961
rect 38944 110175 39104 110192
rect 38944 110147 38979 110175
rect 39007 110147 39041 110175
rect 39069 110147 39104 110175
rect 38944 110113 39104 110147
rect 38944 110085 38979 110113
rect 39007 110085 39041 110113
rect 39069 110085 39104 110113
rect 38944 110051 39104 110085
rect 38944 110023 38979 110051
rect 39007 110023 39041 110051
rect 39069 110023 39104 110051
rect 38944 109989 39104 110023
rect 38944 109961 38979 109989
rect 39007 109961 39041 109989
rect 39069 109961 39104 109989
rect 38944 109944 39104 109961
rect 48789 110175 49099 118961
rect 48789 110147 48837 110175
rect 48865 110147 48899 110175
rect 48927 110147 48961 110175
rect 48989 110147 49023 110175
rect 49051 110147 49099 110175
rect 48789 110113 49099 110147
rect 48789 110085 48837 110113
rect 48865 110085 48899 110113
rect 48927 110085 48961 110113
rect 48989 110085 49023 110113
rect 49051 110085 49099 110113
rect 48789 110051 49099 110085
rect 48789 110023 48837 110051
rect 48865 110023 48899 110051
rect 48927 110023 48961 110051
rect 48989 110023 49023 110051
rect 49051 110023 49099 110051
rect 48789 109989 49099 110023
rect 48789 109961 48837 109989
rect 48865 109961 48899 109989
rect 48927 109961 48961 109989
rect 48989 109961 49023 109989
rect 49051 109961 49099 109989
rect 35289 104147 35337 104175
rect 35365 104147 35399 104175
rect 35427 104147 35461 104175
rect 35489 104147 35523 104175
rect 35551 104147 35599 104175
rect 35289 104113 35599 104147
rect 35289 104085 35337 104113
rect 35365 104085 35399 104113
rect 35427 104085 35461 104113
rect 35489 104085 35523 104113
rect 35551 104085 35599 104113
rect 35289 104051 35599 104085
rect 35289 104023 35337 104051
rect 35365 104023 35399 104051
rect 35427 104023 35461 104051
rect 35489 104023 35523 104051
rect 35551 104023 35599 104051
rect 35289 103989 35599 104023
rect 35289 103961 35337 103989
rect 35365 103961 35399 103989
rect 35427 103961 35461 103989
rect 35489 103961 35523 103989
rect 35551 103961 35599 103989
rect 35289 95175 35599 103961
rect 46624 104175 46784 104192
rect 46624 104147 46659 104175
rect 46687 104147 46721 104175
rect 46749 104147 46784 104175
rect 46624 104113 46784 104147
rect 46624 104085 46659 104113
rect 46687 104085 46721 104113
rect 46749 104085 46784 104113
rect 46624 104051 46784 104085
rect 46624 104023 46659 104051
rect 46687 104023 46721 104051
rect 46749 104023 46784 104051
rect 46624 103989 46784 104023
rect 46624 103961 46659 103989
rect 46687 103961 46721 103989
rect 46749 103961 46784 103989
rect 46624 103944 46784 103961
rect 38944 101175 39104 101192
rect 38944 101147 38979 101175
rect 39007 101147 39041 101175
rect 39069 101147 39104 101175
rect 38944 101113 39104 101147
rect 38944 101085 38979 101113
rect 39007 101085 39041 101113
rect 39069 101085 39104 101113
rect 38944 101051 39104 101085
rect 38944 101023 38979 101051
rect 39007 101023 39041 101051
rect 39069 101023 39104 101051
rect 38944 100989 39104 101023
rect 38944 100961 38979 100989
rect 39007 100961 39041 100989
rect 39069 100961 39104 100989
rect 38944 100944 39104 100961
rect 48789 101175 49099 109961
rect 48789 101147 48837 101175
rect 48865 101147 48899 101175
rect 48927 101147 48961 101175
rect 48989 101147 49023 101175
rect 49051 101147 49099 101175
rect 48789 101113 49099 101147
rect 48789 101085 48837 101113
rect 48865 101085 48899 101113
rect 48927 101085 48961 101113
rect 48989 101085 49023 101113
rect 49051 101085 49099 101113
rect 48789 101051 49099 101085
rect 48789 101023 48837 101051
rect 48865 101023 48899 101051
rect 48927 101023 48961 101051
rect 48989 101023 49023 101051
rect 49051 101023 49099 101051
rect 48789 100989 49099 101023
rect 48789 100961 48837 100989
rect 48865 100961 48899 100989
rect 48927 100961 48961 100989
rect 48989 100961 49023 100989
rect 49051 100961 49099 100989
rect 35289 95147 35337 95175
rect 35365 95147 35399 95175
rect 35427 95147 35461 95175
rect 35489 95147 35523 95175
rect 35551 95147 35599 95175
rect 35289 95113 35599 95147
rect 35289 95085 35337 95113
rect 35365 95085 35399 95113
rect 35427 95085 35461 95113
rect 35489 95085 35523 95113
rect 35551 95085 35599 95113
rect 35289 95051 35599 95085
rect 35289 95023 35337 95051
rect 35365 95023 35399 95051
rect 35427 95023 35461 95051
rect 35489 95023 35523 95051
rect 35551 95023 35599 95051
rect 35289 94989 35599 95023
rect 35289 94961 35337 94989
rect 35365 94961 35399 94989
rect 35427 94961 35461 94989
rect 35489 94961 35523 94989
rect 35551 94961 35599 94989
rect 35289 86175 35599 94961
rect 46624 95175 46784 95192
rect 46624 95147 46659 95175
rect 46687 95147 46721 95175
rect 46749 95147 46784 95175
rect 46624 95113 46784 95147
rect 46624 95085 46659 95113
rect 46687 95085 46721 95113
rect 46749 95085 46784 95113
rect 46624 95051 46784 95085
rect 46624 95023 46659 95051
rect 46687 95023 46721 95051
rect 46749 95023 46784 95051
rect 46624 94989 46784 95023
rect 46624 94961 46659 94989
rect 46687 94961 46721 94989
rect 46749 94961 46784 94989
rect 46624 94944 46784 94961
rect 38944 92175 39104 92192
rect 38944 92147 38979 92175
rect 39007 92147 39041 92175
rect 39069 92147 39104 92175
rect 38944 92113 39104 92147
rect 38944 92085 38979 92113
rect 39007 92085 39041 92113
rect 39069 92085 39104 92113
rect 38944 92051 39104 92085
rect 38944 92023 38979 92051
rect 39007 92023 39041 92051
rect 39069 92023 39104 92051
rect 38944 91989 39104 92023
rect 38944 91961 38979 91989
rect 39007 91961 39041 91989
rect 39069 91961 39104 91989
rect 38944 91944 39104 91961
rect 48789 92175 49099 100961
rect 48789 92147 48837 92175
rect 48865 92147 48899 92175
rect 48927 92147 48961 92175
rect 48989 92147 49023 92175
rect 49051 92147 49099 92175
rect 48789 92113 49099 92147
rect 48789 92085 48837 92113
rect 48865 92085 48899 92113
rect 48927 92085 48961 92113
rect 48989 92085 49023 92113
rect 49051 92085 49099 92113
rect 48789 92051 49099 92085
rect 48789 92023 48837 92051
rect 48865 92023 48899 92051
rect 48927 92023 48961 92051
rect 48989 92023 49023 92051
rect 49051 92023 49099 92051
rect 48789 91989 49099 92023
rect 48789 91961 48837 91989
rect 48865 91961 48899 91989
rect 48927 91961 48961 91989
rect 48989 91961 49023 91989
rect 49051 91961 49099 91989
rect 35289 86147 35337 86175
rect 35365 86147 35399 86175
rect 35427 86147 35461 86175
rect 35489 86147 35523 86175
rect 35551 86147 35599 86175
rect 35289 86113 35599 86147
rect 35289 86085 35337 86113
rect 35365 86085 35399 86113
rect 35427 86085 35461 86113
rect 35489 86085 35523 86113
rect 35551 86085 35599 86113
rect 35289 86051 35599 86085
rect 35289 86023 35337 86051
rect 35365 86023 35399 86051
rect 35427 86023 35461 86051
rect 35489 86023 35523 86051
rect 35551 86023 35599 86051
rect 35289 85989 35599 86023
rect 35289 85961 35337 85989
rect 35365 85961 35399 85989
rect 35427 85961 35461 85989
rect 35489 85961 35523 85989
rect 35551 85961 35599 85989
rect 35289 77175 35599 85961
rect 46624 86175 46784 86192
rect 46624 86147 46659 86175
rect 46687 86147 46721 86175
rect 46749 86147 46784 86175
rect 46624 86113 46784 86147
rect 46624 86085 46659 86113
rect 46687 86085 46721 86113
rect 46749 86085 46784 86113
rect 46624 86051 46784 86085
rect 46624 86023 46659 86051
rect 46687 86023 46721 86051
rect 46749 86023 46784 86051
rect 46624 85989 46784 86023
rect 46624 85961 46659 85989
rect 46687 85961 46721 85989
rect 46749 85961 46784 85989
rect 46624 85944 46784 85961
rect 38944 83175 39104 83192
rect 38944 83147 38979 83175
rect 39007 83147 39041 83175
rect 39069 83147 39104 83175
rect 38944 83113 39104 83147
rect 38944 83085 38979 83113
rect 39007 83085 39041 83113
rect 39069 83085 39104 83113
rect 38944 83051 39104 83085
rect 38944 83023 38979 83051
rect 39007 83023 39041 83051
rect 39069 83023 39104 83051
rect 38944 82989 39104 83023
rect 38944 82961 38979 82989
rect 39007 82961 39041 82989
rect 39069 82961 39104 82989
rect 38944 82944 39104 82961
rect 48789 83175 49099 91961
rect 48789 83147 48837 83175
rect 48865 83147 48899 83175
rect 48927 83147 48961 83175
rect 48989 83147 49023 83175
rect 49051 83147 49099 83175
rect 48789 83113 49099 83147
rect 48789 83085 48837 83113
rect 48865 83085 48899 83113
rect 48927 83085 48961 83113
rect 48989 83085 49023 83113
rect 49051 83085 49099 83113
rect 48789 83051 49099 83085
rect 48789 83023 48837 83051
rect 48865 83023 48899 83051
rect 48927 83023 48961 83051
rect 48989 83023 49023 83051
rect 49051 83023 49099 83051
rect 48789 82989 49099 83023
rect 48789 82961 48837 82989
rect 48865 82961 48899 82989
rect 48927 82961 48961 82989
rect 48989 82961 49023 82989
rect 49051 82961 49099 82989
rect 35289 77147 35337 77175
rect 35365 77147 35399 77175
rect 35427 77147 35461 77175
rect 35489 77147 35523 77175
rect 35551 77147 35599 77175
rect 35289 77113 35599 77147
rect 35289 77085 35337 77113
rect 35365 77085 35399 77113
rect 35427 77085 35461 77113
rect 35489 77085 35523 77113
rect 35551 77085 35599 77113
rect 35289 77051 35599 77085
rect 35289 77023 35337 77051
rect 35365 77023 35399 77051
rect 35427 77023 35461 77051
rect 35489 77023 35523 77051
rect 35551 77023 35599 77051
rect 35289 76989 35599 77023
rect 35289 76961 35337 76989
rect 35365 76961 35399 76989
rect 35427 76961 35461 76989
rect 35489 76961 35523 76989
rect 35551 76961 35599 76989
rect 35289 68175 35599 76961
rect 46624 77175 46784 77192
rect 46624 77147 46659 77175
rect 46687 77147 46721 77175
rect 46749 77147 46784 77175
rect 46624 77113 46784 77147
rect 46624 77085 46659 77113
rect 46687 77085 46721 77113
rect 46749 77085 46784 77113
rect 46624 77051 46784 77085
rect 46624 77023 46659 77051
rect 46687 77023 46721 77051
rect 46749 77023 46784 77051
rect 46624 76989 46784 77023
rect 46624 76961 46659 76989
rect 46687 76961 46721 76989
rect 46749 76961 46784 76989
rect 46624 76944 46784 76961
rect 38944 74175 39104 74192
rect 38944 74147 38979 74175
rect 39007 74147 39041 74175
rect 39069 74147 39104 74175
rect 38944 74113 39104 74147
rect 38944 74085 38979 74113
rect 39007 74085 39041 74113
rect 39069 74085 39104 74113
rect 38944 74051 39104 74085
rect 38944 74023 38979 74051
rect 39007 74023 39041 74051
rect 39069 74023 39104 74051
rect 38944 73989 39104 74023
rect 38944 73961 38979 73989
rect 39007 73961 39041 73989
rect 39069 73961 39104 73989
rect 38944 73944 39104 73961
rect 48789 74175 49099 82961
rect 48789 74147 48837 74175
rect 48865 74147 48899 74175
rect 48927 74147 48961 74175
rect 48989 74147 49023 74175
rect 49051 74147 49099 74175
rect 48789 74113 49099 74147
rect 48789 74085 48837 74113
rect 48865 74085 48899 74113
rect 48927 74085 48961 74113
rect 48989 74085 49023 74113
rect 49051 74085 49099 74113
rect 48789 74051 49099 74085
rect 48789 74023 48837 74051
rect 48865 74023 48899 74051
rect 48927 74023 48961 74051
rect 48989 74023 49023 74051
rect 49051 74023 49099 74051
rect 48789 73989 49099 74023
rect 48789 73961 48837 73989
rect 48865 73961 48899 73989
rect 48927 73961 48961 73989
rect 48989 73961 49023 73989
rect 49051 73961 49099 73989
rect 35289 68147 35337 68175
rect 35365 68147 35399 68175
rect 35427 68147 35461 68175
rect 35489 68147 35523 68175
rect 35551 68147 35599 68175
rect 35289 68113 35599 68147
rect 35289 68085 35337 68113
rect 35365 68085 35399 68113
rect 35427 68085 35461 68113
rect 35489 68085 35523 68113
rect 35551 68085 35599 68113
rect 35289 68051 35599 68085
rect 35289 68023 35337 68051
rect 35365 68023 35399 68051
rect 35427 68023 35461 68051
rect 35489 68023 35523 68051
rect 35551 68023 35599 68051
rect 35289 67989 35599 68023
rect 35289 67961 35337 67989
rect 35365 67961 35399 67989
rect 35427 67961 35461 67989
rect 35489 67961 35523 67989
rect 35551 67961 35599 67989
rect 35289 59175 35599 67961
rect 46624 68175 46784 68192
rect 46624 68147 46659 68175
rect 46687 68147 46721 68175
rect 46749 68147 46784 68175
rect 46624 68113 46784 68147
rect 46624 68085 46659 68113
rect 46687 68085 46721 68113
rect 46749 68085 46784 68113
rect 46624 68051 46784 68085
rect 46624 68023 46659 68051
rect 46687 68023 46721 68051
rect 46749 68023 46784 68051
rect 46624 67989 46784 68023
rect 46624 67961 46659 67989
rect 46687 67961 46721 67989
rect 46749 67961 46784 67989
rect 46624 67944 46784 67961
rect 38944 65175 39104 65192
rect 38944 65147 38979 65175
rect 39007 65147 39041 65175
rect 39069 65147 39104 65175
rect 38944 65113 39104 65147
rect 38944 65085 38979 65113
rect 39007 65085 39041 65113
rect 39069 65085 39104 65113
rect 38944 65051 39104 65085
rect 38944 65023 38979 65051
rect 39007 65023 39041 65051
rect 39069 65023 39104 65051
rect 38944 64989 39104 65023
rect 38944 64961 38979 64989
rect 39007 64961 39041 64989
rect 39069 64961 39104 64989
rect 38944 64944 39104 64961
rect 48789 65175 49099 73961
rect 48789 65147 48837 65175
rect 48865 65147 48899 65175
rect 48927 65147 48961 65175
rect 48989 65147 49023 65175
rect 49051 65147 49099 65175
rect 48789 65113 49099 65147
rect 48789 65085 48837 65113
rect 48865 65085 48899 65113
rect 48927 65085 48961 65113
rect 48989 65085 49023 65113
rect 49051 65085 49099 65113
rect 48789 65051 49099 65085
rect 48789 65023 48837 65051
rect 48865 65023 48899 65051
rect 48927 65023 48961 65051
rect 48989 65023 49023 65051
rect 49051 65023 49099 65051
rect 48789 64989 49099 65023
rect 48789 64961 48837 64989
rect 48865 64961 48899 64989
rect 48927 64961 48961 64989
rect 48989 64961 49023 64989
rect 49051 64961 49099 64989
rect 35289 59147 35337 59175
rect 35365 59147 35399 59175
rect 35427 59147 35461 59175
rect 35489 59147 35523 59175
rect 35551 59147 35599 59175
rect 35289 59113 35599 59147
rect 35289 59085 35337 59113
rect 35365 59085 35399 59113
rect 35427 59085 35461 59113
rect 35489 59085 35523 59113
rect 35551 59085 35599 59113
rect 35289 59051 35599 59085
rect 35289 59023 35337 59051
rect 35365 59023 35399 59051
rect 35427 59023 35461 59051
rect 35489 59023 35523 59051
rect 35551 59023 35599 59051
rect 35289 58989 35599 59023
rect 35289 58961 35337 58989
rect 35365 58961 35399 58989
rect 35427 58961 35461 58989
rect 35489 58961 35523 58989
rect 35551 58961 35599 58989
rect 35289 50175 35599 58961
rect 46624 59175 46784 59192
rect 46624 59147 46659 59175
rect 46687 59147 46721 59175
rect 46749 59147 46784 59175
rect 46624 59113 46784 59147
rect 46624 59085 46659 59113
rect 46687 59085 46721 59113
rect 46749 59085 46784 59113
rect 46624 59051 46784 59085
rect 46624 59023 46659 59051
rect 46687 59023 46721 59051
rect 46749 59023 46784 59051
rect 46624 58989 46784 59023
rect 46624 58961 46659 58989
rect 46687 58961 46721 58989
rect 46749 58961 46784 58989
rect 46624 58944 46784 58961
rect 38944 56175 39104 56192
rect 38944 56147 38979 56175
rect 39007 56147 39041 56175
rect 39069 56147 39104 56175
rect 38944 56113 39104 56147
rect 38944 56085 38979 56113
rect 39007 56085 39041 56113
rect 39069 56085 39104 56113
rect 38944 56051 39104 56085
rect 38944 56023 38979 56051
rect 39007 56023 39041 56051
rect 39069 56023 39104 56051
rect 38944 55989 39104 56023
rect 38944 55961 38979 55989
rect 39007 55961 39041 55989
rect 39069 55961 39104 55989
rect 38944 55944 39104 55961
rect 48789 56175 49099 64961
rect 48789 56147 48837 56175
rect 48865 56147 48899 56175
rect 48927 56147 48961 56175
rect 48989 56147 49023 56175
rect 49051 56147 49099 56175
rect 48789 56113 49099 56147
rect 48789 56085 48837 56113
rect 48865 56085 48899 56113
rect 48927 56085 48961 56113
rect 48989 56085 49023 56113
rect 49051 56085 49099 56113
rect 48789 56051 49099 56085
rect 48789 56023 48837 56051
rect 48865 56023 48899 56051
rect 48927 56023 48961 56051
rect 48989 56023 49023 56051
rect 49051 56023 49099 56051
rect 48789 55989 49099 56023
rect 48789 55961 48837 55989
rect 48865 55961 48899 55989
rect 48927 55961 48961 55989
rect 48989 55961 49023 55989
rect 49051 55961 49099 55989
rect 35289 50147 35337 50175
rect 35365 50147 35399 50175
rect 35427 50147 35461 50175
rect 35489 50147 35523 50175
rect 35551 50147 35599 50175
rect 35289 50113 35599 50147
rect 35289 50085 35337 50113
rect 35365 50085 35399 50113
rect 35427 50085 35461 50113
rect 35489 50085 35523 50113
rect 35551 50085 35599 50113
rect 35289 50051 35599 50085
rect 35289 50023 35337 50051
rect 35365 50023 35399 50051
rect 35427 50023 35461 50051
rect 35489 50023 35523 50051
rect 35551 50023 35599 50051
rect 35289 49989 35599 50023
rect 35289 49961 35337 49989
rect 35365 49961 35399 49989
rect 35427 49961 35461 49989
rect 35489 49961 35523 49989
rect 35551 49961 35599 49989
rect 35289 41175 35599 49961
rect 46624 50175 46784 50192
rect 46624 50147 46659 50175
rect 46687 50147 46721 50175
rect 46749 50147 46784 50175
rect 46624 50113 46784 50147
rect 46624 50085 46659 50113
rect 46687 50085 46721 50113
rect 46749 50085 46784 50113
rect 46624 50051 46784 50085
rect 46624 50023 46659 50051
rect 46687 50023 46721 50051
rect 46749 50023 46784 50051
rect 46624 49989 46784 50023
rect 46624 49961 46659 49989
rect 46687 49961 46721 49989
rect 46749 49961 46784 49989
rect 46624 49944 46784 49961
rect 38944 47175 39104 47192
rect 38944 47147 38979 47175
rect 39007 47147 39041 47175
rect 39069 47147 39104 47175
rect 38944 47113 39104 47147
rect 38944 47085 38979 47113
rect 39007 47085 39041 47113
rect 39069 47085 39104 47113
rect 38944 47051 39104 47085
rect 38944 47023 38979 47051
rect 39007 47023 39041 47051
rect 39069 47023 39104 47051
rect 38944 46989 39104 47023
rect 38944 46961 38979 46989
rect 39007 46961 39041 46989
rect 39069 46961 39104 46989
rect 38944 46944 39104 46961
rect 48789 47175 49099 55961
rect 48789 47147 48837 47175
rect 48865 47147 48899 47175
rect 48927 47147 48961 47175
rect 48989 47147 49023 47175
rect 49051 47147 49099 47175
rect 48789 47113 49099 47147
rect 48789 47085 48837 47113
rect 48865 47085 48899 47113
rect 48927 47085 48961 47113
rect 48989 47085 49023 47113
rect 49051 47085 49099 47113
rect 48789 47051 49099 47085
rect 48789 47023 48837 47051
rect 48865 47023 48899 47051
rect 48927 47023 48961 47051
rect 48989 47023 49023 47051
rect 49051 47023 49099 47051
rect 48789 46989 49099 47023
rect 48789 46961 48837 46989
rect 48865 46961 48899 46989
rect 48927 46961 48961 46989
rect 48989 46961 49023 46989
rect 49051 46961 49099 46989
rect 35289 41147 35337 41175
rect 35365 41147 35399 41175
rect 35427 41147 35461 41175
rect 35489 41147 35523 41175
rect 35551 41147 35599 41175
rect 35289 41113 35599 41147
rect 35289 41085 35337 41113
rect 35365 41085 35399 41113
rect 35427 41085 35461 41113
rect 35489 41085 35523 41113
rect 35551 41085 35599 41113
rect 35289 41051 35599 41085
rect 35289 41023 35337 41051
rect 35365 41023 35399 41051
rect 35427 41023 35461 41051
rect 35489 41023 35523 41051
rect 35551 41023 35599 41051
rect 35289 40989 35599 41023
rect 35289 40961 35337 40989
rect 35365 40961 35399 40989
rect 35427 40961 35461 40989
rect 35489 40961 35523 40989
rect 35551 40961 35599 40989
rect 35289 32175 35599 40961
rect 46624 41175 46784 41192
rect 46624 41147 46659 41175
rect 46687 41147 46721 41175
rect 46749 41147 46784 41175
rect 46624 41113 46784 41147
rect 46624 41085 46659 41113
rect 46687 41085 46721 41113
rect 46749 41085 46784 41113
rect 46624 41051 46784 41085
rect 46624 41023 46659 41051
rect 46687 41023 46721 41051
rect 46749 41023 46784 41051
rect 46624 40989 46784 41023
rect 46624 40961 46659 40989
rect 46687 40961 46721 40989
rect 46749 40961 46784 40989
rect 46624 40944 46784 40961
rect 38944 38175 39104 38192
rect 38944 38147 38979 38175
rect 39007 38147 39041 38175
rect 39069 38147 39104 38175
rect 38944 38113 39104 38147
rect 38944 38085 38979 38113
rect 39007 38085 39041 38113
rect 39069 38085 39104 38113
rect 38944 38051 39104 38085
rect 38944 38023 38979 38051
rect 39007 38023 39041 38051
rect 39069 38023 39104 38051
rect 38944 37989 39104 38023
rect 38944 37961 38979 37989
rect 39007 37961 39041 37989
rect 39069 37961 39104 37989
rect 38944 37944 39104 37961
rect 48789 38175 49099 46961
rect 48789 38147 48837 38175
rect 48865 38147 48899 38175
rect 48927 38147 48961 38175
rect 48989 38147 49023 38175
rect 49051 38147 49099 38175
rect 48789 38113 49099 38147
rect 48789 38085 48837 38113
rect 48865 38085 48899 38113
rect 48927 38085 48961 38113
rect 48989 38085 49023 38113
rect 49051 38085 49099 38113
rect 48789 38051 49099 38085
rect 48789 38023 48837 38051
rect 48865 38023 48899 38051
rect 48927 38023 48961 38051
rect 48989 38023 49023 38051
rect 49051 38023 49099 38051
rect 48789 37989 49099 38023
rect 48789 37961 48837 37989
rect 48865 37961 48899 37989
rect 48927 37961 48961 37989
rect 48989 37961 49023 37989
rect 49051 37961 49099 37989
rect 35289 32147 35337 32175
rect 35365 32147 35399 32175
rect 35427 32147 35461 32175
rect 35489 32147 35523 32175
rect 35551 32147 35599 32175
rect 35289 32113 35599 32147
rect 35289 32085 35337 32113
rect 35365 32085 35399 32113
rect 35427 32085 35461 32113
rect 35489 32085 35523 32113
rect 35551 32085 35599 32113
rect 35289 32051 35599 32085
rect 35289 32023 35337 32051
rect 35365 32023 35399 32051
rect 35427 32023 35461 32051
rect 35489 32023 35523 32051
rect 35551 32023 35599 32051
rect 35289 31989 35599 32023
rect 35289 31961 35337 31989
rect 35365 31961 35399 31989
rect 35427 31961 35461 31989
rect 35489 31961 35523 31989
rect 35551 31961 35599 31989
rect 35289 23175 35599 31961
rect 46624 32175 46784 32192
rect 46624 32147 46659 32175
rect 46687 32147 46721 32175
rect 46749 32147 46784 32175
rect 46624 32113 46784 32147
rect 46624 32085 46659 32113
rect 46687 32085 46721 32113
rect 46749 32085 46784 32113
rect 46624 32051 46784 32085
rect 46624 32023 46659 32051
rect 46687 32023 46721 32051
rect 46749 32023 46784 32051
rect 46624 31989 46784 32023
rect 46624 31961 46659 31989
rect 46687 31961 46721 31989
rect 46749 31961 46784 31989
rect 46624 31944 46784 31961
rect 38944 29175 39104 29192
rect 38944 29147 38979 29175
rect 39007 29147 39041 29175
rect 39069 29147 39104 29175
rect 38944 29113 39104 29147
rect 38944 29085 38979 29113
rect 39007 29085 39041 29113
rect 39069 29085 39104 29113
rect 38944 29051 39104 29085
rect 38944 29023 38979 29051
rect 39007 29023 39041 29051
rect 39069 29023 39104 29051
rect 38944 28989 39104 29023
rect 38944 28961 38979 28989
rect 39007 28961 39041 28989
rect 39069 28961 39104 28989
rect 38944 28944 39104 28961
rect 48789 29175 49099 37961
rect 48789 29147 48837 29175
rect 48865 29147 48899 29175
rect 48927 29147 48961 29175
rect 48989 29147 49023 29175
rect 49051 29147 49099 29175
rect 48789 29113 49099 29147
rect 48789 29085 48837 29113
rect 48865 29085 48899 29113
rect 48927 29085 48961 29113
rect 48989 29085 49023 29113
rect 49051 29085 49099 29113
rect 48789 29051 49099 29085
rect 48789 29023 48837 29051
rect 48865 29023 48899 29051
rect 48927 29023 48961 29051
rect 48989 29023 49023 29051
rect 49051 29023 49099 29051
rect 48789 28989 49099 29023
rect 48789 28961 48837 28989
rect 48865 28961 48899 28989
rect 48927 28961 48961 28989
rect 48989 28961 49023 28989
rect 49051 28961 49099 28989
rect 35289 23147 35337 23175
rect 35365 23147 35399 23175
rect 35427 23147 35461 23175
rect 35489 23147 35523 23175
rect 35551 23147 35599 23175
rect 35289 23113 35599 23147
rect 35289 23085 35337 23113
rect 35365 23085 35399 23113
rect 35427 23085 35461 23113
rect 35489 23085 35523 23113
rect 35551 23085 35599 23113
rect 35289 23051 35599 23085
rect 35289 23023 35337 23051
rect 35365 23023 35399 23051
rect 35427 23023 35461 23051
rect 35489 23023 35523 23051
rect 35551 23023 35599 23051
rect 35289 22989 35599 23023
rect 35289 22961 35337 22989
rect 35365 22961 35399 22989
rect 35427 22961 35461 22989
rect 35489 22961 35523 22989
rect 35551 22961 35599 22989
rect 35289 14175 35599 22961
rect 46624 23175 46784 23192
rect 46624 23147 46659 23175
rect 46687 23147 46721 23175
rect 46749 23147 46784 23175
rect 46624 23113 46784 23147
rect 46624 23085 46659 23113
rect 46687 23085 46721 23113
rect 46749 23085 46784 23113
rect 46624 23051 46784 23085
rect 46624 23023 46659 23051
rect 46687 23023 46721 23051
rect 46749 23023 46784 23051
rect 46624 22989 46784 23023
rect 46624 22961 46659 22989
rect 46687 22961 46721 22989
rect 46749 22961 46784 22989
rect 46624 22944 46784 22961
rect 38944 20175 39104 20192
rect 38944 20147 38979 20175
rect 39007 20147 39041 20175
rect 39069 20147 39104 20175
rect 38944 20113 39104 20147
rect 38944 20085 38979 20113
rect 39007 20085 39041 20113
rect 39069 20085 39104 20113
rect 38944 20051 39104 20085
rect 38944 20023 38979 20051
rect 39007 20023 39041 20051
rect 39069 20023 39104 20051
rect 38944 19989 39104 20023
rect 38944 19961 38979 19989
rect 39007 19961 39041 19989
rect 39069 19961 39104 19989
rect 38944 19944 39104 19961
rect 48789 20175 49099 28961
rect 48789 20147 48837 20175
rect 48865 20147 48899 20175
rect 48927 20147 48961 20175
rect 48989 20147 49023 20175
rect 49051 20147 49099 20175
rect 48789 20113 49099 20147
rect 48789 20085 48837 20113
rect 48865 20085 48899 20113
rect 48927 20085 48961 20113
rect 48989 20085 49023 20113
rect 49051 20085 49099 20113
rect 48789 20051 49099 20085
rect 48789 20023 48837 20051
rect 48865 20023 48899 20051
rect 48927 20023 48961 20051
rect 48989 20023 49023 20051
rect 49051 20023 49099 20051
rect 48789 19989 49099 20023
rect 48789 19961 48837 19989
rect 48865 19961 48899 19989
rect 48927 19961 48961 19989
rect 48989 19961 49023 19989
rect 49051 19961 49099 19989
rect 35289 14147 35337 14175
rect 35365 14147 35399 14175
rect 35427 14147 35461 14175
rect 35489 14147 35523 14175
rect 35551 14147 35599 14175
rect 35289 14113 35599 14147
rect 35289 14085 35337 14113
rect 35365 14085 35399 14113
rect 35427 14085 35461 14113
rect 35489 14085 35523 14113
rect 35551 14085 35599 14113
rect 35289 14051 35599 14085
rect 35289 14023 35337 14051
rect 35365 14023 35399 14051
rect 35427 14023 35461 14051
rect 35489 14023 35523 14051
rect 35551 14023 35599 14051
rect 35289 13989 35599 14023
rect 35289 13961 35337 13989
rect 35365 13961 35399 13989
rect 35427 13961 35461 13989
rect 35489 13961 35523 13989
rect 35551 13961 35599 13989
rect 35289 5175 35599 13961
rect 46624 14175 46784 14192
rect 46624 14147 46659 14175
rect 46687 14147 46721 14175
rect 46749 14147 46784 14175
rect 46624 14113 46784 14147
rect 46624 14085 46659 14113
rect 46687 14085 46721 14113
rect 46749 14085 46784 14113
rect 46624 14051 46784 14085
rect 46624 14023 46659 14051
rect 46687 14023 46721 14051
rect 46749 14023 46784 14051
rect 46624 13989 46784 14023
rect 46624 13961 46659 13989
rect 46687 13961 46721 13989
rect 46749 13961 46784 13989
rect 46624 13944 46784 13961
rect 38944 11175 39104 11192
rect 38944 11147 38979 11175
rect 39007 11147 39041 11175
rect 39069 11147 39104 11175
rect 38944 11113 39104 11147
rect 38944 11085 38979 11113
rect 39007 11085 39041 11113
rect 39069 11085 39104 11113
rect 38944 11051 39104 11085
rect 38944 11023 38979 11051
rect 39007 11023 39041 11051
rect 39069 11023 39104 11051
rect 38944 10989 39104 11023
rect 38944 10961 38979 10989
rect 39007 10961 39041 10989
rect 39069 10961 39104 10989
rect 38944 10944 39104 10961
rect 48789 11175 49099 19961
rect 48789 11147 48837 11175
rect 48865 11147 48899 11175
rect 48927 11147 48961 11175
rect 48989 11147 49023 11175
rect 49051 11147 49099 11175
rect 48789 11113 49099 11147
rect 48789 11085 48837 11113
rect 48865 11085 48899 11113
rect 48927 11085 48961 11113
rect 48989 11085 49023 11113
rect 49051 11085 49099 11113
rect 48789 11051 49099 11085
rect 48789 11023 48837 11051
rect 48865 11023 48899 11051
rect 48927 11023 48961 11051
rect 48989 11023 49023 11051
rect 49051 11023 49099 11051
rect 48789 10989 49099 11023
rect 48789 10961 48837 10989
rect 48865 10961 48899 10989
rect 48927 10961 48961 10989
rect 48989 10961 49023 10989
rect 49051 10961 49099 10989
rect 35289 5147 35337 5175
rect 35365 5147 35399 5175
rect 35427 5147 35461 5175
rect 35489 5147 35523 5175
rect 35551 5147 35599 5175
rect 35289 5113 35599 5147
rect 35289 5085 35337 5113
rect 35365 5085 35399 5113
rect 35427 5085 35461 5113
rect 35489 5085 35523 5113
rect 35551 5085 35599 5113
rect 35289 5051 35599 5085
rect 35289 5023 35337 5051
rect 35365 5023 35399 5051
rect 35427 5023 35461 5051
rect 35489 5023 35523 5051
rect 35551 5023 35599 5051
rect 35289 4989 35599 5023
rect 35289 4961 35337 4989
rect 35365 4961 35399 4989
rect 35427 4961 35461 4989
rect 35489 4961 35523 4989
rect 35551 4961 35599 4989
rect 35289 -560 35599 4961
rect 46624 5175 46784 5192
rect 46624 5147 46659 5175
rect 46687 5147 46721 5175
rect 46749 5147 46784 5175
rect 46624 5113 46784 5147
rect 46624 5085 46659 5113
rect 46687 5085 46721 5113
rect 46749 5085 46784 5113
rect 46624 5051 46784 5085
rect 46624 5023 46659 5051
rect 46687 5023 46721 5051
rect 46749 5023 46784 5051
rect 46624 4989 46784 5023
rect 46624 4961 46659 4989
rect 46687 4961 46721 4989
rect 46749 4961 46784 4989
rect 46624 4944 46784 4961
rect 35289 -588 35337 -560
rect 35365 -588 35399 -560
rect 35427 -588 35461 -560
rect 35489 -588 35523 -560
rect 35551 -588 35599 -560
rect 35289 -622 35599 -588
rect 35289 -650 35337 -622
rect 35365 -650 35399 -622
rect 35427 -650 35461 -622
rect 35489 -650 35523 -622
rect 35551 -650 35599 -622
rect 35289 -684 35599 -650
rect 35289 -712 35337 -684
rect 35365 -712 35399 -684
rect 35427 -712 35461 -684
rect 35489 -712 35523 -684
rect 35551 -712 35599 -684
rect 35289 -746 35599 -712
rect 35289 -774 35337 -746
rect 35365 -774 35399 -746
rect 35427 -774 35461 -746
rect 35489 -774 35523 -746
rect 35551 -774 35599 -746
rect 35289 -822 35599 -774
rect 48789 2175 49099 10961
rect 48789 2147 48837 2175
rect 48865 2147 48899 2175
rect 48927 2147 48961 2175
rect 48989 2147 49023 2175
rect 49051 2147 49099 2175
rect 48789 2113 49099 2147
rect 48789 2085 48837 2113
rect 48865 2085 48899 2113
rect 48927 2085 48961 2113
rect 48989 2085 49023 2113
rect 49051 2085 49099 2113
rect 48789 2051 49099 2085
rect 48789 2023 48837 2051
rect 48865 2023 48899 2051
rect 48927 2023 48961 2051
rect 48989 2023 49023 2051
rect 49051 2023 49099 2051
rect 48789 1989 49099 2023
rect 48789 1961 48837 1989
rect 48865 1961 48899 1989
rect 48927 1961 48961 1989
rect 48989 1961 49023 1989
rect 49051 1961 49099 1989
rect 48789 -80 49099 1961
rect 48789 -108 48837 -80
rect 48865 -108 48899 -80
rect 48927 -108 48961 -80
rect 48989 -108 49023 -80
rect 49051 -108 49099 -80
rect 48789 -142 49099 -108
rect 48789 -170 48837 -142
rect 48865 -170 48899 -142
rect 48927 -170 48961 -142
rect 48989 -170 49023 -142
rect 49051 -170 49099 -142
rect 48789 -204 49099 -170
rect 48789 -232 48837 -204
rect 48865 -232 48899 -204
rect 48927 -232 48961 -204
rect 48989 -232 49023 -204
rect 49051 -232 49099 -204
rect 48789 -266 49099 -232
rect 48789 -294 48837 -266
rect 48865 -294 48899 -266
rect 48927 -294 48961 -266
rect 48989 -294 49023 -266
rect 49051 -294 49099 -266
rect 48789 -822 49099 -294
rect 50649 299086 50959 299134
rect 50649 299058 50697 299086
rect 50725 299058 50759 299086
rect 50787 299058 50821 299086
rect 50849 299058 50883 299086
rect 50911 299058 50959 299086
rect 50649 299024 50959 299058
rect 50649 298996 50697 299024
rect 50725 298996 50759 299024
rect 50787 298996 50821 299024
rect 50849 298996 50883 299024
rect 50911 298996 50959 299024
rect 50649 298962 50959 298996
rect 50649 298934 50697 298962
rect 50725 298934 50759 298962
rect 50787 298934 50821 298962
rect 50849 298934 50883 298962
rect 50911 298934 50959 298962
rect 50649 298900 50959 298934
rect 50649 298872 50697 298900
rect 50725 298872 50759 298900
rect 50787 298872 50821 298900
rect 50849 298872 50883 298900
rect 50911 298872 50959 298900
rect 50649 293175 50959 298872
rect 50649 293147 50697 293175
rect 50725 293147 50759 293175
rect 50787 293147 50821 293175
rect 50849 293147 50883 293175
rect 50911 293147 50959 293175
rect 50649 293113 50959 293147
rect 50649 293085 50697 293113
rect 50725 293085 50759 293113
rect 50787 293085 50821 293113
rect 50849 293085 50883 293113
rect 50911 293085 50959 293113
rect 50649 293051 50959 293085
rect 50649 293023 50697 293051
rect 50725 293023 50759 293051
rect 50787 293023 50821 293051
rect 50849 293023 50883 293051
rect 50911 293023 50959 293051
rect 50649 292989 50959 293023
rect 50649 292961 50697 292989
rect 50725 292961 50759 292989
rect 50787 292961 50821 292989
rect 50849 292961 50883 292989
rect 50911 292961 50959 292989
rect 50649 284175 50959 292961
rect 50649 284147 50697 284175
rect 50725 284147 50759 284175
rect 50787 284147 50821 284175
rect 50849 284147 50883 284175
rect 50911 284147 50959 284175
rect 50649 284113 50959 284147
rect 50649 284085 50697 284113
rect 50725 284085 50759 284113
rect 50787 284085 50821 284113
rect 50849 284085 50883 284113
rect 50911 284085 50959 284113
rect 50649 284051 50959 284085
rect 50649 284023 50697 284051
rect 50725 284023 50759 284051
rect 50787 284023 50821 284051
rect 50849 284023 50883 284051
rect 50911 284023 50959 284051
rect 50649 283989 50959 284023
rect 50649 283961 50697 283989
rect 50725 283961 50759 283989
rect 50787 283961 50821 283989
rect 50849 283961 50883 283989
rect 50911 283961 50959 283989
rect 50649 275175 50959 283961
rect 50649 275147 50697 275175
rect 50725 275147 50759 275175
rect 50787 275147 50821 275175
rect 50849 275147 50883 275175
rect 50911 275147 50959 275175
rect 50649 275113 50959 275147
rect 50649 275085 50697 275113
rect 50725 275085 50759 275113
rect 50787 275085 50821 275113
rect 50849 275085 50883 275113
rect 50911 275085 50959 275113
rect 50649 275051 50959 275085
rect 50649 275023 50697 275051
rect 50725 275023 50759 275051
rect 50787 275023 50821 275051
rect 50849 275023 50883 275051
rect 50911 275023 50959 275051
rect 50649 274989 50959 275023
rect 50649 274961 50697 274989
rect 50725 274961 50759 274989
rect 50787 274961 50821 274989
rect 50849 274961 50883 274989
rect 50911 274961 50959 274989
rect 50649 266175 50959 274961
rect 50649 266147 50697 266175
rect 50725 266147 50759 266175
rect 50787 266147 50821 266175
rect 50849 266147 50883 266175
rect 50911 266147 50959 266175
rect 50649 266113 50959 266147
rect 50649 266085 50697 266113
rect 50725 266085 50759 266113
rect 50787 266085 50821 266113
rect 50849 266085 50883 266113
rect 50911 266085 50959 266113
rect 50649 266051 50959 266085
rect 50649 266023 50697 266051
rect 50725 266023 50759 266051
rect 50787 266023 50821 266051
rect 50849 266023 50883 266051
rect 50911 266023 50959 266051
rect 50649 265989 50959 266023
rect 50649 265961 50697 265989
rect 50725 265961 50759 265989
rect 50787 265961 50821 265989
rect 50849 265961 50883 265989
rect 50911 265961 50959 265989
rect 50649 257175 50959 265961
rect 50649 257147 50697 257175
rect 50725 257147 50759 257175
rect 50787 257147 50821 257175
rect 50849 257147 50883 257175
rect 50911 257147 50959 257175
rect 50649 257113 50959 257147
rect 50649 257085 50697 257113
rect 50725 257085 50759 257113
rect 50787 257085 50821 257113
rect 50849 257085 50883 257113
rect 50911 257085 50959 257113
rect 50649 257051 50959 257085
rect 50649 257023 50697 257051
rect 50725 257023 50759 257051
rect 50787 257023 50821 257051
rect 50849 257023 50883 257051
rect 50911 257023 50959 257051
rect 50649 256989 50959 257023
rect 50649 256961 50697 256989
rect 50725 256961 50759 256989
rect 50787 256961 50821 256989
rect 50849 256961 50883 256989
rect 50911 256961 50959 256989
rect 50649 248175 50959 256961
rect 50649 248147 50697 248175
rect 50725 248147 50759 248175
rect 50787 248147 50821 248175
rect 50849 248147 50883 248175
rect 50911 248147 50959 248175
rect 50649 248113 50959 248147
rect 50649 248085 50697 248113
rect 50725 248085 50759 248113
rect 50787 248085 50821 248113
rect 50849 248085 50883 248113
rect 50911 248085 50959 248113
rect 50649 248051 50959 248085
rect 50649 248023 50697 248051
rect 50725 248023 50759 248051
rect 50787 248023 50821 248051
rect 50849 248023 50883 248051
rect 50911 248023 50959 248051
rect 50649 247989 50959 248023
rect 50649 247961 50697 247989
rect 50725 247961 50759 247989
rect 50787 247961 50821 247989
rect 50849 247961 50883 247989
rect 50911 247961 50959 247989
rect 50649 239175 50959 247961
rect 50649 239147 50697 239175
rect 50725 239147 50759 239175
rect 50787 239147 50821 239175
rect 50849 239147 50883 239175
rect 50911 239147 50959 239175
rect 50649 239113 50959 239147
rect 50649 239085 50697 239113
rect 50725 239085 50759 239113
rect 50787 239085 50821 239113
rect 50849 239085 50883 239113
rect 50911 239085 50959 239113
rect 50649 239051 50959 239085
rect 50649 239023 50697 239051
rect 50725 239023 50759 239051
rect 50787 239023 50821 239051
rect 50849 239023 50883 239051
rect 50911 239023 50959 239051
rect 50649 238989 50959 239023
rect 50649 238961 50697 238989
rect 50725 238961 50759 238989
rect 50787 238961 50821 238989
rect 50849 238961 50883 238989
rect 50911 238961 50959 238989
rect 50649 230175 50959 238961
rect 50649 230147 50697 230175
rect 50725 230147 50759 230175
rect 50787 230147 50821 230175
rect 50849 230147 50883 230175
rect 50911 230147 50959 230175
rect 50649 230113 50959 230147
rect 50649 230085 50697 230113
rect 50725 230085 50759 230113
rect 50787 230085 50821 230113
rect 50849 230085 50883 230113
rect 50911 230085 50959 230113
rect 50649 230051 50959 230085
rect 50649 230023 50697 230051
rect 50725 230023 50759 230051
rect 50787 230023 50821 230051
rect 50849 230023 50883 230051
rect 50911 230023 50959 230051
rect 50649 229989 50959 230023
rect 50649 229961 50697 229989
rect 50725 229961 50759 229989
rect 50787 229961 50821 229989
rect 50849 229961 50883 229989
rect 50911 229961 50959 229989
rect 50649 221175 50959 229961
rect 50649 221147 50697 221175
rect 50725 221147 50759 221175
rect 50787 221147 50821 221175
rect 50849 221147 50883 221175
rect 50911 221147 50959 221175
rect 50649 221113 50959 221147
rect 50649 221085 50697 221113
rect 50725 221085 50759 221113
rect 50787 221085 50821 221113
rect 50849 221085 50883 221113
rect 50911 221085 50959 221113
rect 50649 221051 50959 221085
rect 50649 221023 50697 221051
rect 50725 221023 50759 221051
rect 50787 221023 50821 221051
rect 50849 221023 50883 221051
rect 50911 221023 50959 221051
rect 50649 220989 50959 221023
rect 50649 220961 50697 220989
rect 50725 220961 50759 220989
rect 50787 220961 50821 220989
rect 50849 220961 50883 220989
rect 50911 220961 50959 220989
rect 50649 212175 50959 220961
rect 50649 212147 50697 212175
rect 50725 212147 50759 212175
rect 50787 212147 50821 212175
rect 50849 212147 50883 212175
rect 50911 212147 50959 212175
rect 50649 212113 50959 212147
rect 50649 212085 50697 212113
rect 50725 212085 50759 212113
rect 50787 212085 50821 212113
rect 50849 212085 50883 212113
rect 50911 212085 50959 212113
rect 50649 212051 50959 212085
rect 50649 212023 50697 212051
rect 50725 212023 50759 212051
rect 50787 212023 50821 212051
rect 50849 212023 50883 212051
rect 50911 212023 50959 212051
rect 50649 211989 50959 212023
rect 50649 211961 50697 211989
rect 50725 211961 50759 211989
rect 50787 211961 50821 211989
rect 50849 211961 50883 211989
rect 50911 211961 50959 211989
rect 50649 203175 50959 211961
rect 50649 203147 50697 203175
rect 50725 203147 50759 203175
rect 50787 203147 50821 203175
rect 50849 203147 50883 203175
rect 50911 203147 50959 203175
rect 50649 203113 50959 203147
rect 50649 203085 50697 203113
rect 50725 203085 50759 203113
rect 50787 203085 50821 203113
rect 50849 203085 50883 203113
rect 50911 203085 50959 203113
rect 50649 203051 50959 203085
rect 50649 203023 50697 203051
rect 50725 203023 50759 203051
rect 50787 203023 50821 203051
rect 50849 203023 50883 203051
rect 50911 203023 50959 203051
rect 50649 202989 50959 203023
rect 50649 202961 50697 202989
rect 50725 202961 50759 202989
rect 50787 202961 50821 202989
rect 50849 202961 50883 202989
rect 50911 202961 50959 202989
rect 50649 194175 50959 202961
rect 50649 194147 50697 194175
rect 50725 194147 50759 194175
rect 50787 194147 50821 194175
rect 50849 194147 50883 194175
rect 50911 194147 50959 194175
rect 50649 194113 50959 194147
rect 50649 194085 50697 194113
rect 50725 194085 50759 194113
rect 50787 194085 50821 194113
rect 50849 194085 50883 194113
rect 50911 194085 50959 194113
rect 50649 194051 50959 194085
rect 50649 194023 50697 194051
rect 50725 194023 50759 194051
rect 50787 194023 50821 194051
rect 50849 194023 50883 194051
rect 50911 194023 50959 194051
rect 50649 193989 50959 194023
rect 50649 193961 50697 193989
rect 50725 193961 50759 193989
rect 50787 193961 50821 193989
rect 50849 193961 50883 193989
rect 50911 193961 50959 193989
rect 50649 185175 50959 193961
rect 50649 185147 50697 185175
rect 50725 185147 50759 185175
rect 50787 185147 50821 185175
rect 50849 185147 50883 185175
rect 50911 185147 50959 185175
rect 50649 185113 50959 185147
rect 50649 185085 50697 185113
rect 50725 185085 50759 185113
rect 50787 185085 50821 185113
rect 50849 185085 50883 185113
rect 50911 185085 50959 185113
rect 50649 185051 50959 185085
rect 50649 185023 50697 185051
rect 50725 185023 50759 185051
rect 50787 185023 50821 185051
rect 50849 185023 50883 185051
rect 50911 185023 50959 185051
rect 50649 184989 50959 185023
rect 50649 184961 50697 184989
rect 50725 184961 50759 184989
rect 50787 184961 50821 184989
rect 50849 184961 50883 184989
rect 50911 184961 50959 184989
rect 50649 176175 50959 184961
rect 50649 176147 50697 176175
rect 50725 176147 50759 176175
rect 50787 176147 50821 176175
rect 50849 176147 50883 176175
rect 50911 176147 50959 176175
rect 50649 176113 50959 176147
rect 50649 176085 50697 176113
rect 50725 176085 50759 176113
rect 50787 176085 50821 176113
rect 50849 176085 50883 176113
rect 50911 176085 50959 176113
rect 50649 176051 50959 176085
rect 50649 176023 50697 176051
rect 50725 176023 50759 176051
rect 50787 176023 50821 176051
rect 50849 176023 50883 176051
rect 50911 176023 50959 176051
rect 50649 175989 50959 176023
rect 50649 175961 50697 175989
rect 50725 175961 50759 175989
rect 50787 175961 50821 175989
rect 50849 175961 50883 175989
rect 50911 175961 50959 175989
rect 50649 167175 50959 175961
rect 64149 298606 64459 299134
rect 64149 298578 64197 298606
rect 64225 298578 64259 298606
rect 64287 298578 64321 298606
rect 64349 298578 64383 298606
rect 64411 298578 64459 298606
rect 64149 298544 64459 298578
rect 64149 298516 64197 298544
rect 64225 298516 64259 298544
rect 64287 298516 64321 298544
rect 64349 298516 64383 298544
rect 64411 298516 64459 298544
rect 64149 298482 64459 298516
rect 64149 298454 64197 298482
rect 64225 298454 64259 298482
rect 64287 298454 64321 298482
rect 64349 298454 64383 298482
rect 64411 298454 64459 298482
rect 64149 298420 64459 298454
rect 64149 298392 64197 298420
rect 64225 298392 64259 298420
rect 64287 298392 64321 298420
rect 64349 298392 64383 298420
rect 64411 298392 64459 298420
rect 64149 290175 64459 298392
rect 64149 290147 64197 290175
rect 64225 290147 64259 290175
rect 64287 290147 64321 290175
rect 64349 290147 64383 290175
rect 64411 290147 64459 290175
rect 64149 290113 64459 290147
rect 64149 290085 64197 290113
rect 64225 290085 64259 290113
rect 64287 290085 64321 290113
rect 64349 290085 64383 290113
rect 64411 290085 64459 290113
rect 64149 290051 64459 290085
rect 64149 290023 64197 290051
rect 64225 290023 64259 290051
rect 64287 290023 64321 290051
rect 64349 290023 64383 290051
rect 64411 290023 64459 290051
rect 64149 289989 64459 290023
rect 64149 289961 64197 289989
rect 64225 289961 64259 289989
rect 64287 289961 64321 289989
rect 64349 289961 64383 289989
rect 64411 289961 64459 289989
rect 64149 281175 64459 289961
rect 64149 281147 64197 281175
rect 64225 281147 64259 281175
rect 64287 281147 64321 281175
rect 64349 281147 64383 281175
rect 64411 281147 64459 281175
rect 64149 281113 64459 281147
rect 64149 281085 64197 281113
rect 64225 281085 64259 281113
rect 64287 281085 64321 281113
rect 64349 281085 64383 281113
rect 64411 281085 64459 281113
rect 64149 281051 64459 281085
rect 64149 281023 64197 281051
rect 64225 281023 64259 281051
rect 64287 281023 64321 281051
rect 64349 281023 64383 281051
rect 64411 281023 64459 281051
rect 64149 280989 64459 281023
rect 64149 280961 64197 280989
rect 64225 280961 64259 280989
rect 64287 280961 64321 280989
rect 64349 280961 64383 280989
rect 64411 280961 64459 280989
rect 64149 272175 64459 280961
rect 64149 272147 64197 272175
rect 64225 272147 64259 272175
rect 64287 272147 64321 272175
rect 64349 272147 64383 272175
rect 64411 272147 64459 272175
rect 64149 272113 64459 272147
rect 64149 272085 64197 272113
rect 64225 272085 64259 272113
rect 64287 272085 64321 272113
rect 64349 272085 64383 272113
rect 64411 272085 64459 272113
rect 64149 272051 64459 272085
rect 64149 272023 64197 272051
rect 64225 272023 64259 272051
rect 64287 272023 64321 272051
rect 64349 272023 64383 272051
rect 64411 272023 64459 272051
rect 64149 271989 64459 272023
rect 64149 271961 64197 271989
rect 64225 271961 64259 271989
rect 64287 271961 64321 271989
rect 64349 271961 64383 271989
rect 64411 271961 64459 271989
rect 64149 263175 64459 271961
rect 64149 263147 64197 263175
rect 64225 263147 64259 263175
rect 64287 263147 64321 263175
rect 64349 263147 64383 263175
rect 64411 263147 64459 263175
rect 64149 263113 64459 263147
rect 64149 263085 64197 263113
rect 64225 263085 64259 263113
rect 64287 263085 64321 263113
rect 64349 263085 64383 263113
rect 64411 263085 64459 263113
rect 64149 263051 64459 263085
rect 64149 263023 64197 263051
rect 64225 263023 64259 263051
rect 64287 263023 64321 263051
rect 64349 263023 64383 263051
rect 64411 263023 64459 263051
rect 64149 262989 64459 263023
rect 64149 262961 64197 262989
rect 64225 262961 64259 262989
rect 64287 262961 64321 262989
rect 64349 262961 64383 262989
rect 64411 262961 64459 262989
rect 64149 254175 64459 262961
rect 64149 254147 64197 254175
rect 64225 254147 64259 254175
rect 64287 254147 64321 254175
rect 64349 254147 64383 254175
rect 64411 254147 64459 254175
rect 64149 254113 64459 254147
rect 64149 254085 64197 254113
rect 64225 254085 64259 254113
rect 64287 254085 64321 254113
rect 64349 254085 64383 254113
rect 64411 254085 64459 254113
rect 64149 254051 64459 254085
rect 64149 254023 64197 254051
rect 64225 254023 64259 254051
rect 64287 254023 64321 254051
rect 64349 254023 64383 254051
rect 64411 254023 64459 254051
rect 64149 253989 64459 254023
rect 64149 253961 64197 253989
rect 64225 253961 64259 253989
rect 64287 253961 64321 253989
rect 64349 253961 64383 253989
rect 64411 253961 64459 253989
rect 64149 245175 64459 253961
rect 64149 245147 64197 245175
rect 64225 245147 64259 245175
rect 64287 245147 64321 245175
rect 64349 245147 64383 245175
rect 64411 245147 64459 245175
rect 64149 245113 64459 245147
rect 64149 245085 64197 245113
rect 64225 245085 64259 245113
rect 64287 245085 64321 245113
rect 64349 245085 64383 245113
rect 64411 245085 64459 245113
rect 64149 245051 64459 245085
rect 64149 245023 64197 245051
rect 64225 245023 64259 245051
rect 64287 245023 64321 245051
rect 64349 245023 64383 245051
rect 64411 245023 64459 245051
rect 64149 244989 64459 245023
rect 64149 244961 64197 244989
rect 64225 244961 64259 244989
rect 64287 244961 64321 244989
rect 64349 244961 64383 244989
rect 64411 244961 64459 244989
rect 64149 236175 64459 244961
rect 64149 236147 64197 236175
rect 64225 236147 64259 236175
rect 64287 236147 64321 236175
rect 64349 236147 64383 236175
rect 64411 236147 64459 236175
rect 64149 236113 64459 236147
rect 64149 236085 64197 236113
rect 64225 236085 64259 236113
rect 64287 236085 64321 236113
rect 64349 236085 64383 236113
rect 64411 236085 64459 236113
rect 64149 236051 64459 236085
rect 64149 236023 64197 236051
rect 64225 236023 64259 236051
rect 64287 236023 64321 236051
rect 64349 236023 64383 236051
rect 64411 236023 64459 236051
rect 64149 235989 64459 236023
rect 64149 235961 64197 235989
rect 64225 235961 64259 235989
rect 64287 235961 64321 235989
rect 64349 235961 64383 235989
rect 64411 235961 64459 235989
rect 64149 227175 64459 235961
rect 64149 227147 64197 227175
rect 64225 227147 64259 227175
rect 64287 227147 64321 227175
rect 64349 227147 64383 227175
rect 64411 227147 64459 227175
rect 64149 227113 64459 227147
rect 64149 227085 64197 227113
rect 64225 227085 64259 227113
rect 64287 227085 64321 227113
rect 64349 227085 64383 227113
rect 64411 227085 64459 227113
rect 64149 227051 64459 227085
rect 64149 227023 64197 227051
rect 64225 227023 64259 227051
rect 64287 227023 64321 227051
rect 64349 227023 64383 227051
rect 64411 227023 64459 227051
rect 64149 226989 64459 227023
rect 64149 226961 64197 226989
rect 64225 226961 64259 226989
rect 64287 226961 64321 226989
rect 64349 226961 64383 226989
rect 64411 226961 64459 226989
rect 64149 218175 64459 226961
rect 64149 218147 64197 218175
rect 64225 218147 64259 218175
rect 64287 218147 64321 218175
rect 64349 218147 64383 218175
rect 64411 218147 64459 218175
rect 64149 218113 64459 218147
rect 64149 218085 64197 218113
rect 64225 218085 64259 218113
rect 64287 218085 64321 218113
rect 64349 218085 64383 218113
rect 64411 218085 64459 218113
rect 64149 218051 64459 218085
rect 64149 218023 64197 218051
rect 64225 218023 64259 218051
rect 64287 218023 64321 218051
rect 64349 218023 64383 218051
rect 64411 218023 64459 218051
rect 64149 217989 64459 218023
rect 64149 217961 64197 217989
rect 64225 217961 64259 217989
rect 64287 217961 64321 217989
rect 64349 217961 64383 217989
rect 64411 217961 64459 217989
rect 64149 209175 64459 217961
rect 64149 209147 64197 209175
rect 64225 209147 64259 209175
rect 64287 209147 64321 209175
rect 64349 209147 64383 209175
rect 64411 209147 64459 209175
rect 64149 209113 64459 209147
rect 64149 209085 64197 209113
rect 64225 209085 64259 209113
rect 64287 209085 64321 209113
rect 64349 209085 64383 209113
rect 64411 209085 64459 209113
rect 64149 209051 64459 209085
rect 64149 209023 64197 209051
rect 64225 209023 64259 209051
rect 64287 209023 64321 209051
rect 64349 209023 64383 209051
rect 64411 209023 64459 209051
rect 64149 208989 64459 209023
rect 64149 208961 64197 208989
rect 64225 208961 64259 208989
rect 64287 208961 64321 208989
rect 64349 208961 64383 208989
rect 64411 208961 64459 208989
rect 64149 200175 64459 208961
rect 64149 200147 64197 200175
rect 64225 200147 64259 200175
rect 64287 200147 64321 200175
rect 64349 200147 64383 200175
rect 64411 200147 64459 200175
rect 64149 200113 64459 200147
rect 64149 200085 64197 200113
rect 64225 200085 64259 200113
rect 64287 200085 64321 200113
rect 64349 200085 64383 200113
rect 64411 200085 64459 200113
rect 64149 200051 64459 200085
rect 64149 200023 64197 200051
rect 64225 200023 64259 200051
rect 64287 200023 64321 200051
rect 64349 200023 64383 200051
rect 64411 200023 64459 200051
rect 64149 199989 64459 200023
rect 64149 199961 64197 199989
rect 64225 199961 64259 199989
rect 64287 199961 64321 199989
rect 64349 199961 64383 199989
rect 64411 199961 64459 199989
rect 64149 191175 64459 199961
rect 64149 191147 64197 191175
rect 64225 191147 64259 191175
rect 64287 191147 64321 191175
rect 64349 191147 64383 191175
rect 64411 191147 64459 191175
rect 64149 191113 64459 191147
rect 64149 191085 64197 191113
rect 64225 191085 64259 191113
rect 64287 191085 64321 191113
rect 64349 191085 64383 191113
rect 64411 191085 64459 191113
rect 64149 191051 64459 191085
rect 64149 191023 64197 191051
rect 64225 191023 64259 191051
rect 64287 191023 64321 191051
rect 64349 191023 64383 191051
rect 64411 191023 64459 191051
rect 64149 190989 64459 191023
rect 64149 190961 64197 190989
rect 64225 190961 64259 190989
rect 64287 190961 64321 190989
rect 64349 190961 64383 190989
rect 64411 190961 64459 190989
rect 64149 182175 64459 190961
rect 64149 182147 64197 182175
rect 64225 182147 64259 182175
rect 64287 182147 64321 182175
rect 64349 182147 64383 182175
rect 64411 182147 64459 182175
rect 64149 182113 64459 182147
rect 64149 182085 64197 182113
rect 64225 182085 64259 182113
rect 64287 182085 64321 182113
rect 64349 182085 64383 182113
rect 64411 182085 64459 182113
rect 64149 182051 64459 182085
rect 64149 182023 64197 182051
rect 64225 182023 64259 182051
rect 64287 182023 64321 182051
rect 64349 182023 64383 182051
rect 64411 182023 64459 182051
rect 64149 181989 64459 182023
rect 64149 181961 64197 181989
rect 64225 181961 64259 181989
rect 64287 181961 64321 181989
rect 64349 181961 64383 181989
rect 64411 181961 64459 181989
rect 54304 173175 54464 173192
rect 54304 173147 54339 173175
rect 54367 173147 54401 173175
rect 54429 173147 54464 173175
rect 54304 173113 54464 173147
rect 54304 173085 54339 173113
rect 54367 173085 54401 173113
rect 54429 173085 54464 173113
rect 54304 173051 54464 173085
rect 54304 173023 54339 173051
rect 54367 173023 54401 173051
rect 54429 173023 54464 173051
rect 54304 172989 54464 173023
rect 54304 172961 54339 172989
rect 54367 172961 54401 172989
rect 54429 172961 54464 172989
rect 54304 172944 54464 172961
rect 64149 173175 64459 181961
rect 64149 173147 64197 173175
rect 64225 173147 64259 173175
rect 64287 173147 64321 173175
rect 64349 173147 64383 173175
rect 64411 173147 64459 173175
rect 64149 173113 64459 173147
rect 64149 173085 64197 173113
rect 64225 173085 64259 173113
rect 64287 173085 64321 173113
rect 64349 173085 64383 173113
rect 64411 173085 64459 173113
rect 64149 173051 64459 173085
rect 64149 173023 64197 173051
rect 64225 173023 64259 173051
rect 64287 173023 64321 173051
rect 64349 173023 64383 173051
rect 64411 173023 64459 173051
rect 64149 172989 64459 173023
rect 64149 172961 64197 172989
rect 64225 172961 64259 172989
rect 64287 172961 64321 172989
rect 64349 172961 64383 172989
rect 64411 172961 64459 172989
rect 50649 167147 50697 167175
rect 50725 167147 50759 167175
rect 50787 167147 50821 167175
rect 50849 167147 50883 167175
rect 50911 167147 50959 167175
rect 50649 167113 50959 167147
rect 50649 167085 50697 167113
rect 50725 167085 50759 167113
rect 50787 167085 50821 167113
rect 50849 167085 50883 167113
rect 50911 167085 50959 167113
rect 50649 167051 50959 167085
rect 50649 167023 50697 167051
rect 50725 167023 50759 167051
rect 50787 167023 50821 167051
rect 50849 167023 50883 167051
rect 50911 167023 50959 167051
rect 50649 166989 50959 167023
rect 50649 166961 50697 166989
rect 50725 166961 50759 166989
rect 50787 166961 50821 166989
rect 50849 166961 50883 166989
rect 50911 166961 50959 166989
rect 50649 158175 50959 166961
rect 61984 167175 62144 167192
rect 61984 167147 62019 167175
rect 62047 167147 62081 167175
rect 62109 167147 62144 167175
rect 61984 167113 62144 167147
rect 61984 167085 62019 167113
rect 62047 167085 62081 167113
rect 62109 167085 62144 167113
rect 61984 167051 62144 167085
rect 61984 167023 62019 167051
rect 62047 167023 62081 167051
rect 62109 167023 62144 167051
rect 61984 166989 62144 167023
rect 61984 166961 62019 166989
rect 62047 166961 62081 166989
rect 62109 166961 62144 166989
rect 61984 166944 62144 166961
rect 54304 164175 54464 164192
rect 54304 164147 54339 164175
rect 54367 164147 54401 164175
rect 54429 164147 54464 164175
rect 54304 164113 54464 164147
rect 54304 164085 54339 164113
rect 54367 164085 54401 164113
rect 54429 164085 54464 164113
rect 54304 164051 54464 164085
rect 54304 164023 54339 164051
rect 54367 164023 54401 164051
rect 54429 164023 54464 164051
rect 54304 163989 54464 164023
rect 54304 163961 54339 163989
rect 54367 163961 54401 163989
rect 54429 163961 54464 163989
rect 54304 163944 54464 163961
rect 64149 164175 64459 172961
rect 64149 164147 64197 164175
rect 64225 164147 64259 164175
rect 64287 164147 64321 164175
rect 64349 164147 64383 164175
rect 64411 164147 64459 164175
rect 64149 164113 64459 164147
rect 64149 164085 64197 164113
rect 64225 164085 64259 164113
rect 64287 164085 64321 164113
rect 64349 164085 64383 164113
rect 64411 164085 64459 164113
rect 64149 164051 64459 164085
rect 64149 164023 64197 164051
rect 64225 164023 64259 164051
rect 64287 164023 64321 164051
rect 64349 164023 64383 164051
rect 64411 164023 64459 164051
rect 64149 163989 64459 164023
rect 64149 163961 64197 163989
rect 64225 163961 64259 163989
rect 64287 163961 64321 163989
rect 64349 163961 64383 163989
rect 64411 163961 64459 163989
rect 50649 158147 50697 158175
rect 50725 158147 50759 158175
rect 50787 158147 50821 158175
rect 50849 158147 50883 158175
rect 50911 158147 50959 158175
rect 50649 158113 50959 158147
rect 50649 158085 50697 158113
rect 50725 158085 50759 158113
rect 50787 158085 50821 158113
rect 50849 158085 50883 158113
rect 50911 158085 50959 158113
rect 50649 158051 50959 158085
rect 50649 158023 50697 158051
rect 50725 158023 50759 158051
rect 50787 158023 50821 158051
rect 50849 158023 50883 158051
rect 50911 158023 50959 158051
rect 50649 157989 50959 158023
rect 50649 157961 50697 157989
rect 50725 157961 50759 157989
rect 50787 157961 50821 157989
rect 50849 157961 50883 157989
rect 50911 157961 50959 157989
rect 50649 149175 50959 157961
rect 61984 158175 62144 158192
rect 61984 158147 62019 158175
rect 62047 158147 62081 158175
rect 62109 158147 62144 158175
rect 61984 158113 62144 158147
rect 61984 158085 62019 158113
rect 62047 158085 62081 158113
rect 62109 158085 62144 158113
rect 61984 158051 62144 158085
rect 61984 158023 62019 158051
rect 62047 158023 62081 158051
rect 62109 158023 62144 158051
rect 61984 157989 62144 158023
rect 61984 157961 62019 157989
rect 62047 157961 62081 157989
rect 62109 157961 62144 157989
rect 61984 157944 62144 157961
rect 54304 155175 54464 155192
rect 54304 155147 54339 155175
rect 54367 155147 54401 155175
rect 54429 155147 54464 155175
rect 54304 155113 54464 155147
rect 54304 155085 54339 155113
rect 54367 155085 54401 155113
rect 54429 155085 54464 155113
rect 54304 155051 54464 155085
rect 54304 155023 54339 155051
rect 54367 155023 54401 155051
rect 54429 155023 54464 155051
rect 54304 154989 54464 155023
rect 54304 154961 54339 154989
rect 54367 154961 54401 154989
rect 54429 154961 54464 154989
rect 54304 154944 54464 154961
rect 64149 155175 64459 163961
rect 64149 155147 64197 155175
rect 64225 155147 64259 155175
rect 64287 155147 64321 155175
rect 64349 155147 64383 155175
rect 64411 155147 64459 155175
rect 64149 155113 64459 155147
rect 64149 155085 64197 155113
rect 64225 155085 64259 155113
rect 64287 155085 64321 155113
rect 64349 155085 64383 155113
rect 64411 155085 64459 155113
rect 64149 155051 64459 155085
rect 64149 155023 64197 155051
rect 64225 155023 64259 155051
rect 64287 155023 64321 155051
rect 64349 155023 64383 155051
rect 64411 155023 64459 155051
rect 64149 154989 64459 155023
rect 64149 154961 64197 154989
rect 64225 154961 64259 154989
rect 64287 154961 64321 154989
rect 64349 154961 64383 154989
rect 64411 154961 64459 154989
rect 50649 149147 50697 149175
rect 50725 149147 50759 149175
rect 50787 149147 50821 149175
rect 50849 149147 50883 149175
rect 50911 149147 50959 149175
rect 50649 149113 50959 149147
rect 50649 149085 50697 149113
rect 50725 149085 50759 149113
rect 50787 149085 50821 149113
rect 50849 149085 50883 149113
rect 50911 149085 50959 149113
rect 50649 149051 50959 149085
rect 50649 149023 50697 149051
rect 50725 149023 50759 149051
rect 50787 149023 50821 149051
rect 50849 149023 50883 149051
rect 50911 149023 50959 149051
rect 50649 148989 50959 149023
rect 50649 148961 50697 148989
rect 50725 148961 50759 148989
rect 50787 148961 50821 148989
rect 50849 148961 50883 148989
rect 50911 148961 50959 148989
rect 50649 140175 50959 148961
rect 61984 149175 62144 149192
rect 61984 149147 62019 149175
rect 62047 149147 62081 149175
rect 62109 149147 62144 149175
rect 61984 149113 62144 149147
rect 61984 149085 62019 149113
rect 62047 149085 62081 149113
rect 62109 149085 62144 149113
rect 61984 149051 62144 149085
rect 61984 149023 62019 149051
rect 62047 149023 62081 149051
rect 62109 149023 62144 149051
rect 61984 148989 62144 149023
rect 61984 148961 62019 148989
rect 62047 148961 62081 148989
rect 62109 148961 62144 148989
rect 61984 148944 62144 148961
rect 54304 146175 54464 146192
rect 54304 146147 54339 146175
rect 54367 146147 54401 146175
rect 54429 146147 54464 146175
rect 54304 146113 54464 146147
rect 54304 146085 54339 146113
rect 54367 146085 54401 146113
rect 54429 146085 54464 146113
rect 54304 146051 54464 146085
rect 54304 146023 54339 146051
rect 54367 146023 54401 146051
rect 54429 146023 54464 146051
rect 54304 145989 54464 146023
rect 54304 145961 54339 145989
rect 54367 145961 54401 145989
rect 54429 145961 54464 145989
rect 54304 145944 54464 145961
rect 64149 146175 64459 154961
rect 64149 146147 64197 146175
rect 64225 146147 64259 146175
rect 64287 146147 64321 146175
rect 64349 146147 64383 146175
rect 64411 146147 64459 146175
rect 64149 146113 64459 146147
rect 64149 146085 64197 146113
rect 64225 146085 64259 146113
rect 64287 146085 64321 146113
rect 64349 146085 64383 146113
rect 64411 146085 64459 146113
rect 64149 146051 64459 146085
rect 64149 146023 64197 146051
rect 64225 146023 64259 146051
rect 64287 146023 64321 146051
rect 64349 146023 64383 146051
rect 64411 146023 64459 146051
rect 64149 145989 64459 146023
rect 64149 145961 64197 145989
rect 64225 145961 64259 145989
rect 64287 145961 64321 145989
rect 64349 145961 64383 145989
rect 64411 145961 64459 145989
rect 50649 140147 50697 140175
rect 50725 140147 50759 140175
rect 50787 140147 50821 140175
rect 50849 140147 50883 140175
rect 50911 140147 50959 140175
rect 50649 140113 50959 140147
rect 50649 140085 50697 140113
rect 50725 140085 50759 140113
rect 50787 140085 50821 140113
rect 50849 140085 50883 140113
rect 50911 140085 50959 140113
rect 50649 140051 50959 140085
rect 50649 140023 50697 140051
rect 50725 140023 50759 140051
rect 50787 140023 50821 140051
rect 50849 140023 50883 140051
rect 50911 140023 50959 140051
rect 50649 139989 50959 140023
rect 50649 139961 50697 139989
rect 50725 139961 50759 139989
rect 50787 139961 50821 139989
rect 50849 139961 50883 139989
rect 50911 139961 50959 139989
rect 50649 131175 50959 139961
rect 61984 140175 62144 140192
rect 61984 140147 62019 140175
rect 62047 140147 62081 140175
rect 62109 140147 62144 140175
rect 61984 140113 62144 140147
rect 61984 140085 62019 140113
rect 62047 140085 62081 140113
rect 62109 140085 62144 140113
rect 61984 140051 62144 140085
rect 61984 140023 62019 140051
rect 62047 140023 62081 140051
rect 62109 140023 62144 140051
rect 61984 139989 62144 140023
rect 61984 139961 62019 139989
rect 62047 139961 62081 139989
rect 62109 139961 62144 139989
rect 61984 139944 62144 139961
rect 54304 137175 54464 137192
rect 54304 137147 54339 137175
rect 54367 137147 54401 137175
rect 54429 137147 54464 137175
rect 54304 137113 54464 137147
rect 54304 137085 54339 137113
rect 54367 137085 54401 137113
rect 54429 137085 54464 137113
rect 54304 137051 54464 137085
rect 54304 137023 54339 137051
rect 54367 137023 54401 137051
rect 54429 137023 54464 137051
rect 54304 136989 54464 137023
rect 54304 136961 54339 136989
rect 54367 136961 54401 136989
rect 54429 136961 54464 136989
rect 54304 136944 54464 136961
rect 64149 137175 64459 145961
rect 64149 137147 64197 137175
rect 64225 137147 64259 137175
rect 64287 137147 64321 137175
rect 64349 137147 64383 137175
rect 64411 137147 64459 137175
rect 64149 137113 64459 137147
rect 64149 137085 64197 137113
rect 64225 137085 64259 137113
rect 64287 137085 64321 137113
rect 64349 137085 64383 137113
rect 64411 137085 64459 137113
rect 64149 137051 64459 137085
rect 64149 137023 64197 137051
rect 64225 137023 64259 137051
rect 64287 137023 64321 137051
rect 64349 137023 64383 137051
rect 64411 137023 64459 137051
rect 64149 136989 64459 137023
rect 64149 136961 64197 136989
rect 64225 136961 64259 136989
rect 64287 136961 64321 136989
rect 64349 136961 64383 136989
rect 64411 136961 64459 136989
rect 50649 131147 50697 131175
rect 50725 131147 50759 131175
rect 50787 131147 50821 131175
rect 50849 131147 50883 131175
rect 50911 131147 50959 131175
rect 50649 131113 50959 131147
rect 50649 131085 50697 131113
rect 50725 131085 50759 131113
rect 50787 131085 50821 131113
rect 50849 131085 50883 131113
rect 50911 131085 50959 131113
rect 50649 131051 50959 131085
rect 50649 131023 50697 131051
rect 50725 131023 50759 131051
rect 50787 131023 50821 131051
rect 50849 131023 50883 131051
rect 50911 131023 50959 131051
rect 50649 130989 50959 131023
rect 50649 130961 50697 130989
rect 50725 130961 50759 130989
rect 50787 130961 50821 130989
rect 50849 130961 50883 130989
rect 50911 130961 50959 130989
rect 50649 122175 50959 130961
rect 61984 131175 62144 131192
rect 61984 131147 62019 131175
rect 62047 131147 62081 131175
rect 62109 131147 62144 131175
rect 61984 131113 62144 131147
rect 61984 131085 62019 131113
rect 62047 131085 62081 131113
rect 62109 131085 62144 131113
rect 61984 131051 62144 131085
rect 61984 131023 62019 131051
rect 62047 131023 62081 131051
rect 62109 131023 62144 131051
rect 61984 130989 62144 131023
rect 61984 130961 62019 130989
rect 62047 130961 62081 130989
rect 62109 130961 62144 130989
rect 61984 130944 62144 130961
rect 54304 128175 54464 128192
rect 54304 128147 54339 128175
rect 54367 128147 54401 128175
rect 54429 128147 54464 128175
rect 54304 128113 54464 128147
rect 54304 128085 54339 128113
rect 54367 128085 54401 128113
rect 54429 128085 54464 128113
rect 54304 128051 54464 128085
rect 54304 128023 54339 128051
rect 54367 128023 54401 128051
rect 54429 128023 54464 128051
rect 54304 127989 54464 128023
rect 54304 127961 54339 127989
rect 54367 127961 54401 127989
rect 54429 127961 54464 127989
rect 54304 127944 54464 127961
rect 64149 128175 64459 136961
rect 64149 128147 64197 128175
rect 64225 128147 64259 128175
rect 64287 128147 64321 128175
rect 64349 128147 64383 128175
rect 64411 128147 64459 128175
rect 64149 128113 64459 128147
rect 64149 128085 64197 128113
rect 64225 128085 64259 128113
rect 64287 128085 64321 128113
rect 64349 128085 64383 128113
rect 64411 128085 64459 128113
rect 64149 128051 64459 128085
rect 64149 128023 64197 128051
rect 64225 128023 64259 128051
rect 64287 128023 64321 128051
rect 64349 128023 64383 128051
rect 64411 128023 64459 128051
rect 64149 127989 64459 128023
rect 64149 127961 64197 127989
rect 64225 127961 64259 127989
rect 64287 127961 64321 127989
rect 64349 127961 64383 127989
rect 64411 127961 64459 127989
rect 50649 122147 50697 122175
rect 50725 122147 50759 122175
rect 50787 122147 50821 122175
rect 50849 122147 50883 122175
rect 50911 122147 50959 122175
rect 50649 122113 50959 122147
rect 50649 122085 50697 122113
rect 50725 122085 50759 122113
rect 50787 122085 50821 122113
rect 50849 122085 50883 122113
rect 50911 122085 50959 122113
rect 50649 122051 50959 122085
rect 50649 122023 50697 122051
rect 50725 122023 50759 122051
rect 50787 122023 50821 122051
rect 50849 122023 50883 122051
rect 50911 122023 50959 122051
rect 50649 121989 50959 122023
rect 50649 121961 50697 121989
rect 50725 121961 50759 121989
rect 50787 121961 50821 121989
rect 50849 121961 50883 121989
rect 50911 121961 50959 121989
rect 50649 113175 50959 121961
rect 61984 122175 62144 122192
rect 61984 122147 62019 122175
rect 62047 122147 62081 122175
rect 62109 122147 62144 122175
rect 61984 122113 62144 122147
rect 61984 122085 62019 122113
rect 62047 122085 62081 122113
rect 62109 122085 62144 122113
rect 61984 122051 62144 122085
rect 61984 122023 62019 122051
rect 62047 122023 62081 122051
rect 62109 122023 62144 122051
rect 61984 121989 62144 122023
rect 61984 121961 62019 121989
rect 62047 121961 62081 121989
rect 62109 121961 62144 121989
rect 61984 121944 62144 121961
rect 54304 119175 54464 119192
rect 54304 119147 54339 119175
rect 54367 119147 54401 119175
rect 54429 119147 54464 119175
rect 54304 119113 54464 119147
rect 54304 119085 54339 119113
rect 54367 119085 54401 119113
rect 54429 119085 54464 119113
rect 54304 119051 54464 119085
rect 54304 119023 54339 119051
rect 54367 119023 54401 119051
rect 54429 119023 54464 119051
rect 54304 118989 54464 119023
rect 54304 118961 54339 118989
rect 54367 118961 54401 118989
rect 54429 118961 54464 118989
rect 54304 118944 54464 118961
rect 64149 119175 64459 127961
rect 64149 119147 64197 119175
rect 64225 119147 64259 119175
rect 64287 119147 64321 119175
rect 64349 119147 64383 119175
rect 64411 119147 64459 119175
rect 64149 119113 64459 119147
rect 64149 119085 64197 119113
rect 64225 119085 64259 119113
rect 64287 119085 64321 119113
rect 64349 119085 64383 119113
rect 64411 119085 64459 119113
rect 64149 119051 64459 119085
rect 64149 119023 64197 119051
rect 64225 119023 64259 119051
rect 64287 119023 64321 119051
rect 64349 119023 64383 119051
rect 64411 119023 64459 119051
rect 64149 118989 64459 119023
rect 64149 118961 64197 118989
rect 64225 118961 64259 118989
rect 64287 118961 64321 118989
rect 64349 118961 64383 118989
rect 64411 118961 64459 118989
rect 50649 113147 50697 113175
rect 50725 113147 50759 113175
rect 50787 113147 50821 113175
rect 50849 113147 50883 113175
rect 50911 113147 50959 113175
rect 50649 113113 50959 113147
rect 50649 113085 50697 113113
rect 50725 113085 50759 113113
rect 50787 113085 50821 113113
rect 50849 113085 50883 113113
rect 50911 113085 50959 113113
rect 50649 113051 50959 113085
rect 50649 113023 50697 113051
rect 50725 113023 50759 113051
rect 50787 113023 50821 113051
rect 50849 113023 50883 113051
rect 50911 113023 50959 113051
rect 50649 112989 50959 113023
rect 50649 112961 50697 112989
rect 50725 112961 50759 112989
rect 50787 112961 50821 112989
rect 50849 112961 50883 112989
rect 50911 112961 50959 112989
rect 50649 104175 50959 112961
rect 61984 113175 62144 113192
rect 61984 113147 62019 113175
rect 62047 113147 62081 113175
rect 62109 113147 62144 113175
rect 61984 113113 62144 113147
rect 61984 113085 62019 113113
rect 62047 113085 62081 113113
rect 62109 113085 62144 113113
rect 61984 113051 62144 113085
rect 61984 113023 62019 113051
rect 62047 113023 62081 113051
rect 62109 113023 62144 113051
rect 61984 112989 62144 113023
rect 61984 112961 62019 112989
rect 62047 112961 62081 112989
rect 62109 112961 62144 112989
rect 61984 112944 62144 112961
rect 54304 110175 54464 110192
rect 54304 110147 54339 110175
rect 54367 110147 54401 110175
rect 54429 110147 54464 110175
rect 54304 110113 54464 110147
rect 54304 110085 54339 110113
rect 54367 110085 54401 110113
rect 54429 110085 54464 110113
rect 54304 110051 54464 110085
rect 54304 110023 54339 110051
rect 54367 110023 54401 110051
rect 54429 110023 54464 110051
rect 54304 109989 54464 110023
rect 54304 109961 54339 109989
rect 54367 109961 54401 109989
rect 54429 109961 54464 109989
rect 54304 109944 54464 109961
rect 64149 110175 64459 118961
rect 64149 110147 64197 110175
rect 64225 110147 64259 110175
rect 64287 110147 64321 110175
rect 64349 110147 64383 110175
rect 64411 110147 64459 110175
rect 64149 110113 64459 110147
rect 64149 110085 64197 110113
rect 64225 110085 64259 110113
rect 64287 110085 64321 110113
rect 64349 110085 64383 110113
rect 64411 110085 64459 110113
rect 64149 110051 64459 110085
rect 64149 110023 64197 110051
rect 64225 110023 64259 110051
rect 64287 110023 64321 110051
rect 64349 110023 64383 110051
rect 64411 110023 64459 110051
rect 64149 109989 64459 110023
rect 64149 109961 64197 109989
rect 64225 109961 64259 109989
rect 64287 109961 64321 109989
rect 64349 109961 64383 109989
rect 64411 109961 64459 109989
rect 50649 104147 50697 104175
rect 50725 104147 50759 104175
rect 50787 104147 50821 104175
rect 50849 104147 50883 104175
rect 50911 104147 50959 104175
rect 50649 104113 50959 104147
rect 50649 104085 50697 104113
rect 50725 104085 50759 104113
rect 50787 104085 50821 104113
rect 50849 104085 50883 104113
rect 50911 104085 50959 104113
rect 50649 104051 50959 104085
rect 50649 104023 50697 104051
rect 50725 104023 50759 104051
rect 50787 104023 50821 104051
rect 50849 104023 50883 104051
rect 50911 104023 50959 104051
rect 50649 103989 50959 104023
rect 50649 103961 50697 103989
rect 50725 103961 50759 103989
rect 50787 103961 50821 103989
rect 50849 103961 50883 103989
rect 50911 103961 50959 103989
rect 50649 95175 50959 103961
rect 61984 104175 62144 104192
rect 61984 104147 62019 104175
rect 62047 104147 62081 104175
rect 62109 104147 62144 104175
rect 61984 104113 62144 104147
rect 61984 104085 62019 104113
rect 62047 104085 62081 104113
rect 62109 104085 62144 104113
rect 61984 104051 62144 104085
rect 61984 104023 62019 104051
rect 62047 104023 62081 104051
rect 62109 104023 62144 104051
rect 61984 103989 62144 104023
rect 61984 103961 62019 103989
rect 62047 103961 62081 103989
rect 62109 103961 62144 103989
rect 61984 103944 62144 103961
rect 54304 101175 54464 101192
rect 54304 101147 54339 101175
rect 54367 101147 54401 101175
rect 54429 101147 54464 101175
rect 54304 101113 54464 101147
rect 54304 101085 54339 101113
rect 54367 101085 54401 101113
rect 54429 101085 54464 101113
rect 54304 101051 54464 101085
rect 54304 101023 54339 101051
rect 54367 101023 54401 101051
rect 54429 101023 54464 101051
rect 54304 100989 54464 101023
rect 54304 100961 54339 100989
rect 54367 100961 54401 100989
rect 54429 100961 54464 100989
rect 54304 100944 54464 100961
rect 64149 101175 64459 109961
rect 64149 101147 64197 101175
rect 64225 101147 64259 101175
rect 64287 101147 64321 101175
rect 64349 101147 64383 101175
rect 64411 101147 64459 101175
rect 64149 101113 64459 101147
rect 64149 101085 64197 101113
rect 64225 101085 64259 101113
rect 64287 101085 64321 101113
rect 64349 101085 64383 101113
rect 64411 101085 64459 101113
rect 64149 101051 64459 101085
rect 64149 101023 64197 101051
rect 64225 101023 64259 101051
rect 64287 101023 64321 101051
rect 64349 101023 64383 101051
rect 64411 101023 64459 101051
rect 64149 100989 64459 101023
rect 64149 100961 64197 100989
rect 64225 100961 64259 100989
rect 64287 100961 64321 100989
rect 64349 100961 64383 100989
rect 64411 100961 64459 100989
rect 50649 95147 50697 95175
rect 50725 95147 50759 95175
rect 50787 95147 50821 95175
rect 50849 95147 50883 95175
rect 50911 95147 50959 95175
rect 50649 95113 50959 95147
rect 50649 95085 50697 95113
rect 50725 95085 50759 95113
rect 50787 95085 50821 95113
rect 50849 95085 50883 95113
rect 50911 95085 50959 95113
rect 50649 95051 50959 95085
rect 50649 95023 50697 95051
rect 50725 95023 50759 95051
rect 50787 95023 50821 95051
rect 50849 95023 50883 95051
rect 50911 95023 50959 95051
rect 50649 94989 50959 95023
rect 50649 94961 50697 94989
rect 50725 94961 50759 94989
rect 50787 94961 50821 94989
rect 50849 94961 50883 94989
rect 50911 94961 50959 94989
rect 50649 86175 50959 94961
rect 61984 95175 62144 95192
rect 61984 95147 62019 95175
rect 62047 95147 62081 95175
rect 62109 95147 62144 95175
rect 61984 95113 62144 95147
rect 61984 95085 62019 95113
rect 62047 95085 62081 95113
rect 62109 95085 62144 95113
rect 61984 95051 62144 95085
rect 61984 95023 62019 95051
rect 62047 95023 62081 95051
rect 62109 95023 62144 95051
rect 61984 94989 62144 95023
rect 61984 94961 62019 94989
rect 62047 94961 62081 94989
rect 62109 94961 62144 94989
rect 61984 94944 62144 94961
rect 54304 92175 54464 92192
rect 54304 92147 54339 92175
rect 54367 92147 54401 92175
rect 54429 92147 54464 92175
rect 54304 92113 54464 92147
rect 54304 92085 54339 92113
rect 54367 92085 54401 92113
rect 54429 92085 54464 92113
rect 54304 92051 54464 92085
rect 54304 92023 54339 92051
rect 54367 92023 54401 92051
rect 54429 92023 54464 92051
rect 54304 91989 54464 92023
rect 54304 91961 54339 91989
rect 54367 91961 54401 91989
rect 54429 91961 54464 91989
rect 54304 91944 54464 91961
rect 64149 92175 64459 100961
rect 64149 92147 64197 92175
rect 64225 92147 64259 92175
rect 64287 92147 64321 92175
rect 64349 92147 64383 92175
rect 64411 92147 64459 92175
rect 64149 92113 64459 92147
rect 64149 92085 64197 92113
rect 64225 92085 64259 92113
rect 64287 92085 64321 92113
rect 64349 92085 64383 92113
rect 64411 92085 64459 92113
rect 64149 92051 64459 92085
rect 64149 92023 64197 92051
rect 64225 92023 64259 92051
rect 64287 92023 64321 92051
rect 64349 92023 64383 92051
rect 64411 92023 64459 92051
rect 64149 91989 64459 92023
rect 64149 91961 64197 91989
rect 64225 91961 64259 91989
rect 64287 91961 64321 91989
rect 64349 91961 64383 91989
rect 64411 91961 64459 91989
rect 50649 86147 50697 86175
rect 50725 86147 50759 86175
rect 50787 86147 50821 86175
rect 50849 86147 50883 86175
rect 50911 86147 50959 86175
rect 50649 86113 50959 86147
rect 50649 86085 50697 86113
rect 50725 86085 50759 86113
rect 50787 86085 50821 86113
rect 50849 86085 50883 86113
rect 50911 86085 50959 86113
rect 50649 86051 50959 86085
rect 50649 86023 50697 86051
rect 50725 86023 50759 86051
rect 50787 86023 50821 86051
rect 50849 86023 50883 86051
rect 50911 86023 50959 86051
rect 50649 85989 50959 86023
rect 50649 85961 50697 85989
rect 50725 85961 50759 85989
rect 50787 85961 50821 85989
rect 50849 85961 50883 85989
rect 50911 85961 50959 85989
rect 50649 77175 50959 85961
rect 61984 86175 62144 86192
rect 61984 86147 62019 86175
rect 62047 86147 62081 86175
rect 62109 86147 62144 86175
rect 61984 86113 62144 86147
rect 61984 86085 62019 86113
rect 62047 86085 62081 86113
rect 62109 86085 62144 86113
rect 61984 86051 62144 86085
rect 61984 86023 62019 86051
rect 62047 86023 62081 86051
rect 62109 86023 62144 86051
rect 61984 85989 62144 86023
rect 61984 85961 62019 85989
rect 62047 85961 62081 85989
rect 62109 85961 62144 85989
rect 61984 85944 62144 85961
rect 54304 83175 54464 83192
rect 54304 83147 54339 83175
rect 54367 83147 54401 83175
rect 54429 83147 54464 83175
rect 54304 83113 54464 83147
rect 54304 83085 54339 83113
rect 54367 83085 54401 83113
rect 54429 83085 54464 83113
rect 54304 83051 54464 83085
rect 54304 83023 54339 83051
rect 54367 83023 54401 83051
rect 54429 83023 54464 83051
rect 54304 82989 54464 83023
rect 54304 82961 54339 82989
rect 54367 82961 54401 82989
rect 54429 82961 54464 82989
rect 54304 82944 54464 82961
rect 64149 83175 64459 91961
rect 64149 83147 64197 83175
rect 64225 83147 64259 83175
rect 64287 83147 64321 83175
rect 64349 83147 64383 83175
rect 64411 83147 64459 83175
rect 64149 83113 64459 83147
rect 64149 83085 64197 83113
rect 64225 83085 64259 83113
rect 64287 83085 64321 83113
rect 64349 83085 64383 83113
rect 64411 83085 64459 83113
rect 64149 83051 64459 83085
rect 64149 83023 64197 83051
rect 64225 83023 64259 83051
rect 64287 83023 64321 83051
rect 64349 83023 64383 83051
rect 64411 83023 64459 83051
rect 64149 82989 64459 83023
rect 64149 82961 64197 82989
rect 64225 82961 64259 82989
rect 64287 82961 64321 82989
rect 64349 82961 64383 82989
rect 64411 82961 64459 82989
rect 50649 77147 50697 77175
rect 50725 77147 50759 77175
rect 50787 77147 50821 77175
rect 50849 77147 50883 77175
rect 50911 77147 50959 77175
rect 50649 77113 50959 77147
rect 50649 77085 50697 77113
rect 50725 77085 50759 77113
rect 50787 77085 50821 77113
rect 50849 77085 50883 77113
rect 50911 77085 50959 77113
rect 50649 77051 50959 77085
rect 50649 77023 50697 77051
rect 50725 77023 50759 77051
rect 50787 77023 50821 77051
rect 50849 77023 50883 77051
rect 50911 77023 50959 77051
rect 50649 76989 50959 77023
rect 50649 76961 50697 76989
rect 50725 76961 50759 76989
rect 50787 76961 50821 76989
rect 50849 76961 50883 76989
rect 50911 76961 50959 76989
rect 50649 68175 50959 76961
rect 61984 77175 62144 77192
rect 61984 77147 62019 77175
rect 62047 77147 62081 77175
rect 62109 77147 62144 77175
rect 61984 77113 62144 77147
rect 61984 77085 62019 77113
rect 62047 77085 62081 77113
rect 62109 77085 62144 77113
rect 61984 77051 62144 77085
rect 61984 77023 62019 77051
rect 62047 77023 62081 77051
rect 62109 77023 62144 77051
rect 61984 76989 62144 77023
rect 61984 76961 62019 76989
rect 62047 76961 62081 76989
rect 62109 76961 62144 76989
rect 61984 76944 62144 76961
rect 54304 74175 54464 74192
rect 54304 74147 54339 74175
rect 54367 74147 54401 74175
rect 54429 74147 54464 74175
rect 54304 74113 54464 74147
rect 54304 74085 54339 74113
rect 54367 74085 54401 74113
rect 54429 74085 54464 74113
rect 54304 74051 54464 74085
rect 54304 74023 54339 74051
rect 54367 74023 54401 74051
rect 54429 74023 54464 74051
rect 54304 73989 54464 74023
rect 54304 73961 54339 73989
rect 54367 73961 54401 73989
rect 54429 73961 54464 73989
rect 54304 73944 54464 73961
rect 64149 74175 64459 82961
rect 64149 74147 64197 74175
rect 64225 74147 64259 74175
rect 64287 74147 64321 74175
rect 64349 74147 64383 74175
rect 64411 74147 64459 74175
rect 64149 74113 64459 74147
rect 64149 74085 64197 74113
rect 64225 74085 64259 74113
rect 64287 74085 64321 74113
rect 64349 74085 64383 74113
rect 64411 74085 64459 74113
rect 64149 74051 64459 74085
rect 64149 74023 64197 74051
rect 64225 74023 64259 74051
rect 64287 74023 64321 74051
rect 64349 74023 64383 74051
rect 64411 74023 64459 74051
rect 64149 73989 64459 74023
rect 64149 73961 64197 73989
rect 64225 73961 64259 73989
rect 64287 73961 64321 73989
rect 64349 73961 64383 73989
rect 64411 73961 64459 73989
rect 50649 68147 50697 68175
rect 50725 68147 50759 68175
rect 50787 68147 50821 68175
rect 50849 68147 50883 68175
rect 50911 68147 50959 68175
rect 50649 68113 50959 68147
rect 50649 68085 50697 68113
rect 50725 68085 50759 68113
rect 50787 68085 50821 68113
rect 50849 68085 50883 68113
rect 50911 68085 50959 68113
rect 50649 68051 50959 68085
rect 50649 68023 50697 68051
rect 50725 68023 50759 68051
rect 50787 68023 50821 68051
rect 50849 68023 50883 68051
rect 50911 68023 50959 68051
rect 50649 67989 50959 68023
rect 50649 67961 50697 67989
rect 50725 67961 50759 67989
rect 50787 67961 50821 67989
rect 50849 67961 50883 67989
rect 50911 67961 50959 67989
rect 50649 59175 50959 67961
rect 61984 68175 62144 68192
rect 61984 68147 62019 68175
rect 62047 68147 62081 68175
rect 62109 68147 62144 68175
rect 61984 68113 62144 68147
rect 61984 68085 62019 68113
rect 62047 68085 62081 68113
rect 62109 68085 62144 68113
rect 61984 68051 62144 68085
rect 61984 68023 62019 68051
rect 62047 68023 62081 68051
rect 62109 68023 62144 68051
rect 61984 67989 62144 68023
rect 61984 67961 62019 67989
rect 62047 67961 62081 67989
rect 62109 67961 62144 67989
rect 61984 67944 62144 67961
rect 54304 65175 54464 65192
rect 54304 65147 54339 65175
rect 54367 65147 54401 65175
rect 54429 65147 54464 65175
rect 54304 65113 54464 65147
rect 54304 65085 54339 65113
rect 54367 65085 54401 65113
rect 54429 65085 54464 65113
rect 54304 65051 54464 65085
rect 54304 65023 54339 65051
rect 54367 65023 54401 65051
rect 54429 65023 54464 65051
rect 54304 64989 54464 65023
rect 54304 64961 54339 64989
rect 54367 64961 54401 64989
rect 54429 64961 54464 64989
rect 54304 64944 54464 64961
rect 64149 65175 64459 73961
rect 64149 65147 64197 65175
rect 64225 65147 64259 65175
rect 64287 65147 64321 65175
rect 64349 65147 64383 65175
rect 64411 65147 64459 65175
rect 64149 65113 64459 65147
rect 64149 65085 64197 65113
rect 64225 65085 64259 65113
rect 64287 65085 64321 65113
rect 64349 65085 64383 65113
rect 64411 65085 64459 65113
rect 64149 65051 64459 65085
rect 64149 65023 64197 65051
rect 64225 65023 64259 65051
rect 64287 65023 64321 65051
rect 64349 65023 64383 65051
rect 64411 65023 64459 65051
rect 64149 64989 64459 65023
rect 64149 64961 64197 64989
rect 64225 64961 64259 64989
rect 64287 64961 64321 64989
rect 64349 64961 64383 64989
rect 64411 64961 64459 64989
rect 50649 59147 50697 59175
rect 50725 59147 50759 59175
rect 50787 59147 50821 59175
rect 50849 59147 50883 59175
rect 50911 59147 50959 59175
rect 50649 59113 50959 59147
rect 50649 59085 50697 59113
rect 50725 59085 50759 59113
rect 50787 59085 50821 59113
rect 50849 59085 50883 59113
rect 50911 59085 50959 59113
rect 50649 59051 50959 59085
rect 50649 59023 50697 59051
rect 50725 59023 50759 59051
rect 50787 59023 50821 59051
rect 50849 59023 50883 59051
rect 50911 59023 50959 59051
rect 50649 58989 50959 59023
rect 50649 58961 50697 58989
rect 50725 58961 50759 58989
rect 50787 58961 50821 58989
rect 50849 58961 50883 58989
rect 50911 58961 50959 58989
rect 50649 50175 50959 58961
rect 61984 59175 62144 59192
rect 61984 59147 62019 59175
rect 62047 59147 62081 59175
rect 62109 59147 62144 59175
rect 61984 59113 62144 59147
rect 61984 59085 62019 59113
rect 62047 59085 62081 59113
rect 62109 59085 62144 59113
rect 61984 59051 62144 59085
rect 61984 59023 62019 59051
rect 62047 59023 62081 59051
rect 62109 59023 62144 59051
rect 61984 58989 62144 59023
rect 61984 58961 62019 58989
rect 62047 58961 62081 58989
rect 62109 58961 62144 58989
rect 61984 58944 62144 58961
rect 54304 56175 54464 56192
rect 54304 56147 54339 56175
rect 54367 56147 54401 56175
rect 54429 56147 54464 56175
rect 54304 56113 54464 56147
rect 54304 56085 54339 56113
rect 54367 56085 54401 56113
rect 54429 56085 54464 56113
rect 54304 56051 54464 56085
rect 54304 56023 54339 56051
rect 54367 56023 54401 56051
rect 54429 56023 54464 56051
rect 54304 55989 54464 56023
rect 54304 55961 54339 55989
rect 54367 55961 54401 55989
rect 54429 55961 54464 55989
rect 54304 55944 54464 55961
rect 64149 56175 64459 64961
rect 64149 56147 64197 56175
rect 64225 56147 64259 56175
rect 64287 56147 64321 56175
rect 64349 56147 64383 56175
rect 64411 56147 64459 56175
rect 64149 56113 64459 56147
rect 64149 56085 64197 56113
rect 64225 56085 64259 56113
rect 64287 56085 64321 56113
rect 64349 56085 64383 56113
rect 64411 56085 64459 56113
rect 64149 56051 64459 56085
rect 64149 56023 64197 56051
rect 64225 56023 64259 56051
rect 64287 56023 64321 56051
rect 64349 56023 64383 56051
rect 64411 56023 64459 56051
rect 64149 55989 64459 56023
rect 64149 55961 64197 55989
rect 64225 55961 64259 55989
rect 64287 55961 64321 55989
rect 64349 55961 64383 55989
rect 64411 55961 64459 55989
rect 50649 50147 50697 50175
rect 50725 50147 50759 50175
rect 50787 50147 50821 50175
rect 50849 50147 50883 50175
rect 50911 50147 50959 50175
rect 50649 50113 50959 50147
rect 50649 50085 50697 50113
rect 50725 50085 50759 50113
rect 50787 50085 50821 50113
rect 50849 50085 50883 50113
rect 50911 50085 50959 50113
rect 50649 50051 50959 50085
rect 50649 50023 50697 50051
rect 50725 50023 50759 50051
rect 50787 50023 50821 50051
rect 50849 50023 50883 50051
rect 50911 50023 50959 50051
rect 50649 49989 50959 50023
rect 50649 49961 50697 49989
rect 50725 49961 50759 49989
rect 50787 49961 50821 49989
rect 50849 49961 50883 49989
rect 50911 49961 50959 49989
rect 50649 41175 50959 49961
rect 61984 50175 62144 50192
rect 61984 50147 62019 50175
rect 62047 50147 62081 50175
rect 62109 50147 62144 50175
rect 61984 50113 62144 50147
rect 61984 50085 62019 50113
rect 62047 50085 62081 50113
rect 62109 50085 62144 50113
rect 61984 50051 62144 50085
rect 61984 50023 62019 50051
rect 62047 50023 62081 50051
rect 62109 50023 62144 50051
rect 61984 49989 62144 50023
rect 61984 49961 62019 49989
rect 62047 49961 62081 49989
rect 62109 49961 62144 49989
rect 61984 49944 62144 49961
rect 54304 47175 54464 47192
rect 54304 47147 54339 47175
rect 54367 47147 54401 47175
rect 54429 47147 54464 47175
rect 54304 47113 54464 47147
rect 54304 47085 54339 47113
rect 54367 47085 54401 47113
rect 54429 47085 54464 47113
rect 54304 47051 54464 47085
rect 54304 47023 54339 47051
rect 54367 47023 54401 47051
rect 54429 47023 54464 47051
rect 54304 46989 54464 47023
rect 54304 46961 54339 46989
rect 54367 46961 54401 46989
rect 54429 46961 54464 46989
rect 54304 46944 54464 46961
rect 64149 47175 64459 55961
rect 64149 47147 64197 47175
rect 64225 47147 64259 47175
rect 64287 47147 64321 47175
rect 64349 47147 64383 47175
rect 64411 47147 64459 47175
rect 64149 47113 64459 47147
rect 64149 47085 64197 47113
rect 64225 47085 64259 47113
rect 64287 47085 64321 47113
rect 64349 47085 64383 47113
rect 64411 47085 64459 47113
rect 64149 47051 64459 47085
rect 64149 47023 64197 47051
rect 64225 47023 64259 47051
rect 64287 47023 64321 47051
rect 64349 47023 64383 47051
rect 64411 47023 64459 47051
rect 64149 46989 64459 47023
rect 64149 46961 64197 46989
rect 64225 46961 64259 46989
rect 64287 46961 64321 46989
rect 64349 46961 64383 46989
rect 64411 46961 64459 46989
rect 50649 41147 50697 41175
rect 50725 41147 50759 41175
rect 50787 41147 50821 41175
rect 50849 41147 50883 41175
rect 50911 41147 50959 41175
rect 50649 41113 50959 41147
rect 50649 41085 50697 41113
rect 50725 41085 50759 41113
rect 50787 41085 50821 41113
rect 50849 41085 50883 41113
rect 50911 41085 50959 41113
rect 50649 41051 50959 41085
rect 50649 41023 50697 41051
rect 50725 41023 50759 41051
rect 50787 41023 50821 41051
rect 50849 41023 50883 41051
rect 50911 41023 50959 41051
rect 50649 40989 50959 41023
rect 50649 40961 50697 40989
rect 50725 40961 50759 40989
rect 50787 40961 50821 40989
rect 50849 40961 50883 40989
rect 50911 40961 50959 40989
rect 50649 32175 50959 40961
rect 61984 41175 62144 41192
rect 61984 41147 62019 41175
rect 62047 41147 62081 41175
rect 62109 41147 62144 41175
rect 61984 41113 62144 41147
rect 61984 41085 62019 41113
rect 62047 41085 62081 41113
rect 62109 41085 62144 41113
rect 61984 41051 62144 41085
rect 61984 41023 62019 41051
rect 62047 41023 62081 41051
rect 62109 41023 62144 41051
rect 61984 40989 62144 41023
rect 61984 40961 62019 40989
rect 62047 40961 62081 40989
rect 62109 40961 62144 40989
rect 61984 40944 62144 40961
rect 54304 38175 54464 38192
rect 54304 38147 54339 38175
rect 54367 38147 54401 38175
rect 54429 38147 54464 38175
rect 54304 38113 54464 38147
rect 54304 38085 54339 38113
rect 54367 38085 54401 38113
rect 54429 38085 54464 38113
rect 54304 38051 54464 38085
rect 54304 38023 54339 38051
rect 54367 38023 54401 38051
rect 54429 38023 54464 38051
rect 54304 37989 54464 38023
rect 54304 37961 54339 37989
rect 54367 37961 54401 37989
rect 54429 37961 54464 37989
rect 54304 37944 54464 37961
rect 64149 38175 64459 46961
rect 64149 38147 64197 38175
rect 64225 38147 64259 38175
rect 64287 38147 64321 38175
rect 64349 38147 64383 38175
rect 64411 38147 64459 38175
rect 64149 38113 64459 38147
rect 64149 38085 64197 38113
rect 64225 38085 64259 38113
rect 64287 38085 64321 38113
rect 64349 38085 64383 38113
rect 64411 38085 64459 38113
rect 64149 38051 64459 38085
rect 64149 38023 64197 38051
rect 64225 38023 64259 38051
rect 64287 38023 64321 38051
rect 64349 38023 64383 38051
rect 64411 38023 64459 38051
rect 64149 37989 64459 38023
rect 64149 37961 64197 37989
rect 64225 37961 64259 37989
rect 64287 37961 64321 37989
rect 64349 37961 64383 37989
rect 64411 37961 64459 37989
rect 50649 32147 50697 32175
rect 50725 32147 50759 32175
rect 50787 32147 50821 32175
rect 50849 32147 50883 32175
rect 50911 32147 50959 32175
rect 50649 32113 50959 32147
rect 50649 32085 50697 32113
rect 50725 32085 50759 32113
rect 50787 32085 50821 32113
rect 50849 32085 50883 32113
rect 50911 32085 50959 32113
rect 50649 32051 50959 32085
rect 50649 32023 50697 32051
rect 50725 32023 50759 32051
rect 50787 32023 50821 32051
rect 50849 32023 50883 32051
rect 50911 32023 50959 32051
rect 50649 31989 50959 32023
rect 50649 31961 50697 31989
rect 50725 31961 50759 31989
rect 50787 31961 50821 31989
rect 50849 31961 50883 31989
rect 50911 31961 50959 31989
rect 50649 23175 50959 31961
rect 61984 32175 62144 32192
rect 61984 32147 62019 32175
rect 62047 32147 62081 32175
rect 62109 32147 62144 32175
rect 61984 32113 62144 32147
rect 61984 32085 62019 32113
rect 62047 32085 62081 32113
rect 62109 32085 62144 32113
rect 61984 32051 62144 32085
rect 61984 32023 62019 32051
rect 62047 32023 62081 32051
rect 62109 32023 62144 32051
rect 61984 31989 62144 32023
rect 61984 31961 62019 31989
rect 62047 31961 62081 31989
rect 62109 31961 62144 31989
rect 61984 31944 62144 31961
rect 54304 29175 54464 29192
rect 54304 29147 54339 29175
rect 54367 29147 54401 29175
rect 54429 29147 54464 29175
rect 54304 29113 54464 29147
rect 54304 29085 54339 29113
rect 54367 29085 54401 29113
rect 54429 29085 54464 29113
rect 54304 29051 54464 29085
rect 54304 29023 54339 29051
rect 54367 29023 54401 29051
rect 54429 29023 54464 29051
rect 54304 28989 54464 29023
rect 54304 28961 54339 28989
rect 54367 28961 54401 28989
rect 54429 28961 54464 28989
rect 54304 28944 54464 28961
rect 64149 29175 64459 37961
rect 64149 29147 64197 29175
rect 64225 29147 64259 29175
rect 64287 29147 64321 29175
rect 64349 29147 64383 29175
rect 64411 29147 64459 29175
rect 64149 29113 64459 29147
rect 64149 29085 64197 29113
rect 64225 29085 64259 29113
rect 64287 29085 64321 29113
rect 64349 29085 64383 29113
rect 64411 29085 64459 29113
rect 64149 29051 64459 29085
rect 64149 29023 64197 29051
rect 64225 29023 64259 29051
rect 64287 29023 64321 29051
rect 64349 29023 64383 29051
rect 64411 29023 64459 29051
rect 64149 28989 64459 29023
rect 64149 28961 64197 28989
rect 64225 28961 64259 28989
rect 64287 28961 64321 28989
rect 64349 28961 64383 28989
rect 64411 28961 64459 28989
rect 50649 23147 50697 23175
rect 50725 23147 50759 23175
rect 50787 23147 50821 23175
rect 50849 23147 50883 23175
rect 50911 23147 50959 23175
rect 50649 23113 50959 23147
rect 50649 23085 50697 23113
rect 50725 23085 50759 23113
rect 50787 23085 50821 23113
rect 50849 23085 50883 23113
rect 50911 23085 50959 23113
rect 50649 23051 50959 23085
rect 50649 23023 50697 23051
rect 50725 23023 50759 23051
rect 50787 23023 50821 23051
rect 50849 23023 50883 23051
rect 50911 23023 50959 23051
rect 50649 22989 50959 23023
rect 50649 22961 50697 22989
rect 50725 22961 50759 22989
rect 50787 22961 50821 22989
rect 50849 22961 50883 22989
rect 50911 22961 50959 22989
rect 50649 14175 50959 22961
rect 61984 23175 62144 23192
rect 61984 23147 62019 23175
rect 62047 23147 62081 23175
rect 62109 23147 62144 23175
rect 61984 23113 62144 23147
rect 61984 23085 62019 23113
rect 62047 23085 62081 23113
rect 62109 23085 62144 23113
rect 61984 23051 62144 23085
rect 61984 23023 62019 23051
rect 62047 23023 62081 23051
rect 62109 23023 62144 23051
rect 61984 22989 62144 23023
rect 61984 22961 62019 22989
rect 62047 22961 62081 22989
rect 62109 22961 62144 22989
rect 61984 22944 62144 22961
rect 54304 20175 54464 20192
rect 54304 20147 54339 20175
rect 54367 20147 54401 20175
rect 54429 20147 54464 20175
rect 54304 20113 54464 20147
rect 54304 20085 54339 20113
rect 54367 20085 54401 20113
rect 54429 20085 54464 20113
rect 54304 20051 54464 20085
rect 54304 20023 54339 20051
rect 54367 20023 54401 20051
rect 54429 20023 54464 20051
rect 54304 19989 54464 20023
rect 54304 19961 54339 19989
rect 54367 19961 54401 19989
rect 54429 19961 54464 19989
rect 54304 19944 54464 19961
rect 64149 20175 64459 28961
rect 64149 20147 64197 20175
rect 64225 20147 64259 20175
rect 64287 20147 64321 20175
rect 64349 20147 64383 20175
rect 64411 20147 64459 20175
rect 64149 20113 64459 20147
rect 64149 20085 64197 20113
rect 64225 20085 64259 20113
rect 64287 20085 64321 20113
rect 64349 20085 64383 20113
rect 64411 20085 64459 20113
rect 64149 20051 64459 20085
rect 64149 20023 64197 20051
rect 64225 20023 64259 20051
rect 64287 20023 64321 20051
rect 64349 20023 64383 20051
rect 64411 20023 64459 20051
rect 64149 19989 64459 20023
rect 64149 19961 64197 19989
rect 64225 19961 64259 19989
rect 64287 19961 64321 19989
rect 64349 19961 64383 19989
rect 64411 19961 64459 19989
rect 50649 14147 50697 14175
rect 50725 14147 50759 14175
rect 50787 14147 50821 14175
rect 50849 14147 50883 14175
rect 50911 14147 50959 14175
rect 50649 14113 50959 14147
rect 50649 14085 50697 14113
rect 50725 14085 50759 14113
rect 50787 14085 50821 14113
rect 50849 14085 50883 14113
rect 50911 14085 50959 14113
rect 50649 14051 50959 14085
rect 50649 14023 50697 14051
rect 50725 14023 50759 14051
rect 50787 14023 50821 14051
rect 50849 14023 50883 14051
rect 50911 14023 50959 14051
rect 50649 13989 50959 14023
rect 50649 13961 50697 13989
rect 50725 13961 50759 13989
rect 50787 13961 50821 13989
rect 50849 13961 50883 13989
rect 50911 13961 50959 13989
rect 50649 5175 50959 13961
rect 61984 14175 62144 14192
rect 61984 14147 62019 14175
rect 62047 14147 62081 14175
rect 62109 14147 62144 14175
rect 61984 14113 62144 14147
rect 61984 14085 62019 14113
rect 62047 14085 62081 14113
rect 62109 14085 62144 14113
rect 61984 14051 62144 14085
rect 61984 14023 62019 14051
rect 62047 14023 62081 14051
rect 62109 14023 62144 14051
rect 61984 13989 62144 14023
rect 61984 13961 62019 13989
rect 62047 13961 62081 13989
rect 62109 13961 62144 13989
rect 61984 13944 62144 13961
rect 54304 11175 54464 11192
rect 54304 11147 54339 11175
rect 54367 11147 54401 11175
rect 54429 11147 54464 11175
rect 54304 11113 54464 11147
rect 54304 11085 54339 11113
rect 54367 11085 54401 11113
rect 54429 11085 54464 11113
rect 54304 11051 54464 11085
rect 54304 11023 54339 11051
rect 54367 11023 54401 11051
rect 54429 11023 54464 11051
rect 54304 10989 54464 11023
rect 54304 10961 54339 10989
rect 54367 10961 54401 10989
rect 54429 10961 54464 10989
rect 54304 10944 54464 10961
rect 64149 11175 64459 19961
rect 64149 11147 64197 11175
rect 64225 11147 64259 11175
rect 64287 11147 64321 11175
rect 64349 11147 64383 11175
rect 64411 11147 64459 11175
rect 64149 11113 64459 11147
rect 64149 11085 64197 11113
rect 64225 11085 64259 11113
rect 64287 11085 64321 11113
rect 64349 11085 64383 11113
rect 64411 11085 64459 11113
rect 64149 11051 64459 11085
rect 64149 11023 64197 11051
rect 64225 11023 64259 11051
rect 64287 11023 64321 11051
rect 64349 11023 64383 11051
rect 64411 11023 64459 11051
rect 64149 10989 64459 11023
rect 64149 10961 64197 10989
rect 64225 10961 64259 10989
rect 64287 10961 64321 10989
rect 64349 10961 64383 10989
rect 64411 10961 64459 10989
rect 50649 5147 50697 5175
rect 50725 5147 50759 5175
rect 50787 5147 50821 5175
rect 50849 5147 50883 5175
rect 50911 5147 50959 5175
rect 50649 5113 50959 5147
rect 50649 5085 50697 5113
rect 50725 5085 50759 5113
rect 50787 5085 50821 5113
rect 50849 5085 50883 5113
rect 50911 5085 50959 5113
rect 50649 5051 50959 5085
rect 50649 5023 50697 5051
rect 50725 5023 50759 5051
rect 50787 5023 50821 5051
rect 50849 5023 50883 5051
rect 50911 5023 50959 5051
rect 50649 4989 50959 5023
rect 50649 4961 50697 4989
rect 50725 4961 50759 4989
rect 50787 4961 50821 4989
rect 50849 4961 50883 4989
rect 50911 4961 50959 4989
rect 50649 -560 50959 4961
rect 61984 5175 62144 5192
rect 61984 5147 62019 5175
rect 62047 5147 62081 5175
rect 62109 5147 62144 5175
rect 61984 5113 62144 5147
rect 61984 5085 62019 5113
rect 62047 5085 62081 5113
rect 62109 5085 62144 5113
rect 61984 5051 62144 5085
rect 61984 5023 62019 5051
rect 62047 5023 62081 5051
rect 62109 5023 62144 5051
rect 61984 4989 62144 5023
rect 61984 4961 62019 4989
rect 62047 4961 62081 4989
rect 62109 4961 62144 4989
rect 61984 4944 62144 4961
rect 50649 -588 50697 -560
rect 50725 -588 50759 -560
rect 50787 -588 50821 -560
rect 50849 -588 50883 -560
rect 50911 -588 50959 -560
rect 50649 -622 50959 -588
rect 50649 -650 50697 -622
rect 50725 -650 50759 -622
rect 50787 -650 50821 -622
rect 50849 -650 50883 -622
rect 50911 -650 50959 -622
rect 50649 -684 50959 -650
rect 50649 -712 50697 -684
rect 50725 -712 50759 -684
rect 50787 -712 50821 -684
rect 50849 -712 50883 -684
rect 50911 -712 50959 -684
rect 50649 -746 50959 -712
rect 50649 -774 50697 -746
rect 50725 -774 50759 -746
rect 50787 -774 50821 -746
rect 50849 -774 50883 -746
rect 50911 -774 50959 -746
rect 50649 -822 50959 -774
rect 64149 2175 64459 10961
rect 64149 2147 64197 2175
rect 64225 2147 64259 2175
rect 64287 2147 64321 2175
rect 64349 2147 64383 2175
rect 64411 2147 64459 2175
rect 64149 2113 64459 2147
rect 64149 2085 64197 2113
rect 64225 2085 64259 2113
rect 64287 2085 64321 2113
rect 64349 2085 64383 2113
rect 64411 2085 64459 2113
rect 64149 2051 64459 2085
rect 64149 2023 64197 2051
rect 64225 2023 64259 2051
rect 64287 2023 64321 2051
rect 64349 2023 64383 2051
rect 64411 2023 64459 2051
rect 64149 1989 64459 2023
rect 64149 1961 64197 1989
rect 64225 1961 64259 1989
rect 64287 1961 64321 1989
rect 64349 1961 64383 1989
rect 64411 1961 64459 1989
rect 64149 -80 64459 1961
rect 64149 -108 64197 -80
rect 64225 -108 64259 -80
rect 64287 -108 64321 -80
rect 64349 -108 64383 -80
rect 64411 -108 64459 -80
rect 64149 -142 64459 -108
rect 64149 -170 64197 -142
rect 64225 -170 64259 -142
rect 64287 -170 64321 -142
rect 64349 -170 64383 -142
rect 64411 -170 64459 -142
rect 64149 -204 64459 -170
rect 64149 -232 64197 -204
rect 64225 -232 64259 -204
rect 64287 -232 64321 -204
rect 64349 -232 64383 -204
rect 64411 -232 64459 -204
rect 64149 -266 64459 -232
rect 64149 -294 64197 -266
rect 64225 -294 64259 -266
rect 64287 -294 64321 -266
rect 64349 -294 64383 -266
rect 64411 -294 64459 -266
rect 64149 -822 64459 -294
rect 66009 299086 66319 299134
rect 66009 299058 66057 299086
rect 66085 299058 66119 299086
rect 66147 299058 66181 299086
rect 66209 299058 66243 299086
rect 66271 299058 66319 299086
rect 66009 299024 66319 299058
rect 66009 298996 66057 299024
rect 66085 298996 66119 299024
rect 66147 298996 66181 299024
rect 66209 298996 66243 299024
rect 66271 298996 66319 299024
rect 66009 298962 66319 298996
rect 66009 298934 66057 298962
rect 66085 298934 66119 298962
rect 66147 298934 66181 298962
rect 66209 298934 66243 298962
rect 66271 298934 66319 298962
rect 66009 298900 66319 298934
rect 66009 298872 66057 298900
rect 66085 298872 66119 298900
rect 66147 298872 66181 298900
rect 66209 298872 66243 298900
rect 66271 298872 66319 298900
rect 66009 293175 66319 298872
rect 66009 293147 66057 293175
rect 66085 293147 66119 293175
rect 66147 293147 66181 293175
rect 66209 293147 66243 293175
rect 66271 293147 66319 293175
rect 66009 293113 66319 293147
rect 66009 293085 66057 293113
rect 66085 293085 66119 293113
rect 66147 293085 66181 293113
rect 66209 293085 66243 293113
rect 66271 293085 66319 293113
rect 66009 293051 66319 293085
rect 66009 293023 66057 293051
rect 66085 293023 66119 293051
rect 66147 293023 66181 293051
rect 66209 293023 66243 293051
rect 66271 293023 66319 293051
rect 66009 292989 66319 293023
rect 66009 292961 66057 292989
rect 66085 292961 66119 292989
rect 66147 292961 66181 292989
rect 66209 292961 66243 292989
rect 66271 292961 66319 292989
rect 66009 284175 66319 292961
rect 66009 284147 66057 284175
rect 66085 284147 66119 284175
rect 66147 284147 66181 284175
rect 66209 284147 66243 284175
rect 66271 284147 66319 284175
rect 66009 284113 66319 284147
rect 66009 284085 66057 284113
rect 66085 284085 66119 284113
rect 66147 284085 66181 284113
rect 66209 284085 66243 284113
rect 66271 284085 66319 284113
rect 66009 284051 66319 284085
rect 66009 284023 66057 284051
rect 66085 284023 66119 284051
rect 66147 284023 66181 284051
rect 66209 284023 66243 284051
rect 66271 284023 66319 284051
rect 66009 283989 66319 284023
rect 66009 283961 66057 283989
rect 66085 283961 66119 283989
rect 66147 283961 66181 283989
rect 66209 283961 66243 283989
rect 66271 283961 66319 283989
rect 66009 275175 66319 283961
rect 66009 275147 66057 275175
rect 66085 275147 66119 275175
rect 66147 275147 66181 275175
rect 66209 275147 66243 275175
rect 66271 275147 66319 275175
rect 66009 275113 66319 275147
rect 66009 275085 66057 275113
rect 66085 275085 66119 275113
rect 66147 275085 66181 275113
rect 66209 275085 66243 275113
rect 66271 275085 66319 275113
rect 66009 275051 66319 275085
rect 66009 275023 66057 275051
rect 66085 275023 66119 275051
rect 66147 275023 66181 275051
rect 66209 275023 66243 275051
rect 66271 275023 66319 275051
rect 66009 274989 66319 275023
rect 66009 274961 66057 274989
rect 66085 274961 66119 274989
rect 66147 274961 66181 274989
rect 66209 274961 66243 274989
rect 66271 274961 66319 274989
rect 66009 266175 66319 274961
rect 66009 266147 66057 266175
rect 66085 266147 66119 266175
rect 66147 266147 66181 266175
rect 66209 266147 66243 266175
rect 66271 266147 66319 266175
rect 66009 266113 66319 266147
rect 66009 266085 66057 266113
rect 66085 266085 66119 266113
rect 66147 266085 66181 266113
rect 66209 266085 66243 266113
rect 66271 266085 66319 266113
rect 66009 266051 66319 266085
rect 66009 266023 66057 266051
rect 66085 266023 66119 266051
rect 66147 266023 66181 266051
rect 66209 266023 66243 266051
rect 66271 266023 66319 266051
rect 66009 265989 66319 266023
rect 66009 265961 66057 265989
rect 66085 265961 66119 265989
rect 66147 265961 66181 265989
rect 66209 265961 66243 265989
rect 66271 265961 66319 265989
rect 66009 257175 66319 265961
rect 66009 257147 66057 257175
rect 66085 257147 66119 257175
rect 66147 257147 66181 257175
rect 66209 257147 66243 257175
rect 66271 257147 66319 257175
rect 66009 257113 66319 257147
rect 66009 257085 66057 257113
rect 66085 257085 66119 257113
rect 66147 257085 66181 257113
rect 66209 257085 66243 257113
rect 66271 257085 66319 257113
rect 66009 257051 66319 257085
rect 66009 257023 66057 257051
rect 66085 257023 66119 257051
rect 66147 257023 66181 257051
rect 66209 257023 66243 257051
rect 66271 257023 66319 257051
rect 66009 256989 66319 257023
rect 66009 256961 66057 256989
rect 66085 256961 66119 256989
rect 66147 256961 66181 256989
rect 66209 256961 66243 256989
rect 66271 256961 66319 256989
rect 66009 248175 66319 256961
rect 66009 248147 66057 248175
rect 66085 248147 66119 248175
rect 66147 248147 66181 248175
rect 66209 248147 66243 248175
rect 66271 248147 66319 248175
rect 66009 248113 66319 248147
rect 66009 248085 66057 248113
rect 66085 248085 66119 248113
rect 66147 248085 66181 248113
rect 66209 248085 66243 248113
rect 66271 248085 66319 248113
rect 66009 248051 66319 248085
rect 66009 248023 66057 248051
rect 66085 248023 66119 248051
rect 66147 248023 66181 248051
rect 66209 248023 66243 248051
rect 66271 248023 66319 248051
rect 66009 247989 66319 248023
rect 66009 247961 66057 247989
rect 66085 247961 66119 247989
rect 66147 247961 66181 247989
rect 66209 247961 66243 247989
rect 66271 247961 66319 247989
rect 66009 239175 66319 247961
rect 66009 239147 66057 239175
rect 66085 239147 66119 239175
rect 66147 239147 66181 239175
rect 66209 239147 66243 239175
rect 66271 239147 66319 239175
rect 66009 239113 66319 239147
rect 66009 239085 66057 239113
rect 66085 239085 66119 239113
rect 66147 239085 66181 239113
rect 66209 239085 66243 239113
rect 66271 239085 66319 239113
rect 66009 239051 66319 239085
rect 66009 239023 66057 239051
rect 66085 239023 66119 239051
rect 66147 239023 66181 239051
rect 66209 239023 66243 239051
rect 66271 239023 66319 239051
rect 66009 238989 66319 239023
rect 66009 238961 66057 238989
rect 66085 238961 66119 238989
rect 66147 238961 66181 238989
rect 66209 238961 66243 238989
rect 66271 238961 66319 238989
rect 66009 230175 66319 238961
rect 66009 230147 66057 230175
rect 66085 230147 66119 230175
rect 66147 230147 66181 230175
rect 66209 230147 66243 230175
rect 66271 230147 66319 230175
rect 66009 230113 66319 230147
rect 66009 230085 66057 230113
rect 66085 230085 66119 230113
rect 66147 230085 66181 230113
rect 66209 230085 66243 230113
rect 66271 230085 66319 230113
rect 66009 230051 66319 230085
rect 66009 230023 66057 230051
rect 66085 230023 66119 230051
rect 66147 230023 66181 230051
rect 66209 230023 66243 230051
rect 66271 230023 66319 230051
rect 66009 229989 66319 230023
rect 66009 229961 66057 229989
rect 66085 229961 66119 229989
rect 66147 229961 66181 229989
rect 66209 229961 66243 229989
rect 66271 229961 66319 229989
rect 66009 221175 66319 229961
rect 66009 221147 66057 221175
rect 66085 221147 66119 221175
rect 66147 221147 66181 221175
rect 66209 221147 66243 221175
rect 66271 221147 66319 221175
rect 66009 221113 66319 221147
rect 66009 221085 66057 221113
rect 66085 221085 66119 221113
rect 66147 221085 66181 221113
rect 66209 221085 66243 221113
rect 66271 221085 66319 221113
rect 66009 221051 66319 221085
rect 66009 221023 66057 221051
rect 66085 221023 66119 221051
rect 66147 221023 66181 221051
rect 66209 221023 66243 221051
rect 66271 221023 66319 221051
rect 66009 220989 66319 221023
rect 66009 220961 66057 220989
rect 66085 220961 66119 220989
rect 66147 220961 66181 220989
rect 66209 220961 66243 220989
rect 66271 220961 66319 220989
rect 66009 212175 66319 220961
rect 66009 212147 66057 212175
rect 66085 212147 66119 212175
rect 66147 212147 66181 212175
rect 66209 212147 66243 212175
rect 66271 212147 66319 212175
rect 66009 212113 66319 212147
rect 66009 212085 66057 212113
rect 66085 212085 66119 212113
rect 66147 212085 66181 212113
rect 66209 212085 66243 212113
rect 66271 212085 66319 212113
rect 66009 212051 66319 212085
rect 66009 212023 66057 212051
rect 66085 212023 66119 212051
rect 66147 212023 66181 212051
rect 66209 212023 66243 212051
rect 66271 212023 66319 212051
rect 66009 211989 66319 212023
rect 66009 211961 66057 211989
rect 66085 211961 66119 211989
rect 66147 211961 66181 211989
rect 66209 211961 66243 211989
rect 66271 211961 66319 211989
rect 66009 203175 66319 211961
rect 66009 203147 66057 203175
rect 66085 203147 66119 203175
rect 66147 203147 66181 203175
rect 66209 203147 66243 203175
rect 66271 203147 66319 203175
rect 66009 203113 66319 203147
rect 66009 203085 66057 203113
rect 66085 203085 66119 203113
rect 66147 203085 66181 203113
rect 66209 203085 66243 203113
rect 66271 203085 66319 203113
rect 66009 203051 66319 203085
rect 66009 203023 66057 203051
rect 66085 203023 66119 203051
rect 66147 203023 66181 203051
rect 66209 203023 66243 203051
rect 66271 203023 66319 203051
rect 66009 202989 66319 203023
rect 66009 202961 66057 202989
rect 66085 202961 66119 202989
rect 66147 202961 66181 202989
rect 66209 202961 66243 202989
rect 66271 202961 66319 202989
rect 66009 194175 66319 202961
rect 66009 194147 66057 194175
rect 66085 194147 66119 194175
rect 66147 194147 66181 194175
rect 66209 194147 66243 194175
rect 66271 194147 66319 194175
rect 66009 194113 66319 194147
rect 66009 194085 66057 194113
rect 66085 194085 66119 194113
rect 66147 194085 66181 194113
rect 66209 194085 66243 194113
rect 66271 194085 66319 194113
rect 66009 194051 66319 194085
rect 66009 194023 66057 194051
rect 66085 194023 66119 194051
rect 66147 194023 66181 194051
rect 66209 194023 66243 194051
rect 66271 194023 66319 194051
rect 66009 193989 66319 194023
rect 66009 193961 66057 193989
rect 66085 193961 66119 193989
rect 66147 193961 66181 193989
rect 66209 193961 66243 193989
rect 66271 193961 66319 193989
rect 66009 185175 66319 193961
rect 66009 185147 66057 185175
rect 66085 185147 66119 185175
rect 66147 185147 66181 185175
rect 66209 185147 66243 185175
rect 66271 185147 66319 185175
rect 66009 185113 66319 185147
rect 66009 185085 66057 185113
rect 66085 185085 66119 185113
rect 66147 185085 66181 185113
rect 66209 185085 66243 185113
rect 66271 185085 66319 185113
rect 66009 185051 66319 185085
rect 66009 185023 66057 185051
rect 66085 185023 66119 185051
rect 66147 185023 66181 185051
rect 66209 185023 66243 185051
rect 66271 185023 66319 185051
rect 66009 184989 66319 185023
rect 66009 184961 66057 184989
rect 66085 184961 66119 184989
rect 66147 184961 66181 184989
rect 66209 184961 66243 184989
rect 66271 184961 66319 184989
rect 66009 176175 66319 184961
rect 66009 176147 66057 176175
rect 66085 176147 66119 176175
rect 66147 176147 66181 176175
rect 66209 176147 66243 176175
rect 66271 176147 66319 176175
rect 66009 176113 66319 176147
rect 66009 176085 66057 176113
rect 66085 176085 66119 176113
rect 66147 176085 66181 176113
rect 66209 176085 66243 176113
rect 66271 176085 66319 176113
rect 66009 176051 66319 176085
rect 66009 176023 66057 176051
rect 66085 176023 66119 176051
rect 66147 176023 66181 176051
rect 66209 176023 66243 176051
rect 66271 176023 66319 176051
rect 66009 175989 66319 176023
rect 66009 175961 66057 175989
rect 66085 175961 66119 175989
rect 66147 175961 66181 175989
rect 66209 175961 66243 175989
rect 66271 175961 66319 175989
rect 66009 167175 66319 175961
rect 79509 298606 79819 299134
rect 79509 298578 79557 298606
rect 79585 298578 79619 298606
rect 79647 298578 79681 298606
rect 79709 298578 79743 298606
rect 79771 298578 79819 298606
rect 79509 298544 79819 298578
rect 79509 298516 79557 298544
rect 79585 298516 79619 298544
rect 79647 298516 79681 298544
rect 79709 298516 79743 298544
rect 79771 298516 79819 298544
rect 79509 298482 79819 298516
rect 79509 298454 79557 298482
rect 79585 298454 79619 298482
rect 79647 298454 79681 298482
rect 79709 298454 79743 298482
rect 79771 298454 79819 298482
rect 79509 298420 79819 298454
rect 79509 298392 79557 298420
rect 79585 298392 79619 298420
rect 79647 298392 79681 298420
rect 79709 298392 79743 298420
rect 79771 298392 79819 298420
rect 79509 290175 79819 298392
rect 79509 290147 79557 290175
rect 79585 290147 79619 290175
rect 79647 290147 79681 290175
rect 79709 290147 79743 290175
rect 79771 290147 79819 290175
rect 79509 290113 79819 290147
rect 79509 290085 79557 290113
rect 79585 290085 79619 290113
rect 79647 290085 79681 290113
rect 79709 290085 79743 290113
rect 79771 290085 79819 290113
rect 79509 290051 79819 290085
rect 79509 290023 79557 290051
rect 79585 290023 79619 290051
rect 79647 290023 79681 290051
rect 79709 290023 79743 290051
rect 79771 290023 79819 290051
rect 79509 289989 79819 290023
rect 79509 289961 79557 289989
rect 79585 289961 79619 289989
rect 79647 289961 79681 289989
rect 79709 289961 79743 289989
rect 79771 289961 79819 289989
rect 79509 281175 79819 289961
rect 79509 281147 79557 281175
rect 79585 281147 79619 281175
rect 79647 281147 79681 281175
rect 79709 281147 79743 281175
rect 79771 281147 79819 281175
rect 79509 281113 79819 281147
rect 79509 281085 79557 281113
rect 79585 281085 79619 281113
rect 79647 281085 79681 281113
rect 79709 281085 79743 281113
rect 79771 281085 79819 281113
rect 79509 281051 79819 281085
rect 79509 281023 79557 281051
rect 79585 281023 79619 281051
rect 79647 281023 79681 281051
rect 79709 281023 79743 281051
rect 79771 281023 79819 281051
rect 79509 280989 79819 281023
rect 79509 280961 79557 280989
rect 79585 280961 79619 280989
rect 79647 280961 79681 280989
rect 79709 280961 79743 280989
rect 79771 280961 79819 280989
rect 79509 272175 79819 280961
rect 79509 272147 79557 272175
rect 79585 272147 79619 272175
rect 79647 272147 79681 272175
rect 79709 272147 79743 272175
rect 79771 272147 79819 272175
rect 79509 272113 79819 272147
rect 79509 272085 79557 272113
rect 79585 272085 79619 272113
rect 79647 272085 79681 272113
rect 79709 272085 79743 272113
rect 79771 272085 79819 272113
rect 79509 272051 79819 272085
rect 79509 272023 79557 272051
rect 79585 272023 79619 272051
rect 79647 272023 79681 272051
rect 79709 272023 79743 272051
rect 79771 272023 79819 272051
rect 79509 271989 79819 272023
rect 79509 271961 79557 271989
rect 79585 271961 79619 271989
rect 79647 271961 79681 271989
rect 79709 271961 79743 271989
rect 79771 271961 79819 271989
rect 79509 263175 79819 271961
rect 79509 263147 79557 263175
rect 79585 263147 79619 263175
rect 79647 263147 79681 263175
rect 79709 263147 79743 263175
rect 79771 263147 79819 263175
rect 79509 263113 79819 263147
rect 79509 263085 79557 263113
rect 79585 263085 79619 263113
rect 79647 263085 79681 263113
rect 79709 263085 79743 263113
rect 79771 263085 79819 263113
rect 79509 263051 79819 263085
rect 79509 263023 79557 263051
rect 79585 263023 79619 263051
rect 79647 263023 79681 263051
rect 79709 263023 79743 263051
rect 79771 263023 79819 263051
rect 79509 262989 79819 263023
rect 79509 262961 79557 262989
rect 79585 262961 79619 262989
rect 79647 262961 79681 262989
rect 79709 262961 79743 262989
rect 79771 262961 79819 262989
rect 79509 254175 79819 262961
rect 79509 254147 79557 254175
rect 79585 254147 79619 254175
rect 79647 254147 79681 254175
rect 79709 254147 79743 254175
rect 79771 254147 79819 254175
rect 79509 254113 79819 254147
rect 79509 254085 79557 254113
rect 79585 254085 79619 254113
rect 79647 254085 79681 254113
rect 79709 254085 79743 254113
rect 79771 254085 79819 254113
rect 79509 254051 79819 254085
rect 79509 254023 79557 254051
rect 79585 254023 79619 254051
rect 79647 254023 79681 254051
rect 79709 254023 79743 254051
rect 79771 254023 79819 254051
rect 79509 253989 79819 254023
rect 79509 253961 79557 253989
rect 79585 253961 79619 253989
rect 79647 253961 79681 253989
rect 79709 253961 79743 253989
rect 79771 253961 79819 253989
rect 79509 245175 79819 253961
rect 79509 245147 79557 245175
rect 79585 245147 79619 245175
rect 79647 245147 79681 245175
rect 79709 245147 79743 245175
rect 79771 245147 79819 245175
rect 79509 245113 79819 245147
rect 79509 245085 79557 245113
rect 79585 245085 79619 245113
rect 79647 245085 79681 245113
rect 79709 245085 79743 245113
rect 79771 245085 79819 245113
rect 79509 245051 79819 245085
rect 79509 245023 79557 245051
rect 79585 245023 79619 245051
rect 79647 245023 79681 245051
rect 79709 245023 79743 245051
rect 79771 245023 79819 245051
rect 79509 244989 79819 245023
rect 79509 244961 79557 244989
rect 79585 244961 79619 244989
rect 79647 244961 79681 244989
rect 79709 244961 79743 244989
rect 79771 244961 79819 244989
rect 79509 236175 79819 244961
rect 79509 236147 79557 236175
rect 79585 236147 79619 236175
rect 79647 236147 79681 236175
rect 79709 236147 79743 236175
rect 79771 236147 79819 236175
rect 79509 236113 79819 236147
rect 79509 236085 79557 236113
rect 79585 236085 79619 236113
rect 79647 236085 79681 236113
rect 79709 236085 79743 236113
rect 79771 236085 79819 236113
rect 79509 236051 79819 236085
rect 79509 236023 79557 236051
rect 79585 236023 79619 236051
rect 79647 236023 79681 236051
rect 79709 236023 79743 236051
rect 79771 236023 79819 236051
rect 79509 235989 79819 236023
rect 79509 235961 79557 235989
rect 79585 235961 79619 235989
rect 79647 235961 79681 235989
rect 79709 235961 79743 235989
rect 79771 235961 79819 235989
rect 79509 227175 79819 235961
rect 79509 227147 79557 227175
rect 79585 227147 79619 227175
rect 79647 227147 79681 227175
rect 79709 227147 79743 227175
rect 79771 227147 79819 227175
rect 79509 227113 79819 227147
rect 79509 227085 79557 227113
rect 79585 227085 79619 227113
rect 79647 227085 79681 227113
rect 79709 227085 79743 227113
rect 79771 227085 79819 227113
rect 79509 227051 79819 227085
rect 79509 227023 79557 227051
rect 79585 227023 79619 227051
rect 79647 227023 79681 227051
rect 79709 227023 79743 227051
rect 79771 227023 79819 227051
rect 79509 226989 79819 227023
rect 79509 226961 79557 226989
rect 79585 226961 79619 226989
rect 79647 226961 79681 226989
rect 79709 226961 79743 226989
rect 79771 226961 79819 226989
rect 79509 218175 79819 226961
rect 79509 218147 79557 218175
rect 79585 218147 79619 218175
rect 79647 218147 79681 218175
rect 79709 218147 79743 218175
rect 79771 218147 79819 218175
rect 79509 218113 79819 218147
rect 79509 218085 79557 218113
rect 79585 218085 79619 218113
rect 79647 218085 79681 218113
rect 79709 218085 79743 218113
rect 79771 218085 79819 218113
rect 79509 218051 79819 218085
rect 79509 218023 79557 218051
rect 79585 218023 79619 218051
rect 79647 218023 79681 218051
rect 79709 218023 79743 218051
rect 79771 218023 79819 218051
rect 79509 217989 79819 218023
rect 79509 217961 79557 217989
rect 79585 217961 79619 217989
rect 79647 217961 79681 217989
rect 79709 217961 79743 217989
rect 79771 217961 79819 217989
rect 79509 209175 79819 217961
rect 79509 209147 79557 209175
rect 79585 209147 79619 209175
rect 79647 209147 79681 209175
rect 79709 209147 79743 209175
rect 79771 209147 79819 209175
rect 79509 209113 79819 209147
rect 79509 209085 79557 209113
rect 79585 209085 79619 209113
rect 79647 209085 79681 209113
rect 79709 209085 79743 209113
rect 79771 209085 79819 209113
rect 79509 209051 79819 209085
rect 79509 209023 79557 209051
rect 79585 209023 79619 209051
rect 79647 209023 79681 209051
rect 79709 209023 79743 209051
rect 79771 209023 79819 209051
rect 79509 208989 79819 209023
rect 79509 208961 79557 208989
rect 79585 208961 79619 208989
rect 79647 208961 79681 208989
rect 79709 208961 79743 208989
rect 79771 208961 79819 208989
rect 79509 200175 79819 208961
rect 79509 200147 79557 200175
rect 79585 200147 79619 200175
rect 79647 200147 79681 200175
rect 79709 200147 79743 200175
rect 79771 200147 79819 200175
rect 79509 200113 79819 200147
rect 79509 200085 79557 200113
rect 79585 200085 79619 200113
rect 79647 200085 79681 200113
rect 79709 200085 79743 200113
rect 79771 200085 79819 200113
rect 79509 200051 79819 200085
rect 79509 200023 79557 200051
rect 79585 200023 79619 200051
rect 79647 200023 79681 200051
rect 79709 200023 79743 200051
rect 79771 200023 79819 200051
rect 79509 199989 79819 200023
rect 79509 199961 79557 199989
rect 79585 199961 79619 199989
rect 79647 199961 79681 199989
rect 79709 199961 79743 199989
rect 79771 199961 79819 199989
rect 79509 191175 79819 199961
rect 79509 191147 79557 191175
rect 79585 191147 79619 191175
rect 79647 191147 79681 191175
rect 79709 191147 79743 191175
rect 79771 191147 79819 191175
rect 79509 191113 79819 191147
rect 79509 191085 79557 191113
rect 79585 191085 79619 191113
rect 79647 191085 79681 191113
rect 79709 191085 79743 191113
rect 79771 191085 79819 191113
rect 79509 191051 79819 191085
rect 79509 191023 79557 191051
rect 79585 191023 79619 191051
rect 79647 191023 79681 191051
rect 79709 191023 79743 191051
rect 79771 191023 79819 191051
rect 79509 190989 79819 191023
rect 79509 190961 79557 190989
rect 79585 190961 79619 190989
rect 79647 190961 79681 190989
rect 79709 190961 79743 190989
rect 79771 190961 79819 190989
rect 79509 182175 79819 190961
rect 79509 182147 79557 182175
rect 79585 182147 79619 182175
rect 79647 182147 79681 182175
rect 79709 182147 79743 182175
rect 79771 182147 79819 182175
rect 79509 182113 79819 182147
rect 79509 182085 79557 182113
rect 79585 182085 79619 182113
rect 79647 182085 79681 182113
rect 79709 182085 79743 182113
rect 79771 182085 79819 182113
rect 79509 182051 79819 182085
rect 79509 182023 79557 182051
rect 79585 182023 79619 182051
rect 79647 182023 79681 182051
rect 79709 182023 79743 182051
rect 79771 182023 79819 182051
rect 79509 181989 79819 182023
rect 79509 181961 79557 181989
rect 79585 181961 79619 181989
rect 79647 181961 79681 181989
rect 79709 181961 79743 181989
rect 79771 181961 79819 181989
rect 69664 173175 69824 173192
rect 69664 173147 69699 173175
rect 69727 173147 69761 173175
rect 69789 173147 69824 173175
rect 69664 173113 69824 173147
rect 69664 173085 69699 173113
rect 69727 173085 69761 173113
rect 69789 173085 69824 173113
rect 69664 173051 69824 173085
rect 69664 173023 69699 173051
rect 69727 173023 69761 173051
rect 69789 173023 69824 173051
rect 69664 172989 69824 173023
rect 69664 172961 69699 172989
rect 69727 172961 69761 172989
rect 69789 172961 69824 172989
rect 69664 172944 69824 172961
rect 79509 173175 79819 181961
rect 79509 173147 79557 173175
rect 79585 173147 79619 173175
rect 79647 173147 79681 173175
rect 79709 173147 79743 173175
rect 79771 173147 79819 173175
rect 79509 173113 79819 173147
rect 79509 173085 79557 173113
rect 79585 173085 79619 173113
rect 79647 173085 79681 173113
rect 79709 173085 79743 173113
rect 79771 173085 79819 173113
rect 79509 173051 79819 173085
rect 79509 173023 79557 173051
rect 79585 173023 79619 173051
rect 79647 173023 79681 173051
rect 79709 173023 79743 173051
rect 79771 173023 79819 173051
rect 79509 172989 79819 173023
rect 79509 172961 79557 172989
rect 79585 172961 79619 172989
rect 79647 172961 79681 172989
rect 79709 172961 79743 172989
rect 79771 172961 79819 172989
rect 66009 167147 66057 167175
rect 66085 167147 66119 167175
rect 66147 167147 66181 167175
rect 66209 167147 66243 167175
rect 66271 167147 66319 167175
rect 66009 167113 66319 167147
rect 66009 167085 66057 167113
rect 66085 167085 66119 167113
rect 66147 167085 66181 167113
rect 66209 167085 66243 167113
rect 66271 167085 66319 167113
rect 66009 167051 66319 167085
rect 66009 167023 66057 167051
rect 66085 167023 66119 167051
rect 66147 167023 66181 167051
rect 66209 167023 66243 167051
rect 66271 167023 66319 167051
rect 66009 166989 66319 167023
rect 66009 166961 66057 166989
rect 66085 166961 66119 166989
rect 66147 166961 66181 166989
rect 66209 166961 66243 166989
rect 66271 166961 66319 166989
rect 66009 158175 66319 166961
rect 77344 167175 77504 167192
rect 77344 167147 77379 167175
rect 77407 167147 77441 167175
rect 77469 167147 77504 167175
rect 77344 167113 77504 167147
rect 77344 167085 77379 167113
rect 77407 167085 77441 167113
rect 77469 167085 77504 167113
rect 77344 167051 77504 167085
rect 77344 167023 77379 167051
rect 77407 167023 77441 167051
rect 77469 167023 77504 167051
rect 77344 166989 77504 167023
rect 77344 166961 77379 166989
rect 77407 166961 77441 166989
rect 77469 166961 77504 166989
rect 77344 166944 77504 166961
rect 69664 164175 69824 164192
rect 69664 164147 69699 164175
rect 69727 164147 69761 164175
rect 69789 164147 69824 164175
rect 69664 164113 69824 164147
rect 69664 164085 69699 164113
rect 69727 164085 69761 164113
rect 69789 164085 69824 164113
rect 69664 164051 69824 164085
rect 69664 164023 69699 164051
rect 69727 164023 69761 164051
rect 69789 164023 69824 164051
rect 69664 163989 69824 164023
rect 69664 163961 69699 163989
rect 69727 163961 69761 163989
rect 69789 163961 69824 163989
rect 69664 163944 69824 163961
rect 79509 164175 79819 172961
rect 79509 164147 79557 164175
rect 79585 164147 79619 164175
rect 79647 164147 79681 164175
rect 79709 164147 79743 164175
rect 79771 164147 79819 164175
rect 79509 164113 79819 164147
rect 79509 164085 79557 164113
rect 79585 164085 79619 164113
rect 79647 164085 79681 164113
rect 79709 164085 79743 164113
rect 79771 164085 79819 164113
rect 79509 164051 79819 164085
rect 79509 164023 79557 164051
rect 79585 164023 79619 164051
rect 79647 164023 79681 164051
rect 79709 164023 79743 164051
rect 79771 164023 79819 164051
rect 79509 163989 79819 164023
rect 79509 163961 79557 163989
rect 79585 163961 79619 163989
rect 79647 163961 79681 163989
rect 79709 163961 79743 163989
rect 79771 163961 79819 163989
rect 66009 158147 66057 158175
rect 66085 158147 66119 158175
rect 66147 158147 66181 158175
rect 66209 158147 66243 158175
rect 66271 158147 66319 158175
rect 66009 158113 66319 158147
rect 66009 158085 66057 158113
rect 66085 158085 66119 158113
rect 66147 158085 66181 158113
rect 66209 158085 66243 158113
rect 66271 158085 66319 158113
rect 66009 158051 66319 158085
rect 66009 158023 66057 158051
rect 66085 158023 66119 158051
rect 66147 158023 66181 158051
rect 66209 158023 66243 158051
rect 66271 158023 66319 158051
rect 66009 157989 66319 158023
rect 66009 157961 66057 157989
rect 66085 157961 66119 157989
rect 66147 157961 66181 157989
rect 66209 157961 66243 157989
rect 66271 157961 66319 157989
rect 66009 149175 66319 157961
rect 77344 158175 77504 158192
rect 77344 158147 77379 158175
rect 77407 158147 77441 158175
rect 77469 158147 77504 158175
rect 77344 158113 77504 158147
rect 77344 158085 77379 158113
rect 77407 158085 77441 158113
rect 77469 158085 77504 158113
rect 77344 158051 77504 158085
rect 77344 158023 77379 158051
rect 77407 158023 77441 158051
rect 77469 158023 77504 158051
rect 77344 157989 77504 158023
rect 77344 157961 77379 157989
rect 77407 157961 77441 157989
rect 77469 157961 77504 157989
rect 77344 157944 77504 157961
rect 69664 155175 69824 155192
rect 69664 155147 69699 155175
rect 69727 155147 69761 155175
rect 69789 155147 69824 155175
rect 69664 155113 69824 155147
rect 69664 155085 69699 155113
rect 69727 155085 69761 155113
rect 69789 155085 69824 155113
rect 69664 155051 69824 155085
rect 69664 155023 69699 155051
rect 69727 155023 69761 155051
rect 69789 155023 69824 155051
rect 69664 154989 69824 155023
rect 69664 154961 69699 154989
rect 69727 154961 69761 154989
rect 69789 154961 69824 154989
rect 69664 154944 69824 154961
rect 79509 155175 79819 163961
rect 79509 155147 79557 155175
rect 79585 155147 79619 155175
rect 79647 155147 79681 155175
rect 79709 155147 79743 155175
rect 79771 155147 79819 155175
rect 79509 155113 79819 155147
rect 79509 155085 79557 155113
rect 79585 155085 79619 155113
rect 79647 155085 79681 155113
rect 79709 155085 79743 155113
rect 79771 155085 79819 155113
rect 79509 155051 79819 155085
rect 79509 155023 79557 155051
rect 79585 155023 79619 155051
rect 79647 155023 79681 155051
rect 79709 155023 79743 155051
rect 79771 155023 79819 155051
rect 79509 154989 79819 155023
rect 79509 154961 79557 154989
rect 79585 154961 79619 154989
rect 79647 154961 79681 154989
rect 79709 154961 79743 154989
rect 79771 154961 79819 154989
rect 66009 149147 66057 149175
rect 66085 149147 66119 149175
rect 66147 149147 66181 149175
rect 66209 149147 66243 149175
rect 66271 149147 66319 149175
rect 66009 149113 66319 149147
rect 66009 149085 66057 149113
rect 66085 149085 66119 149113
rect 66147 149085 66181 149113
rect 66209 149085 66243 149113
rect 66271 149085 66319 149113
rect 66009 149051 66319 149085
rect 66009 149023 66057 149051
rect 66085 149023 66119 149051
rect 66147 149023 66181 149051
rect 66209 149023 66243 149051
rect 66271 149023 66319 149051
rect 66009 148989 66319 149023
rect 66009 148961 66057 148989
rect 66085 148961 66119 148989
rect 66147 148961 66181 148989
rect 66209 148961 66243 148989
rect 66271 148961 66319 148989
rect 66009 140175 66319 148961
rect 77344 149175 77504 149192
rect 77344 149147 77379 149175
rect 77407 149147 77441 149175
rect 77469 149147 77504 149175
rect 77344 149113 77504 149147
rect 77344 149085 77379 149113
rect 77407 149085 77441 149113
rect 77469 149085 77504 149113
rect 77344 149051 77504 149085
rect 77344 149023 77379 149051
rect 77407 149023 77441 149051
rect 77469 149023 77504 149051
rect 77344 148989 77504 149023
rect 77344 148961 77379 148989
rect 77407 148961 77441 148989
rect 77469 148961 77504 148989
rect 77344 148944 77504 148961
rect 69664 146175 69824 146192
rect 69664 146147 69699 146175
rect 69727 146147 69761 146175
rect 69789 146147 69824 146175
rect 69664 146113 69824 146147
rect 69664 146085 69699 146113
rect 69727 146085 69761 146113
rect 69789 146085 69824 146113
rect 69664 146051 69824 146085
rect 69664 146023 69699 146051
rect 69727 146023 69761 146051
rect 69789 146023 69824 146051
rect 69664 145989 69824 146023
rect 69664 145961 69699 145989
rect 69727 145961 69761 145989
rect 69789 145961 69824 145989
rect 69664 145944 69824 145961
rect 79509 146175 79819 154961
rect 79509 146147 79557 146175
rect 79585 146147 79619 146175
rect 79647 146147 79681 146175
rect 79709 146147 79743 146175
rect 79771 146147 79819 146175
rect 79509 146113 79819 146147
rect 79509 146085 79557 146113
rect 79585 146085 79619 146113
rect 79647 146085 79681 146113
rect 79709 146085 79743 146113
rect 79771 146085 79819 146113
rect 79509 146051 79819 146085
rect 79509 146023 79557 146051
rect 79585 146023 79619 146051
rect 79647 146023 79681 146051
rect 79709 146023 79743 146051
rect 79771 146023 79819 146051
rect 79509 145989 79819 146023
rect 79509 145961 79557 145989
rect 79585 145961 79619 145989
rect 79647 145961 79681 145989
rect 79709 145961 79743 145989
rect 79771 145961 79819 145989
rect 66009 140147 66057 140175
rect 66085 140147 66119 140175
rect 66147 140147 66181 140175
rect 66209 140147 66243 140175
rect 66271 140147 66319 140175
rect 66009 140113 66319 140147
rect 66009 140085 66057 140113
rect 66085 140085 66119 140113
rect 66147 140085 66181 140113
rect 66209 140085 66243 140113
rect 66271 140085 66319 140113
rect 66009 140051 66319 140085
rect 66009 140023 66057 140051
rect 66085 140023 66119 140051
rect 66147 140023 66181 140051
rect 66209 140023 66243 140051
rect 66271 140023 66319 140051
rect 66009 139989 66319 140023
rect 66009 139961 66057 139989
rect 66085 139961 66119 139989
rect 66147 139961 66181 139989
rect 66209 139961 66243 139989
rect 66271 139961 66319 139989
rect 66009 131175 66319 139961
rect 77344 140175 77504 140192
rect 77344 140147 77379 140175
rect 77407 140147 77441 140175
rect 77469 140147 77504 140175
rect 77344 140113 77504 140147
rect 77344 140085 77379 140113
rect 77407 140085 77441 140113
rect 77469 140085 77504 140113
rect 77344 140051 77504 140085
rect 77344 140023 77379 140051
rect 77407 140023 77441 140051
rect 77469 140023 77504 140051
rect 77344 139989 77504 140023
rect 77344 139961 77379 139989
rect 77407 139961 77441 139989
rect 77469 139961 77504 139989
rect 77344 139944 77504 139961
rect 69664 137175 69824 137192
rect 69664 137147 69699 137175
rect 69727 137147 69761 137175
rect 69789 137147 69824 137175
rect 69664 137113 69824 137147
rect 69664 137085 69699 137113
rect 69727 137085 69761 137113
rect 69789 137085 69824 137113
rect 69664 137051 69824 137085
rect 69664 137023 69699 137051
rect 69727 137023 69761 137051
rect 69789 137023 69824 137051
rect 69664 136989 69824 137023
rect 69664 136961 69699 136989
rect 69727 136961 69761 136989
rect 69789 136961 69824 136989
rect 69664 136944 69824 136961
rect 79509 137175 79819 145961
rect 79509 137147 79557 137175
rect 79585 137147 79619 137175
rect 79647 137147 79681 137175
rect 79709 137147 79743 137175
rect 79771 137147 79819 137175
rect 79509 137113 79819 137147
rect 79509 137085 79557 137113
rect 79585 137085 79619 137113
rect 79647 137085 79681 137113
rect 79709 137085 79743 137113
rect 79771 137085 79819 137113
rect 79509 137051 79819 137085
rect 79509 137023 79557 137051
rect 79585 137023 79619 137051
rect 79647 137023 79681 137051
rect 79709 137023 79743 137051
rect 79771 137023 79819 137051
rect 79509 136989 79819 137023
rect 79509 136961 79557 136989
rect 79585 136961 79619 136989
rect 79647 136961 79681 136989
rect 79709 136961 79743 136989
rect 79771 136961 79819 136989
rect 66009 131147 66057 131175
rect 66085 131147 66119 131175
rect 66147 131147 66181 131175
rect 66209 131147 66243 131175
rect 66271 131147 66319 131175
rect 66009 131113 66319 131147
rect 66009 131085 66057 131113
rect 66085 131085 66119 131113
rect 66147 131085 66181 131113
rect 66209 131085 66243 131113
rect 66271 131085 66319 131113
rect 66009 131051 66319 131085
rect 66009 131023 66057 131051
rect 66085 131023 66119 131051
rect 66147 131023 66181 131051
rect 66209 131023 66243 131051
rect 66271 131023 66319 131051
rect 66009 130989 66319 131023
rect 66009 130961 66057 130989
rect 66085 130961 66119 130989
rect 66147 130961 66181 130989
rect 66209 130961 66243 130989
rect 66271 130961 66319 130989
rect 66009 122175 66319 130961
rect 77344 131175 77504 131192
rect 77344 131147 77379 131175
rect 77407 131147 77441 131175
rect 77469 131147 77504 131175
rect 77344 131113 77504 131147
rect 77344 131085 77379 131113
rect 77407 131085 77441 131113
rect 77469 131085 77504 131113
rect 77344 131051 77504 131085
rect 77344 131023 77379 131051
rect 77407 131023 77441 131051
rect 77469 131023 77504 131051
rect 77344 130989 77504 131023
rect 77344 130961 77379 130989
rect 77407 130961 77441 130989
rect 77469 130961 77504 130989
rect 77344 130944 77504 130961
rect 69664 128175 69824 128192
rect 69664 128147 69699 128175
rect 69727 128147 69761 128175
rect 69789 128147 69824 128175
rect 69664 128113 69824 128147
rect 69664 128085 69699 128113
rect 69727 128085 69761 128113
rect 69789 128085 69824 128113
rect 69664 128051 69824 128085
rect 69664 128023 69699 128051
rect 69727 128023 69761 128051
rect 69789 128023 69824 128051
rect 69664 127989 69824 128023
rect 69664 127961 69699 127989
rect 69727 127961 69761 127989
rect 69789 127961 69824 127989
rect 69664 127944 69824 127961
rect 79509 128175 79819 136961
rect 79509 128147 79557 128175
rect 79585 128147 79619 128175
rect 79647 128147 79681 128175
rect 79709 128147 79743 128175
rect 79771 128147 79819 128175
rect 79509 128113 79819 128147
rect 79509 128085 79557 128113
rect 79585 128085 79619 128113
rect 79647 128085 79681 128113
rect 79709 128085 79743 128113
rect 79771 128085 79819 128113
rect 79509 128051 79819 128085
rect 79509 128023 79557 128051
rect 79585 128023 79619 128051
rect 79647 128023 79681 128051
rect 79709 128023 79743 128051
rect 79771 128023 79819 128051
rect 79509 127989 79819 128023
rect 79509 127961 79557 127989
rect 79585 127961 79619 127989
rect 79647 127961 79681 127989
rect 79709 127961 79743 127989
rect 79771 127961 79819 127989
rect 66009 122147 66057 122175
rect 66085 122147 66119 122175
rect 66147 122147 66181 122175
rect 66209 122147 66243 122175
rect 66271 122147 66319 122175
rect 66009 122113 66319 122147
rect 66009 122085 66057 122113
rect 66085 122085 66119 122113
rect 66147 122085 66181 122113
rect 66209 122085 66243 122113
rect 66271 122085 66319 122113
rect 66009 122051 66319 122085
rect 66009 122023 66057 122051
rect 66085 122023 66119 122051
rect 66147 122023 66181 122051
rect 66209 122023 66243 122051
rect 66271 122023 66319 122051
rect 66009 121989 66319 122023
rect 66009 121961 66057 121989
rect 66085 121961 66119 121989
rect 66147 121961 66181 121989
rect 66209 121961 66243 121989
rect 66271 121961 66319 121989
rect 66009 113175 66319 121961
rect 77344 122175 77504 122192
rect 77344 122147 77379 122175
rect 77407 122147 77441 122175
rect 77469 122147 77504 122175
rect 77344 122113 77504 122147
rect 77344 122085 77379 122113
rect 77407 122085 77441 122113
rect 77469 122085 77504 122113
rect 77344 122051 77504 122085
rect 77344 122023 77379 122051
rect 77407 122023 77441 122051
rect 77469 122023 77504 122051
rect 77344 121989 77504 122023
rect 77344 121961 77379 121989
rect 77407 121961 77441 121989
rect 77469 121961 77504 121989
rect 77344 121944 77504 121961
rect 69664 119175 69824 119192
rect 69664 119147 69699 119175
rect 69727 119147 69761 119175
rect 69789 119147 69824 119175
rect 69664 119113 69824 119147
rect 69664 119085 69699 119113
rect 69727 119085 69761 119113
rect 69789 119085 69824 119113
rect 69664 119051 69824 119085
rect 69664 119023 69699 119051
rect 69727 119023 69761 119051
rect 69789 119023 69824 119051
rect 69664 118989 69824 119023
rect 69664 118961 69699 118989
rect 69727 118961 69761 118989
rect 69789 118961 69824 118989
rect 69664 118944 69824 118961
rect 79509 119175 79819 127961
rect 79509 119147 79557 119175
rect 79585 119147 79619 119175
rect 79647 119147 79681 119175
rect 79709 119147 79743 119175
rect 79771 119147 79819 119175
rect 79509 119113 79819 119147
rect 79509 119085 79557 119113
rect 79585 119085 79619 119113
rect 79647 119085 79681 119113
rect 79709 119085 79743 119113
rect 79771 119085 79819 119113
rect 79509 119051 79819 119085
rect 79509 119023 79557 119051
rect 79585 119023 79619 119051
rect 79647 119023 79681 119051
rect 79709 119023 79743 119051
rect 79771 119023 79819 119051
rect 79509 118989 79819 119023
rect 79509 118961 79557 118989
rect 79585 118961 79619 118989
rect 79647 118961 79681 118989
rect 79709 118961 79743 118989
rect 79771 118961 79819 118989
rect 66009 113147 66057 113175
rect 66085 113147 66119 113175
rect 66147 113147 66181 113175
rect 66209 113147 66243 113175
rect 66271 113147 66319 113175
rect 66009 113113 66319 113147
rect 66009 113085 66057 113113
rect 66085 113085 66119 113113
rect 66147 113085 66181 113113
rect 66209 113085 66243 113113
rect 66271 113085 66319 113113
rect 66009 113051 66319 113085
rect 66009 113023 66057 113051
rect 66085 113023 66119 113051
rect 66147 113023 66181 113051
rect 66209 113023 66243 113051
rect 66271 113023 66319 113051
rect 66009 112989 66319 113023
rect 66009 112961 66057 112989
rect 66085 112961 66119 112989
rect 66147 112961 66181 112989
rect 66209 112961 66243 112989
rect 66271 112961 66319 112989
rect 66009 104175 66319 112961
rect 77344 113175 77504 113192
rect 77344 113147 77379 113175
rect 77407 113147 77441 113175
rect 77469 113147 77504 113175
rect 77344 113113 77504 113147
rect 77344 113085 77379 113113
rect 77407 113085 77441 113113
rect 77469 113085 77504 113113
rect 77344 113051 77504 113085
rect 77344 113023 77379 113051
rect 77407 113023 77441 113051
rect 77469 113023 77504 113051
rect 77344 112989 77504 113023
rect 77344 112961 77379 112989
rect 77407 112961 77441 112989
rect 77469 112961 77504 112989
rect 77344 112944 77504 112961
rect 69664 110175 69824 110192
rect 69664 110147 69699 110175
rect 69727 110147 69761 110175
rect 69789 110147 69824 110175
rect 69664 110113 69824 110147
rect 69664 110085 69699 110113
rect 69727 110085 69761 110113
rect 69789 110085 69824 110113
rect 69664 110051 69824 110085
rect 69664 110023 69699 110051
rect 69727 110023 69761 110051
rect 69789 110023 69824 110051
rect 69664 109989 69824 110023
rect 69664 109961 69699 109989
rect 69727 109961 69761 109989
rect 69789 109961 69824 109989
rect 69664 109944 69824 109961
rect 79509 110175 79819 118961
rect 79509 110147 79557 110175
rect 79585 110147 79619 110175
rect 79647 110147 79681 110175
rect 79709 110147 79743 110175
rect 79771 110147 79819 110175
rect 79509 110113 79819 110147
rect 79509 110085 79557 110113
rect 79585 110085 79619 110113
rect 79647 110085 79681 110113
rect 79709 110085 79743 110113
rect 79771 110085 79819 110113
rect 79509 110051 79819 110085
rect 79509 110023 79557 110051
rect 79585 110023 79619 110051
rect 79647 110023 79681 110051
rect 79709 110023 79743 110051
rect 79771 110023 79819 110051
rect 79509 109989 79819 110023
rect 79509 109961 79557 109989
rect 79585 109961 79619 109989
rect 79647 109961 79681 109989
rect 79709 109961 79743 109989
rect 79771 109961 79819 109989
rect 66009 104147 66057 104175
rect 66085 104147 66119 104175
rect 66147 104147 66181 104175
rect 66209 104147 66243 104175
rect 66271 104147 66319 104175
rect 66009 104113 66319 104147
rect 66009 104085 66057 104113
rect 66085 104085 66119 104113
rect 66147 104085 66181 104113
rect 66209 104085 66243 104113
rect 66271 104085 66319 104113
rect 66009 104051 66319 104085
rect 66009 104023 66057 104051
rect 66085 104023 66119 104051
rect 66147 104023 66181 104051
rect 66209 104023 66243 104051
rect 66271 104023 66319 104051
rect 66009 103989 66319 104023
rect 66009 103961 66057 103989
rect 66085 103961 66119 103989
rect 66147 103961 66181 103989
rect 66209 103961 66243 103989
rect 66271 103961 66319 103989
rect 66009 95175 66319 103961
rect 77344 104175 77504 104192
rect 77344 104147 77379 104175
rect 77407 104147 77441 104175
rect 77469 104147 77504 104175
rect 77344 104113 77504 104147
rect 77344 104085 77379 104113
rect 77407 104085 77441 104113
rect 77469 104085 77504 104113
rect 77344 104051 77504 104085
rect 77344 104023 77379 104051
rect 77407 104023 77441 104051
rect 77469 104023 77504 104051
rect 77344 103989 77504 104023
rect 77344 103961 77379 103989
rect 77407 103961 77441 103989
rect 77469 103961 77504 103989
rect 77344 103944 77504 103961
rect 69664 101175 69824 101192
rect 69664 101147 69699 101175
rect 69727 101147 69761 101175
rect 69789 101147 69824 101175
rect 69664 101113 69824 101147
rect 69664 101085 69699 101113
rect 69727 101085 69761 101113
rect 69789 101085 69824 101113
rect 69664 101051 69824 101085
rect 69664 101023 69699 101051
rect 69727 101023 69761 101051
rect 69789 101023 69824 101051
rect 69664 100989 69824 101023
rect 69664 100961 69699 100989
rect 69727 100961 69761 100989
rect 69789 100961 69824 100989
rect 69664 100944 69824 100961
rect 79509 101175 79819 109961
rect 79509 101147 79557 101175
rect 79585 101147 79619 101175
rect 79647 101147 79681 101175
rect 79709 101147 79743 101175
rect 79771 101147 79819 101175
rect 79509 101113 79819 101147
rect 79509 101085 79557 101113
rect 79585 101085 79619 101113
rect 79647 101085 79681 101113
rect 79709 101085 79743 101113
rect 79771 101085 79819 101113
rect 79509 101051 79819 101085
rect 79509 101023 79557 101051
rect 79585 101023 79619 101051
rect 79647 101023 79681 101051
rect 79709 101023 79743 101051
rect 79771 101023 79819 101051
rect 79509 100989 79819 101023
rect 79509 100961 79557 100989
rect 79585 100961 79619 100989
rect 79647 100961 79681 100989
rect 79709 100961 79743 100989
rect 79771 100961 79819 100989
rect 66009 95147 66057 95175
rect 66085 95147 66119 95175
rect 66147 95147 66181 95175
rect 66209 95147 66243 95175
rect 66271 95147 66319 95175
rect 66009 95113 66319 95147
rect 66009 95085 66057 95113
rect 66085 95085 66119 95113
rect 66147 95085 66181 95113
rect 66209 95085 66243 95113
rect 66271 95085 66319 95113
rect 66009 95051 66319 95085
rect 66009 95023 66057 95051
rect 66085 95023 66119 95051
rect 66147 95023 66181 95051
rect 66209 95023 66243 95051
rect 66271 95023 66319 95051
rect 66009 94989 66319 95023
rect 66009 94961 66057 94989
rect 66085 94961 66119 94989
rect 66147 94961 66181 94989
rect 66209 94961 66243 94989
rect 66271 94961 66319 94989
rect 66009 86175 66319 94961
rect 77344 95175 77504 95192
rect 77344 95147 77379 95175
rect 77407 95147 77441 95175
rect 77469 95147 77504 95175
rect 77344 95113 77504 95147
rect 77344 95085 77379 95113
rect 77407 95085 77441 95113
rect 77469 95085 77504 95113
rect 77344 95051 77504 95085
rect 77344 95023 77379 95051
rect 77407 95023 77441 95051
rect 77469 95023 77504 95051
rect 77344 94989 77504 95023
rect 77344 94961 77379 94989
rect 77407 94961 77441 94989
rect 77469 94961 77504 94989
rect 77344 94944 77504 94961
rect 69664 92175 69824 92192
rect 69664 92147 69699 92175
rect 69727 92147 69761 92175
rect 69789 92147 69824 92175
rect 69664 92113 69824 92147
rect 69664 92085 69699 92113
rect 69727 92085 69761 92113
rect 69789 92085 69824 92113
rect 69664 92051 69824 92085
rect 69664 92023 69699 92051
rect 69727 92023 69761 92051
rect 69789 92023 69824 92051
rect 69664 91989 69824 92023
rect 69664 91961 69699 91989
rect 69727 91961 69761 91989
rect 69789 91961 69824 91989
rect 69664 91944 69824 91961
rect 79509 92175 79819 100961
rect 79509 92147 79557 92175
rect 79585 92147 79619 92175
rect 79647 92147 79681 92175
rect 79709 92147 79743 92175
rect 79771 92147 79819 92175
rect 79509 92113 79819 92147
rect 79509 92085 79557 92113
rect 79585 92085 79619 92113
rect 79647 92085 79681 92113
rect 79709 92085 79743 92113
rect 79771 92085 79819 92113
rect 79509 92051 79819 92085
rect 79509 92023 79557 92051
rect 79585 92023 79619 92051
rect 79647 92023 79681 92051
rect 79709 92023 79743 92051
rect 79771 92023 79819 92051
rect 79509 91989 79819 92023
rect 79509 91961 79557 91989
rect 79585 91961 79619 91989
rect 79647 91961 79681 91989
rect 79709 91961 79743 91989
rect 79771 91961 79819 91989
rect 66009 86147 66057 86175
rect 66085 86147 66119 86175
rect 66147 86147 66181 86175
rect 66209 86147 66243 86175
rect 66271 86147 66319 86175
rect 66009 86113 66319 86147
rect 66009 86085 66057 86113
rect 66085 86085 66119 86113
rect 66147 86085 66181 86113
rect 66209 86085 66243 86113
rect 66271 86085 66319 86113
rect 66009 86051 66319 86085
rect 66009 86023 66057 86051
rect 66085 86023 66119 86051
rect 66147 86023 66181 86051
rect 66209 86023 66243 86051
rect 66271 86023 66319 86051
rect 66009 85989 66319 86023
rect 66009 85961 66057 85989
rect 66085 85961 66119 85989
rect 66147 85961 66181 85989
rect 66209 85961 66243 85989
rect 66271 85961 66319 85989
rect 66009 77175 66319 85961
rect 77344 86175 77504 86192
rect 77344 86147 77379 86175
rect 77407 86147 77441 86175
rect 77469 86147 77504 86175
rect 77344 86113 77504 86147
rect 77344 86085 77379 86113
rect 77407 86085 77441 86113
rect 77469 86085 77504 86113
rect 77344 86051 77504 86085
rect 77344 86023 77379 86051
rect 77407 86023 77441 86051
rect 77469 86023 77504 86051
rect 77344 85989 77504 86023
rect 77344 85961 77379 85989
rect 77407 85961 77441 85989
rect 77469 85961 77504 85989
rect 77344 85944 77504 85961
rect 69664 83175 69824 83192
rect 69664 83147 69699 83175
rect 69727 83147 69761 83175
rect 69789 83147 69824 83175
rect 69664 83113 69824 83147
rect 69664 83085 69699 83113
rect 69727 83085 69761 83113
rect 69789 83085 69824 83113
rect 69664 83051 69824 83085
rect 69664 83023 69699 83051
rect 69727 83023 69761 83051
rect 69789 83023 69824 83051
rect 69664 82989 69824 83023
rect 69664 82961 69699 82989
rect 69727 82961 69761 82989
rect 69789 82961 69824 82989
rect 69664 82944 69824 82961
rect 79509 83175 79819 91961
rect 79509 83147 79557 83175
rect 79585 83147 79619 83175
rect 79647 83147 79681 83175
rect 79709 83147 79743 83175
rect 79771 83147 79819 83175
rect 79509 83113 79819 83147
rect 79509 83085 79557 83113
rect 79585 83085 79619 83113
rect 79647 83085 79681 83113
rect 79709 83085 79743 83113
rect 79771 83085 79819 83113
rect 79509 83051 79819 83085
rect 79509 83023 79557 83051
rect 79585 83023 79619 83051
rect 79647 83023 79681 83051
rect 79709 83023 79743 83051
rect 79771 83023 79819 83051
rect 79509 82989 79819 83023
rect 79509 82961 79557 82989
rect 79585 82961 79619 82989
rect 79647 82961 79681 82989
rect 79709 82961 79743 82989
rect 79771 82961 79819 82989
rect 66009 77147 66057 77175
rect 66085 77147 66119 77175
rect 66147 77147 66181 77175
rect 66209 77147 66243 77175
rect 66271 77147 66319 77175
rect 66009 77113 66319 77147
rect 66009 77085 66057 77113
rect 66085 77085 66119 77113
rect 66147 77085 66181 77113
rect 66209 77085 66243 77113
rect 66271 77085 66319 77113
rect 66009 77051 66319 77085
rect 66009 77023 66057 77051
rect 66085 77023 66119 77051
rect 66147 77023 66181 77051
rect 66209 77023 66243 77051
rect 66271 77023 66319 77051
rect 66009 76989 66319 77023
rect 66009 76961 66057 76989
rect 66085 76961 66119 76989
rect 66147 76961 66181 76989
rect 66209 76961 66243 76989
rect 66271 76961 66319 76989
rect 66009 68175 66319 76961
rect 77344 77175 77504 77192
rect 77344 77147 77379 77175
rect 77407 77147 77441 77175
rect 77469 77147 77504 77175
rect 77344 77113 77504 77147
rect 77344 77085 77379 77113
rect 77407 77085 77441 77113
rect 77469 77085 77504 77113
rect 77344 77051 77504 77085
rect 77344 77023 77379 77051
rect 77407 77023 77441 77051
rect 77469 77023 77504 77051
rect 77344 76989 77504 77023
rect 77344 76961 77379 76989
rect 77407 76961 77441 76989
rect 77469 76961 77504 76989
rect 77344 76944 77504 76961
rect 69664 74175 69824 74192
rect 69664 74147 69699 74175
rect 69727 74147 69761 74175
rect 69789 74147 69824 74175
rect 69664 74113 69824 74147
rect 69664 74085 69699 74113
rect 69727 74085 69761 74113
rect 69789 74085 69824 74113
rect 69664 74051 69824 74085
rect 69664 74023 69699 74051
rect 69727 74023 69761 74051
rect 69789 74023 69824 74051
rect 69664 73989 69824 74023
rect 69664 73961 69699 73989
rect 69727 73961 69761 73989
rect 69789 73961 69824 73989
rect 69664 73944 69824 73961
rect 79509 74175 79819 82961
rect 79509 74147 79557 74175
rect 79585 74147 79619 74175
rect 79647 74147 79681 74175
rect 79709 74147 79743 74175
rect 79771 74147 79819 74175
rect 79509 74113 79819 74147
rect 79509 74085 79557 74113
rect 79585 74085 79619 74113
rect 79647 74085 79681 74113
rect 79709 74085 79743 74113
rect 79771 74085 79819 74113
rect 79509 74051 79819 74085
rect 79509 74023 79557 74051
rect 79585 74023 79619 74051
rect 79647 74023 79681 74051
rect 79709 74023 79743 74051
rect 79771 74023 79819 74051
rect 79509 73989 79819 74023
rect 79509 73961 79557 73989
rect 79585 73961 79619 73989
rect 79647 73961 79681 73989
rect 79709 73961 79743 73989
rect 79771 73961 79819 73989
rect 66009 68147 66057 68175
rect 66085 68147 66119 68175
rect 66147 68147 66181 68175
rect 66209 68147 66243 68175
rect 66271 68147 66319 68175
rect 66009 68113 66319 68147
rect 66009 68085 66057 68113
rect 66085 68085 66119 68113
rect 66147 68085 66181 68113
rect 66209 68085 66243 68113
rect 66271 68085 66319 68113
rect 66009 68051 66319 68085
rect 66009 68023 66057 68051
rect 66085 68023 66119 68051
rect 66147 68023 66181 68051
rect 66209 68023 66243 68051
rect 66271 68023 66319 68051
rect 66009 67989 66319 68023
rect 66009 67961 66057 67989
rect 66085 67961 66119 67989
rect 66147 67961 66181 67989
rect 66209 67961 66243 67989
rect 66271 67961 66319 67989
rect 66009 59175 66319 67961
rect 77344 68175 77504 68192
rect 77344 68147 77379 68175
rect 77407 68147 77441 68175
rect 77469 68147 77504 68175
rect 77344 68113 77504 68147
rect 77344 68085 77379 68113
rect 77407 68085 77441 68113
rect 77469 68085 77504 68113
rect 77344 68051 77504 68085
rect 77344 68023 77379 68051
rect 77407 68023 77441 68051
rect 77469 68023 77504 68051
rect 77344 67989 77504 68023
rect 77344 67961 77379 67989
rect 77407 67961 77441 67989
rect 77469 67961 77504 67989
rect 77344 67944 77504 67961
rect 69664 65175 69824 65192
rect 69664 65147 69699 65175
rect 69727 65147 69761 65175
rect 69789 65147 69824 65175
rect 69664 65113 69824 65147
rect 69664 65085 69699 65113
rect 69727 65085 69761 65113
rect 69789 65085 69824 65113
rect 69664 65051 69824 65085
rect 69664 65023 69699 65051
rect 69727 65023 69761 65051
rect 69789 65023 69824 65051
rect 69664 64989 69824 65023
rect 69664 64961 69699 64989
rect 69727 64961 69761 64989
rect 69789 64961 69824 64989
rect 69664 64944 69824 64961
rect 79509 65175 79819 73961
rect 79509 65147 79557 65175
rect 79585 65147 79619 65175
rect 79647 65147 79681 65175
rect 79709 65147 79743 65175
rect 79771 65147 79819 65175
rect 79509 65113 79819 65147
rect 79509 65085 79557 65113
rect 79585 65085 79619 65113
rect 79647 65085 79681 65113
rect 79709 65085 79743 65113
rect 79771 65085 79819 65113
rect 79509 65051 79819 65085
rect 79509 65023 79557 65051
rect 79585 65023 79619 65051
rect 79647 65023 79681 65051
rect 79709 65023 79743 65051
rect 79771 65023 79819 65051
rect 79509 64989 79819 65023
rect 79509 64961 79557 64989
rect 79585 64961 79619 64989
rect 79647 64961 79681 64989
rect 79709 64961 79743 64989
rect 79771 64961 79819 64989
rect 66009 59147 66057 59175
rect 66085 59147 66119 59175
rect 66147 59147 66181 59175
rect 66209 59147 66243 59175
rect 66271 59147 66319 59175
rect 66009 59113 66319 59147
rect 66009 59085 66057 59113
rect 66085 59085 66119 59113
rect 66147 59085 66181 59113
rect 66209 59085 66243 59113
rect 66271 59085 66319 59113
rect 66009 59051 66319 59085
rect 66009 59023 66057 59051
rect 66085 59023 66119 59051
rect 66147 59023 66181 59051
rect 66209 59023 66243 59051
rect 66271 59023 66319 59051
rect 66009 58989 66319 59023
rect 66009 58961 66057 58989
rect 66085 58961 66119 58989
rect 66147 58961 66181 58989
rect 66209 58961 66243 58989
rect 66271 58961 66319 58989
rect 66009 50175 66319 58961
rect 77344 59175 77504 59192
rect 77344 59147 77379 59175
rect 77407 59147 77441 59175
rect 77469 59147 77504 59175
rect 77344 59113 77504 59147
rect 77344 59085 77379 59113
rect 77407 59085 77441 59113
rect 77469 59085 77504 59113
rect 77344 59051 77504 59085
rect 77344 59023 77379 59051
rect 77407 59023 77441 59051
rect 77469 59023 77504 59051
rect 77344 58989 77504 59023
rect 77344 58961 77379 58989
rect 77407 58961 77441 58989
rect 77469 58961 77504 58989
rect 77344 58944 77504 58961
rect 69664 56175 69824 56192
rect 69664 56147 69699 56175
rect 69727 56147 69761 56175
rect 69789 56147 69824 56175
rect 69664 56113 69824 56147
rect 69664 56085 69699 56113
rect 69727 56085 69761 56113
rect 69789 56085 69824 56113
rect 69664 56051 69824 56085
rect 69664 56023 69699 56051
rect 69727 56023 69761 56051
rect 69789 56023 69824 56051
rect 69664 55989 69824 56023
rect 69664 55961 69699 55989
rect 69727 55961 69761 55989
rect 69789 55961 69824 55989
rect 69664 55944 69824 55961
rect 79509 56175 79819 64961
rect 79509 56147 79557 56175
rect 79585 56147 79619 56175
rect 79647 56147 79681 56175
rect 79709 56147 79743 56175
rect 79771 56147 79819 56175
rect 79509 56113 79819 56147
rect 79509 56085 79557 56113
rect 79585 56085 79619 56113
rect 79647 56085 79681 56113
rect 79709 56085 79743 56113
rect 79771 56085 79819 56113
rect 79509 56051 79819 56085
rect 79509 56023 79557 56051
rect 79585 56023 79619 56051
rect 79647 56023 79681 56051
rect 79709 56023 79743 56051
rect 79771 56023 79819 56051
rect 79509 55989 79819 56023
rect 79509 55961 79557 55989
rect 79585 55961 79619 55989
rect 79647 55961 79681 55989
rect 79709 55961 79743 55989
rect 79771 55961 79819 55989
rect 66009 50147 66057 50175
rect 66085 50147 66119 50175
rect 66147 50147 66181 50175
rect 66209 50147 66243 50175
rect 66271 50147 66319 50175
rect 66009 50113 66319 50147
rect 66009 50085 66057 50113
rect 66085 50085 66119 50113
rect 66147 50085 66181 50113
rect 66209 50085 66243 50113
rect 66271 50085 66319 50113
rect 66009 50051 66319 50085
rect 66009 50023 66057 50051
rect 66085 50023 66119 50051
rect 66147 50023 66181 50051
rect 66209 50023 66243 50051
rect 66271 50023 66319 50051
rect 66009 49989 66319 50023
rect 66009 49961 66057 49989
rect 66085 49961 66119 49989
rect 66147 49961 66181 49989
rect 66209 49961 66243 49989
rect 66271 49961 66319 49989
rect 66009 41175 66319 49961
rect 77344 50175 77504 50192
rect 77344 50147 77379 50175
rect 77407 50147 77441 50175
rect 77469 50147 77504 50175
rect 77344 50113 77504 50147
rect 77344 50085 77379 50113
rect 77407 50085 77441 50113
rect 77469 50085 77504 50113
rect 77344 50051 77504 50085
rect 77344 50023 77379 50051
rect 77407 50023 77441 50051
rect 77469 50023 77504 50051
rect 77344 49989 77504 50023
rect 77344 49961 77379 49989
rect 77407 49961 77441 49989
rect 77469 49961 77504 49989
rect 77344 49944 77504 49961
rect 69664 47175 69824 47192
rect 69664 47147 69699 47175
rect 69727 47147 69761 47175
rect 69789 47147 69824 47175
rect 69664 47113 69824 47147
rect 69664 47085 69699 47113
rect 69727 47085 69761 47113
rect 69789 47085 69824 47113
rect 69664 47051 69824 47085
rect 69664 47023 69699 47051
rect 69727 47023 69761 47051
rect 69789 47023 69824 47051
rect 69664 46989 69824 47023
rect 69664 46961 69699 46989
rect 69727 46961 69761 46989
rect 69789 46961 69824 46989
rect 69664 46944 69824 46961
rect 79509 47175 79819 55961
rect 79509 47147 79557 47175
rect 79585 47147 79619 47175
rect 79647 47147 79681 47175
rect 79709 47147 79743 47175
rect 79771 47147 79819 47175
rect 79509 47113 79819 47147
rect 79509 47085 79557 47113
rect 79585 47085 79619 47113
rect 79647 47085 79681 47113
rect 79709 47085 79743 47113
rect 79771 47085 79819 47113
rect 79509 47051 79819 47085
rect 79509 47023 79557 47051
rect 79585 47023 79619 47051
rect 79647 47023 79681 47051
rect 79709 47023 79743 47051
rect 79771 47023 79819 47051
rect 79509 46989 79819 47023
rect 79509 46961 79557 46989
rect 79585 46961 79619 46989
rect 79647 46961 79681 46989
rect 79709 46961 79743 46989
rect 79771 46961 79819 46989
rect 66009 41147 66057 41175
rect 66085 41147 66119 41175
rect 66147 41147 66181 41175
rect 66209 41147 66243 41175
rect 66271 41147 66319 41175
rect 66009 41113 66319 41147
rect 66009 41085 66057 41113
rect 66085 41085 66119 41113
rect 66147 41085 66181 41113
rect 66209 41085 66243 41113
rect 66271 41085 66319 41113
rect 66009 41051 66319 41085
rect 66009 41023 66057 41051
rect 66085 41023 66119 41051
rect 66147 41023 66181 41051
rect 66209 41023 66243 41051
rect 66271 41023 66319 41051
rect 66009 40989 66319 41023
rect 66009 40961 66057 40989
rect 66085 40961 66119 40989
rect 66147 40961 66181 40989
rect 66209 40961 66243 40989
rect 66271 40961 66319 40989
rect 66009 32175 66319 40961
rect 77344 41175 77504 41192
rect 77344 41147 77379 41175
rect 77407 41147 77441 41175
rect 77469 41147 77504 41175
rect 77344 41113 77504 41147
rect 77344 41085 77379 41113
rect 77407 41085 77441 41113
rect 77469 41085 77504 41113
rect 77344 41051 77504 41085
rect 77344 41023 77379 41051
rect 77407 41023 77441 41051
rect 77469 41023 77504 41051
rect 77344 40989 77504 41023
rect 77344 40961 77379 40989
rect 77407 40961 77441 40989
rect 77469 40961 77504 40989
rect 77344 40944 77504 40961
rect 69664 38175 69824 38192
rect 69664 38147 69699 38175
rect 69727 38147 69761 38175
rect 69789 38147 69824 38175
rect 69664 38113 69824 38147
rect 69664 38085 69699 38113
rect 69727 38085 69761 38113
rect 69789 38085 69824 38113
rect 69664 38051 69824 38085
rect 69664 38023 69699 38051
rect 69727 38023 69761 38051
rect 69789 38023 69824 38051
rect 69664 37989 69824 38023
rect 69664 37961 69699 37989
rect 69727 37961 69761 37989
rect 69789 37961 69824 37989
rect 69664 37944 69824 37961
rect 79509 38175 79819 46961
rect 79509 38147 79557 38175
rect 79585 38147 79619 38175
rect 79647 38147 79681 38175
rect 79709 38147 79743 38175
rect 79771 38147 79819 38175
rect 79509 38113 79819 38147
rect 79509 38085 79557 38113
rect 79585 38085 79619 38113
rect 79647 38085 79681 38113
rect 79709 38085 79743 38113
rect 79771 38085 79819 38113
rect 79509 38051 79819 38085
rect 79509 38023 79557 38051
rect 79585 38023 79619 38051
rect 79647 38023 79681 38051
rect 79709 38023 79743 38051
rect 79771 38023 79819 38051
rect 79509 37989 79819 38023
rect 79509 37961 79557 37989
rect 79585 37961 79619 37989
rect 79647 37961 79681 37989
rect 79709 37961 79743 37989
rect 79771 37961 79819 37989
rect 66009 32147 66057 32175
rect 66085 32147 66119 32175
rect 66147 32147 66181 32175
rect 66209 32147 66243 32175
rect 66271 32147 66319 32175
rect 66009 32113 66319 32147
rect 66009 32085 66057 32113
rect 66085 32085 66119 32113
rect 66147 32085 66181 32113
rect 66209 32085 66243 32113
rect 66271 32085 66319 32113
rect 66009 32051 66319 32085
rect 66009 32023 66057 32051
rect 66085 32023 66119 32051
rect 66147 32023 66181 32051
rect 66209 32023 66243 32051
rect 66271 32023 66319 32051
rect 66009 31989 66319 32023
rect 66009 31961 66057 31989
rect 66085 31961 66119 31989
rect 66147 31961 66181 31989
rect 66209 31961 66243 31989
rect 66271 31961 66319 31989
rect 66009 23175 66319 31961
rect 77344 32175 77504 32192
rect 77344 32147 77379 32175
rect 77407 32147 77441 32175
rect 77469 32147 77504 32175
rect 77344 32113 77504 32147
rect 77344 32085 77379 32113
rect 77407 32085 77441 32113
rect 77469 32085 77504 32113
rect 77344 32051 77504 32085
rect 77344 32023 77379 32051
rect 77407 32023 77441 32051
rect 77469 32023 77504 32051
rect 77344 31989 77504 32023
rect 77344 31961 77379 31989
rect 77407 31961 77441 31989
rect 77469 31961 77504 31989
rect 77344 31944 77504 31961
rect 69664 29175 69824 29192
rect 69664 29147 69699 29175
rect 69727 29147 69761 29175
rect 69789 29147 69824 29175
rect 69664 29113 69824 29147
rect 69664 29085 69699 29113
rect 69727 29085 69761 29113
rect 69789 29085 69824 29113
rect 69664 29051 69824 29085
rect 69664 29023 69699 29051
rect 69727 29023 69761 29051
rect 69789 29023 69824 29051
rect 69664 28989 69824 29023
rect 69664 28961 69699 28989
rect 69727 28961 69761 28989
rect 69789 28961 69824 28989
rect 69664 28944 69824 28961
rect 79509 29175 79819 37961
rect 79509 29147 79557 29175
rect 79585 29147 79619 29175
rect 79647 29147 79681 29175
rect 79709 29147 79743 29175
rect 79771 29147 79819 29175
rect 79509 29113 79819 29147
rect 79509 29085 79557 29113
rect 79585 29085 79619 29113
rect 79647 29085 79681 29113
rect 79709 29085 79743 29113
rect 79771 29085 79819 29113
rect 79509 29051 79819 29085
rect 79509 29023 79557 29051
rect 79585 29023 79619 29051
rect 79647 29023 79681 29051
rect 79709 29023 79743 29051
rect 79771 29023 79819 29051
rect 79509 28989 79819 29023
rect 79509 28961 79557 28989
rect 79585 28961 79619 28989
rect 79647 28961 79681 28989
rect 79709 28961 79743 28989
rect 79771 28961 79819 28989
rect 66009 23147 66057 23175
rect 66085 23147 66119 23175
rect 66147 23147 66181 23175
rect 66209 23147 66243 23175
rect 66271 23147 66319 23175
rect 66009 23113 66319 23147
rect 66009 23085 66057 23113
rect 66085 23085 66119 23113
rect 66147 23085 66181 23113
rect 66209 23085 66243 23113
rect 66271 23085 66319 23113
rect 66009 23051 66319 23085
rect 66009 23023 66057 23051
rect 66085 23023 66119 23051
rect 66147 23023 66181 23051
rect 66209 23023 66243 23051
rect 66271 23023 66319 23051
rect 66009 22989 66319 23023
rect 66009 22961 66057 22989
rect 66085 22961 66119 22989
rect 66147 22961 66181 22989
rect 66209 22961 66243 22989
rect 66271 22961 66319 22989
rect 66009 14175 66319 22961
rect 77344 23175 77504 23192
rect 77344 23147 77379 23175
rect 77407 23147 77441 23175
rect 77469 23147 77504 23175
rect 77344 23113 77504 23147
rect 77344 23085 77379 23113
rect 77407 23085 77441 23113
rect 77469 23085 77504 23113
rect 77344 23051 77504 23085
rect 77344 23023 77379 23051
rect 77407 23023 77441 23051
rect 77469 23023 77504 23051
rect 77344 22989 77504 23023
rect 77344 22961 77379 22989
rect 77407 22961 77441 22989
rect 77469 22961 77504 22989
rect 77344 22944 77504 22961
rect 69664 20175 69824 20192
rect 69664 20147 69699 20175
rect 69727 20147 69761 20175
rect 69789 20147 69824 20175
rect 69664 20113 69824 20147
rect 69664 20085 69699 20113
rect 69727 20085 69761 20113
rect 69789 20085 69824 20113
rect 69664 20051 69824 20085
rect 69664 20023 69699 20051
rect 69727 20023 69761 20051
rect 69789 20023 69824 20051
rect 69664 19989 69824 20023
rect 69664 19961 69699 19989
rect 69727 19961 69761 19989
rect 69789 19961 69824 19989
rect 69664 19944 69824 19961
rect 79509 20175 79819 28961
rect 79509 20147 79557 20175
rect 79585 20147 79619 20175
rect 79647 20147 79681 20175
rect 79709 20147 79743 20175
rect 79771 20147 79819 20175
rect 79509 20113 79819 20147
rect 79509 20085 79557 20113
rect 79585 20085 79619 20113
rect 79647 20085 79681 20113
rect 79709 20085 79743 20113
rect 79771 20085 79819 20113
rect 79509 20051 79819 20085
rect 79509 20023 79557 20051
rect 79585 20023 79619 20051
rect 79647 20023 79681 20051
rect 79709 20023 79743 20051
rect 79771 20023 79819 20051
rect 79509 19989 79819 20023
rect 79509 19961 79557 19989
rect 79585 19961 79619 19989
rect 79647 19961 79681 19989
rect 79709 19961 79743 19989
rect 79771 19961 79819 19989
rect 66009 14147 66057 14175
rect 66085 14147 66119 14175
rect 66147 14147 66181 14175
rect 66209 14147 66243 14175
rect 66271 14147 66319 14175
rect 66009 14113 66319 14147
rect 66009 14085 66057 14113
rect 66085 14085 66119 14113
rect 66147 14085 66181 14113
rect 66209 14085 66243 14113
rect 66271 14085 66319 14113
rect 66009 14051 66319 14085
rect 66009 14023 66057 14051
rect 66085 14023 66119 14051
rect 66147 14023 66181 14051
rect 66209 14023 66243 14051
rect 66271 14023 66319 14051
rect 66009 13989 66319 14023
rect 66009 13961 66057 13989
rect 66085 13961 66119 13989
rect 66147 13961 66181 13989
rect 66209 13961 66243 13989
rect 66271 13961 66319 13989
rect 66009 5175 66319 13961
rect 77344 14175 77504 14192
rect 77344 14147 77379 14175
rect 77407 14147 77441 14175
rect 77469 14147 77504 14175
rect 77344 14113 77504 14147
rect 77344 14085 77379 14113
rect 77407 14085 77441 14113
rect 77469 14085 77504 14113
rect 77344 14051 77504 14085
rect 77344 14023 77379 14051
rect 77407 14023 77441 14051
rect 77469 14023 77504 14051
rect 77344 13989 77504 14023
rect 77344 13961 77379 13989
rect 77407 13961 77441 13989
rect 77469 13961 77504 13989
rect 77344 13944 77504 13961
rect 69664 11175 69824 11192
rect 69664 11147 69699 11175
rect 69727 11147 69761 11175
rect 69789 11147 69824 11175
rect 69664 11113 69824 11147
rect 69664 11085 69699 11113
rect 69727 11085 69761 11113
rect 69789 11085 69824 11113
rect 69664 11051 69824 11085
rect 69664 11023 69699 11051
rect 69727 11023 69761 11051
rect 69789 11023 69824 11051
rect 69664 10989 69824 11023
rect 69664 10961 69699 10989
rect 69727 10961 69761 10989
rect 69789 10961 69824 10989
rect 69664 10944 69824 10961
rect 79509 11175 79819 19961
rect 79509 11147 79557 11175
rect 79585 11147 79619 11175
rect 79647 11147 79681 11175
rect 79709 11147 79743 11175
rect 79771 11147 79819 11175
rect 79509 11113 79819 11147
rect 79509 11085 79557 11113
rect 79585 11085 79619 11113
rect 79647 11085 79681 11113
rect 79709 11085 79743 11113
rect 79771 11085 79819 11113
rect 79509 11051 79819 11085
rect 79509 11023 79557 11051
rect 79585 11023 79619 11051
rect 79647 11023 79681 11051
rect 79709 11023 79743 11051
rect 79771 11023 79819 11051
rect 79509 10989 79819 11023
rect 79509 10961 79557 10989
rect 79585 10961 79619 10989
rect 79647 10961 79681 10989
rect 79709 10961 79743 10989
rect 79771 10961 79819 10989
rect 66009 5147 66057 5175
rect 66085 5147 66119 5175
rect 66147 5147 66181 5175
rect 66209 5147 66243 5175
rect 66271 5147 66319 5175
rect 66009 5113 66319 5147
rect 66009 5085 66057 5113
rect 66085 5085 66119 5113
rect 66147 5085 66181 5113
rect 66209 5085 66243 5113
rect 66271 5085 66319 5113
rect 66009 5051 66319 5085
rect 66009 5023 66057 5051
rect 66085 5023 66119 5051
rect 66147 5023 66181 5051
rect 66209 5023 66243 5051
rect 66271 5023 66319 5051
rect 66009 4989 66319 5023
rect 66009 4961 66057 4989
rect 66085 4961 66119 4989
rect 66147 4961 66181 4989
rect 66209 4961 66243 4989
rect 66271 4961 66319 4989
rect 66009 -560 66319 4961
rect 77344 5175 77504 5192
rect 77344 5147 77379 5175
rect 77407 5147 77441 5175
rect 77469 5147 77504 5175
rect 77344 5113 77504 5147
rect 77344 5085 77379 5113
rect 77407 5085 77441 5113
rect 77469 5085 77504 5113
rect 77344 5051 77504 5085
rect 77344 5023 77379 5051
rect 77407 5023 77441 5051
rect 77469 5023 77504 5051
rect 77344 4989 77504 5023
rect 77344 4961 77379 4989
rect 77407 4961 77441 4989
rect 77469 4961 77504 4989
rect 77344 4944 77504 4961
rect 66009 -588 66057 -560
rect 66085 -588 66119 -560
rect 66147 -588 66181 -560
rect 66209 -588 66243 -560
rect 66271 -588 66319 -560
rect 66009 -622 66319 -588
rect 66009 -650 66057 -622
rect 66085 -650 66119 -622
rect 66147 -650 66181 -622
rect 66209 -650 66243 -622
rect 66271 -650 66319 -622
rect 66009 -684 66319 -650
rect 66009 -712 66057 -684
rect 66085 -712 66119 -684
rect 66147 -712 66181 -684
rect 66209 -712 66243 -684
rect 66271 -712 66319 -684
rect 66009 -746 66319 -712
rect 66009 -774 66057 -746
rect 66085 -774 66119 -746
rect 66147 -774 66181 -746
rect 66209 -774 66243 -746
rect 66271 -774 66319 -746
rect 66009 -822 66319 -774
rect 79509 2175 79819 10961
rect 79509 2147 79557 2175
rect 79585 2147 79619 2175
rect 79647 2147 79681 2175
rect 79709 2147 79743 2175
rect 79771 2147 79819 2175
rect 79509 2113 79819 2147
rect 79509 2085 79557 2113
rect 79585 2085 79619 2113
rect 79647 2085 79681 2113
rect 79709 2085 79743 2113
rect 79771 2085 79819 2113
rect 79509 2051 79819 2085
rect 79509 2023 79557 2051
rect 79585 2023 79619 2051
rect 79647 2023 79681 2051
rect 79709 2023 79743 2051
rect 79771 2023 79819 2051
rect 79509 1989 79819 2023
rect 79509 1961 79557 1989
rect 79585 1961 79619 1989
rect 79647 1961 79681 1989
rect 79709 1961 79743 1989
rect 79771 1961 79819 1989
rect 79509 -80 79819 1961
rect 79509 -108 79557 -80
rect 79585 -108 79619 -80
rect 79647 -108 79681 -80
rect 79709 -108 79743 -80
rect 79771 -108 79819 -80
rect 79509 -142 79819 -108
rect 79509 -170 79557 -142
rect 79585 -170 79619 -142
rect 79647 -170 79681 -142
rect 79709 -170 79743 -142
rect 79771 -170 79819 -142
rect 79509 -204 79819 -170
rect 79509 -232 79557 -204
rect 79585 -232 79619 -204
rect 79647 -232 79681 -204
rect 79709 -232 79743 -204
rect 79771 -232 79819 -204
rect 79509 -266 79819 -232
rect 79509 -294 79557 -266
rect 79585 -294 79619 -266
rect 79647 -294 79681 -266
rect 79709 -294 79743 -266
rect 79771 -294 79819 -266
rect 79509 -822 79819 -294
rect 81369 299086 81679 299134
rect 81369 299058 81417 299086
rect 81445 299058 81479 299086
rect 81507 299058 81541 299086
rect 81569 299058 81603 299086
rect 81631 299058 81679 299086
rect 81369 299024 81679 299058
rect 81369 298996 81417 299024
rect 81445 298996 81479 299024
rect 81507 298996 81541 299024
rect 81569 298996 81603 299024
rect 81631 298996 81679 299024
rect 81369 298962 81679 298996
rect 81369 298934 81417 298962
rect 81445 298934 81479 298962
rect 81507 298934 81541 298962
rect 81569 298934 81603 298962
rect 81631 298934 81679 298962
rect 81369 298900 81679 298934
rect 81369 298872 81417 298900
rect 81445 298872 81479 298900
rect 81507 298872 81541 298900
rect 81569 298872 81603 298900
rect 81631 298872 81679 298900
rect 81369 293175 81679 298872
rect 81369 293147 81417 293175
rect 81445 293147 81479 293175
rect 81507 293147 81541 293175
rect 81569 293147 81603 293175
rect 81631 293147 81679 293175
rect 81369 293113 81679 293147
rect 81369 293085 81417 293113
rect 81445 293085 81479 293113
rect 81507 293085 81541 293113
rect 81569 293085 81603 293113
rect 81631 293085 81679 293113
rect 81369 293051 81679 293085
rect 81369 293023 81417 293051
rect 81445 293023 81479 293051
rect 81507 293023 81541 293051
rect 81569 293023 81603 293051
rect 81631 293023 81679 293051
rect 81369 292989 81679 293023
rect 81369 292961 81417 292989
rect 81445 292961 81479 292989
rect 81507 292961 81541 292989
rect 81569 292961 81603 292989
rect 81631 292961 81679 292989
rect 81369 284175 81679 292961
rect 81369 284147 81417 284175
rect 81445 284147 81479 284175
rect 81507 284147 81541 284175
rect 81569 284147 81603 284175
rect 81631 284147 81679 284175
rect 81369 284113 81679 284147
rect 81369 284085 81417 284113
rect 81445 284085 81479 284113
rect 81507 284085 81541 284113
rect 81569 284085 81603 284113
rect 81631 284085 81679 284113
rect 81369 284051 81679 284085
rect 81369 284023 81417 284051
rect 81445 284023 81479 284051
rect 81507 284023 81541 284051
rect 81569 284023 81603 284051
rect 81631 284023 81679 284051
rect 81369 283989 81679 284023
rect 81369 283961 81417 283989
rect 81445 283961 81479 283989
rect 81507 283961 81541 283989
rect 81569 283961 81603 283989
rect 81631 283961 81679 283989
rect 81369 275175 81679 283961
rect 81369 275147 81417 275175
rect 81445 275147 81479 275175
rect 81507 275147 81541 275175
rect 81569 275147 81603 275175
rect 81631 275147 81679 275175
rect 81369 275113 81679 275147
rect 81369 275085 81417 275113
rect 81445 275085 81479 275113
rect 81507 275085 81541 275113
rect 81569 275085 81603 275113
rect 81631 275085 81679 275113
rect 81369 275051 81679 275085
rect 81369 275023 81417 275051
rect 81445 275023 81479 275051
rect 81507 275023 81541 275051
rect 81569 275023 81603 275051
rect 81631 275023 81679 275051
rect 81369 274989 81679 275023
rect 81369 274961 81417 274989
rect 81445 274961 81479 274989
rect 81507 274961 81541 274989
rect 81569 274961 81603 274989
rect 81631 274961 81679 274989
rect 81369 266175 81679 274961
rect 81369 266147 81417 266175
rect 81445 266147 81479 266175
rect 81507 266147 81541 266175
rect 81569 266147 81603 266175
rect 81631 266147 81679 266175
rect 81369 266113 81679 266147
rect 81369 266085 81417 266113
rect 81445 266085 81479 266113
rect 81507 266085 81541 266113
rect 81569 266085 81603 266113
rect 81631 266085 81679 266113
rect 81369 266051 81679 266085
rect 81369 266023 81417 266051
rect 81445 266023 81479 266051
rect 81507 266023 81541 266051
rect 81569 266023 81603 266051
rect 81631 266023 81679 266051
rect 81369 265989 81679 266023
rect 81369 265961 81417 265989
rect 81445 265961 81479 265989
rect 81507 265961 81541 265989
rect 81569 265961 81603 265989
rect 81631 265961 81679 265989
rect 81369 257175 81679 265961
rect 81369 257147 81417 257175
rect 81445 257147 81479 257175
rect 81507 257147 81541 257175
rect 81569 257147 81603 257175
rect 81631 257147 81679 257175
rect 81369 257113 81679 257147
rect 81369 257085 81417 257113
rect 81445 257085 81479 257113
rect 81507 257085 81541 257113
rect 81569 257085 81603 257113
rect 81631 257085 81679 257113
rect 81369 257051 81679 257085
rect 81369 257023 81417 257051
rect 81445 257023 81479 257051
rect 81507 257023 81541 257051
rect 81569 257023 81603 257051
rect 81631 257023 81679 257051
rect 81369 256989 81679 257023
rect 81369 256961 81417 256989
rect 81445 256961 81479 256989
rect 81507 256961 81541 256989
rect 81569 256961 81603 256989
rect 81631 256961 81679 256989
rect 81369 248175 81679 256961
rect 81369 248147 81417 248175
rect 81445 248147 81479 248175
rect 81507 248147 81541 248175
rect 81569 248147 81603 248175
rect 81631 248147 81679 248175
rect 81369 248113 81679 248147
rect 81369 248085 81417 248113
rect 81445 248085 81479 248113
rect 81507 248085 81541 248113
rect 81569 248085 81603 248113
rect 81631 248085 81679 248113
rect 81369 248051 81679 248085
rect 81369 248023 81417 248051
rect 81445 248023 81479 248051
rect 81507 248023 81541 248051
rect 81569 248023 81603 248051
rect 81631 248023 81679 248051
rect 81369 247989 81679 248023
rect 81369 247961 81417 247989
rect 81445 247961 81479 247989
rect 81507 247961 81541 247989
rect 81569 247961 81603 247989
rect 81631 247961 81679 247989
rect 81369 239175 81679 247961
rect 81369 239147 81417 239175
rect 81445 239147 81479 239175
rect 81507 239147 81541 239175
rect 81569 239147 81603 239175
rect 81631 239147 81679 239175
rect 81369 239113 81679 239147
rect 81369 239085 81417 239113
rect 81445 239085 81479 239113
rect 81507 239085 81541 239113
rect 81569 239085 81603 239113
rect 81631 239085 81679 239113
rect 81369 239051 81679 239085
rect 81369 239023 81417 239051
rect 81445 239023 81479 239051
rect 81507 239023 81541 239051
rect 81569 239023 81603 239051
rect 81631 239023 81679 239051
rect 81369 238989 81679 239023
rect 81369 238961 81417 238989
rect 81445 238961 81479 238989
rect 81507 238961 81541 238989
rect 81569 238961 81603 238989
rect 81631 238961 81679 238989
rect 81369 230175 81679 238961
rect 81369 230147 81417 230175
rect 81445 230147 81479 230175
rect 81507 230147 81541 230175
rect 81569 230147 81603 230175
rect 81631 230147 81679 230175
rect 81369 230113 81679 230147
rect 81369 230085 81417 230113
rect 81445 230085 81479 230113
rect 81507 230085 81541 230113
rect 81569 230085 81603 230113
rect 81631 230085 81679 230113
rect 81369 230051 81679 230085
rect 81369 230023 81417 230051
rect 81445 230023 81479 230051
rect 81507 230023 81541 230051
rect 81569 230023 81603 230051
rect 81631 230023 81679 230051
rect 81369 229989 81679 230023
rect 81369 229961 81417 229989
rect 81445 229961 81479 229989
rect 81507 229961 81541 229989
rect 81569 229961 81603 229989
rect 81631 229961 81679 229989
rect 81369 221175 81679 229961
rect 81369 221147 81417 221175
rect 81445 221147 81479 221175
rect 81507 221147 81541 221175
rect 81569 221147 81603 221175
rect 81631 221147 81679 221175
rect 81369 221113 81679 221147
rect 81369 221085 81417 221113
rect 81445 221085 81479 221113
rect 81507 221085 81541 221113
rect 81569 221085 81603 221113
rect 81631 221085 81679 221113
rect 81369 221051 81679 221085
rect 81369 221023 81417 221051
rect 81445 221023 81479 221051
rect 81507 221023 81541 221051
rect 81569 221023 81603 221051
rect 81631 221023 81679 221051
rect 81369 220989 81679 221023
rect 81369 220961 81417 220989
rect 81445 220961 81479 220989
rect 81507 220961 81541 220989
rect 81569 220961 81603 220989
rect 81631 220961 81679 220989
rect 81369 212175 81679 220961
rect 81369 212147 81417 212175
rect 81445 212147 81479 212175
rect 81507 212147 81541 212175
rect 81569 212147 81603 212175
rect 81631 212147 81679 212175
rect 81369 212113 81679 212147
rect 81369 212085 81417 212113
rect 81445 212085 81479 212113
rect 81507 212085 81541 212113
rect 81569 212085 81603 212113
rect 81631 212085 81679 212113
rect 81369 212051 81679 212085
rect 81369 212023 81417 212051
rect 81445 212023 81479 212051
rect 81507 212023 81541 212051
rect 81569 212023 81603 212051
rect 81631 212023 81679 212051
rect 81369 211989 81679 212023
rect 81369 211961 81417 211989
rect 81445 211961 81479 211989
rect 81507 211961 81541 211989
rect 81569 211961 81603 211989
rect 81631 211961 81679 211989
rect 81369 203175 81679 211961
rect 81369 203147 81417 203175
rect 81445 203147 81479 203175
rect 81507 203147 81541 203175
rect 81569 203147 81603 203175
rect 81631 203147 81679 203175
rect 81369 203113 81679 203147
rect 81369 203085 81417 203113
rect 81445 203085 81479 203113
rect 81507 203085 81541 203113
rect 81569 203085 81603 203113
rect 81631 203085 81679 203113
rect 81369 203051 81679 203085
rect 81369 203023 81417 203051
rect 81445 203023 81479 203051
rect 81507 203023 81541 203051
rect 81569 203023 81603 203051
rect 81631 203023 81679 203051
rect 81369 202989 81679 203023
rect 81369 202961 81417 202989
rect 81445 202961 81479 202989
rect 81507 202961 81541 202989
rect 81569 202961 81603 202989
rect 81631 202961 81679 202989
rect 81369 194175 81679 202961
rect 81369 194147 81417 194175
rect 81445 194147 81479 194175
rect 81507 194147 81541 194175
rect 81569 194147 81603 194175
rect 81631 194147 81679 194175
rect 81369 194113 81679 194147
rect 81369 194085 81417 194113
rect 81445 194085 81479 194113
rect 81507 194085 81541 194113
rect 81569 194085 81603 194113
rect 81631 194085 81679 194113
rect 81369 194051 81679 194085
rect 81369 194023 81417 194051
rect 81445 194023 81479 194051
rect 81507 194023 81541 194051
rect 81569 194023 81603 194051
rect 81631 194023 81679 194051
rect 81369 193989 81679 194023
rect 81369 193961 81417 193989
rect 81445 193961 81479 193989
rect 81507 193961 81541 193989
rect 81569 193961 81603 193989
rect 81631 193961 81679 193989
rect 81369 185175 81679 193961
rect 81369 185147 81417 185175
rect 81445 185147 81479 185175
rect 81507 185147 81541 185175
rect 81569 185147 81603 185175
rect 81631 185147 81679 185175
rect 81369 185113 81679 185147
rect 81369 185085 81417 185113
rect 81445 185085 81479 185113
rect 81507 185085 81541 185113
rect 81569 185085 81603 185113
rect 81631 185085 81679 185113
rect 81369 185051 81679 185085
rect 81369 185023 81417 185051
rect 81445 185023 81479 185051
rect 81507 185023 81541 185051
rect 81569 185023 81603 185051
rect 81631 185023 81679 185051
rect 81369 184989 81679 185023
rect 81369 184961 81417 184989
rect 81445 184961 81479 184989
rect 81507 184961 81541 184989
rect 81569 184961 81603 184989
rect 81631 184961 81679 184989
rect 81369 176175 81679 184961
rect 81369 176147 81417 176175
rect 81445 176147 81479 176175
rect 81507 176147 81541 176175
rect 81569 176147 81603 176175
rect 81631 176147 81679 176175
rect 81369 176113 81679 176147
rect 81369 176085 81417 176113
rect 81445 176085 81479 176113
rect 81507 176085 81541 176113
rect 81569 176085 81603 176113
rect 81631 176085 81679 176113
rect 81369 176051 81679 176085
rect 81369 176023 81417 176051
rect 81445 176023 81479 176051
rect 81507 176023 81541 176051
rect 81569 176023 81603 176051
rect 81631 176023 81679 176051
rect 81369 175989 81679 176023
rect 81369 175961 81417 175989
rect 81445 175961 81479 175989
rect 81507 175961 81541 175989
rect 81569 175961 81603 175989
rect 81631 175961 81679 175989
rect 81369 167175 81679 175961
rect 94869 298606 95179 299134
rect 94869 298578 94917 298606
rect 94945 298578 94979 298606
rect 95007 298578 95041 298606
rect 95069 298578 95103 298606
rect 95131 298578 95179 298606
rect 94869 298544 95179 298578
rect 94869 298516 94917 298544
rect 94945 298516 94979 298544
rect 95007 298516 95041 298544
rect 95069 298516 95103 298544
rect 95131 298516 95179 298544
rect 94869 298482 95179 298516
rect 94869 298454 94917 298482
rect 94945 298454 94979 298482
rect 95007 298454 95041 298482
rect 95069 298454 95103 298482
rect 95131 298454 95179 298482
rect 94869 298420 95179 298454
rect 94869 298392 94917 298420
rect 94945 298392 94979 298420
rect 95007 298392 95041 298420
rect 95069 298392 95103 298420
rect 95131 298392 95179 298420
rect 94869 290175 95179 298392
rect 94869 290147 94917 290175
rect 94945 290147 94979 290175
rect 95007 290147 95041 290175
rect 95069 290147 95103 290175
rect 95131 290147 95179 290175
rect 94869 290113 95179 290147
rect 94869 290085 94917 290113
rect 94945 290085 94979 290113
rect 95007 290085 95041 290113
rect 95069 290085 95103 290113
rect 95131 290085 95179 290113
rect 94869 290051 95179 290085
rect 94869 290023 94917 290051
rect 94945 290023 94979 290051
rect 95007 290023 95041 290051
rect 95069 290023 95103 290051
rect 95131 290023 95179 290051
rect 94869 289989 95179 290023
rect 94869 289961 94917 289989
rect 94945 289961 94979 289989
rect 95007 289961 95041 289989
rect 95069 289961 95103 289989
rect 95131 289961 95179 289989
rect 94869 281175 95179 289961
rect 94869 281147 94917 281175
rect 94945 281147 94979 281175
rect 95007 281147 95041 281175
rect 95069 281147 95103 281175
rect 95131 281147 95179 281175
rect 94869 281113 95179 281147
rect 94869 281085 94917 281113
rect 94945 281085 94979 281113
rect 95007 281085 95041 281113
rect 95069 281085 95103 281113
rect 95131 281085 95179 281113
rect 94869 281051 95179 281085
rect 94869 281023 94917 281051
rect 94945 281023 94979 281051
rect 95007 281023 95041 281051
rect 95069 281023 95103 281051
rect 95131 281023 95179 281051
rect 94869 280989 95179 281023
rect 94869 280961 94917 280989
rect 94945 280961 94979 280989
rect 95007 280961 95041 280989
rect 95069 280961 95103 280989
rect 95131 280961 95179 280989
rect 94869 272175 95179 280961
rect 94869 272147 94917 272175
rect 94945 272147 94979 272175
rect 95007 272147 95041 272175
rect 95069 272147 95103 272175
rect 95131 272147 95179 272175
rect 94869 272113 95179 272147
rect 94869 272085 94917 272113
rect 94945 272085 94979 272113
rect 95007 272085 95041 272113
rect 95069 272085 95103 272113
rect 95131 272085 95179 272113
rect 94869 272051 95179 272085
rect 94869 272023 94917 272051
rect 94945 272023 94979 272051
rect 95007 272023 95041 272051
rect 95069 272023 95103 272051
rect 95131 272023 95179 272051
rect 94869 271989 95179 272023
rect 94869 271961 94917 271989
rect 94945 271961 94979 271989
rect 95007 271961 95041 271989
rect 95069 271961 95103 271989
rect 95131 271961 95179 271989
rect 94869 263175 95179 271961
rect 94869 263147 94917 263175
rect 94945 263147 94979 263175
rect 95007 263147 95041 263175
rect 95069 263147 95103 263175
rect 95131 263147 95179 263175
rect 94869 263113 95179 263147
rect 94869 263085 94917 263113
rect 94945 263085 94979 263113
rect 95007 263085 95041 263113
rect 95069 263085 95103 263113
rect 95131 263085 95179 263113
rect 94869 263051 95179 263085
rect 94869 263023 94917 263051
rect 94945 263023 94979 263051
rect 95007 263023 95041 263051
rect 95069 263023 95103 263051
rect 95131 263023 95179 263051
rect 94869 262989 95179 263023
rect 94869 262961 94917 262989
rect 94945 262961 94979 262989
rect 95007 262961 95041 262989
rect 95069 262961 95103 262989
rect 95131 262961 95179 262989
rect 94869 254175 95179 262961
rect 94869 254147 94917 254175
rect 94945 254147 94979 254175
rect 95007 254147 95041 254175
rect 95069 254147 95103 254175
rect 95131 254147 95179 254175
rect 94869 254113 95179 254147
rect 94869 254085 94917 254113
rect 94945 254085 94979 254113
rect 95007 254085 95041 254113
rect 95069 254085 95103 254113
rect 95131 254085 95179 254113
rect 94869 254051 95179 254085
rect 94869 254023 94917 254051
rect 94945 254023 94979 254051
rect 95007 254023 95041 254051
rect 95069 254023 95103 254051
rect 95131 254023 95179 254051
rect 94869 253989 95179 254023
rect 94869 253961 94917 253989
rect 94945 253961 94979 253989
rect 95007 253961 95041 253989
rect 95069 253961 95103 253989
rect 95131 253961 95179 253989
rect 94869 245175 95179 253961
rect 94869 245147 94917 245175
rect 94945 245147 94979 245175
rect 95007 245147 95041 245175
rect 95069 245147 95103 245175
rect 95131 245147 95179 245175
rect 94869 245113 95179 245147
rect 94869 245085 94917 245113
rect 94945 245085 94979 245113
rect 95007 245085 95041 245113
rect 95069 245085 95103 245113
rect 95131 245085 95179 245113
rect 94869 245051 95179 245085
rect 94869 245023 94917 245051
rect 94945 245023 94979 245051
rect 95007 245023 95041 245051
rect 95069 245023 95103 245051
rect 95131 245023 95179 245051
rect 94869 244989 95179 245023
rect 94869 244961 94917 244989
rect 94945 244961 94979 244989
rect 95007 244961 95041 244989
rect 95069 244961 95103 244989
rect 95131 244961 95179 244989
rect 94869 236175 95179 244961
rect 94869 236147 94917 236175
rect 94945 236147 94979 236175
rect 95007 236147 95041 236175
rect 95069 236147 95103 236175
rect 95131 236147 95179 236175
rect 94869 236113 95179 236147
rect 94869 236085 94917 236113
rect 94945 236085 94979 236113
rect 95007 236085 95041 236113
rect 95069 236085 95103 236113
rect 95131 236085 95179 236113
rect 94869 236051 95179 236085
rect 94869 236023 94917 236051
rect 94945 236023 94979 236051
rect 95007 236023 95041 236051
rect 95069 236023 95103 236051
rect 95131 236023 95179 236051
rect 94869 235989 95179 236023
rect 94869 235961 94917 235989
rect 94945 235961 94979 235989
rect 95007 235961 95041 235989
rect 95069 235961 95103 235989
rect 95131 235961 95179 235989
rect 94869 227175 95179 235961
rect 94869 227147 94917 227175
rect 94945 227147 94979 227175
rect 95007 227147 95041 227175
rect 95069 227147 95103 227175
rect 95131 227147 95179 227175
rect 94869 227113 95179 227147
rect 94869 227085 94917 227113
rect 94945 227085 94979 227113
rect 95007 227085 95041 227113
rect 95069 227085 95103 227113
rect 95131 227085 95179 227113
rect 94869 227051 95179 227085
rect 94869 227023 94917 227051
rect 94945 227023 94979 227051
rect 95007 227023 95041 227051
rect 95069 227023 95103 227051
rect 95131 227023 95179 227051
rect 94869 226989 95179 227023
rect 94869 226961 94917 226989
rect 94945 226961 94979 226989
rect 95007 226961 95041 226989
rect 95069 226961 95103 226989
rect 95131 226961 95179 226989
rect 94869 218175 95179 226961
rect 94869 218147 94917 218175
rect 94945 218147 94979 218175
rect 95007 218147 95041 218175
rect 95069 218147 95103 218175
rect 95131 218147 95179 218175
rect 94869 218113 95179 218147
rect 94869 218085 94917 218113
rect 94945 218085 94979 218113
rect 95007 218085 95041 218113
rect 95069 218085 95103 218113
rect 95131 218085 95179 218113
rect 94869 218051 95179 218085
rect 94869 218023 94917 218051
rect 94945 218023 94979 218051
rect 95007 218023 95041 218051
rect 95069 218023 95103 218051
rect 95131 218023 95179 218051
rect 94869 217989 95179 218023
rect 94869 217961 94917 217989
rect 94945 217961 94979 217989
rect 95007 217961 95041 217989
rect 95069 217961 95103 217989
rect 95131 217961 95179 217989
rect 94869 209175 95179 217961
rect 94869 209147 94917 209175
rect 94945 209147 94979 209175
rect 95007 209147 95041 209175
rect 95069 209147 95103 209175
rect 95131 209147 95179 209175
rect 94869 209113 95179 209147
rect 94869 209085 94917 209113
rect 94945 209085 94979 209113
rect 95007 209085 95041 209113
rect 95069 209085 95103 209113
rect 95131 209085 95179 209113
rect 94869 209051 95179 209085
rect 94869 209023 94917 209051
rect 94945 209023 94979 209051
rect 95007 209023 95041 209051
rect 95069 209023 95103 209051
rect 95131 209023 95179 209051
rect 94869 208989 95179 209023
rect 94869 208961 94917 208989
rect 94945 208961 94979 208989
rect 95007 208961 95041 208989
rect 95069 208961 95103 208989
rect 95131 208961 95179 208989
rect 94869 200175 95179 208961
rect 94869 200147 94917 200175
rect 94945 200147 94979 200175
rect 95007 200147 95041 200175
rect 95069 200147 95103 200175
rect 95131 200147 95179 200175
rect 94869 200113 95179 200147
rect 94869 200085 94917 200113
rect 94945 200085 94979 200113
rect 95007 200085 95041 200113
rect 95069 200085 95103 200113
rect 95131 200085 95179 200113
rect 94869 200051 95179 200085
rect 94869 200023 94917 200051
rect 94945 200023 94979 200051
rect 95007 200023 95041 200051
rect 95069 200023 95103 200051
rect 95131 200023 95179 200051
rect 94869 199989 95179 200023
rect 94869 199961 94917 199989
rect 94945 199961 94979 199989
rect 95007 199961 95041 199989
rect 95069 199961 95103 199989
rect 95131 199961 95179 199989
rect 94869 191175 95179 199961
rect 94869 191147 94917 191175
rect 94945 191147 94979 191175
rect 95007 191147 95041 191175
rect 95069 191147 95103 191175
rect 95131 191147 95179 191175
rect 94869 191113 95179 191147
rect 94869 191085 94917 191113
rect 94945 191085 94979 191113
rect 95007 191085 95041 191113
rect 95069 191085 95103 191113
rect 95131 191085 95179 191113
rect 94869 191051 95179 191085
rect 94869 191023 94917 191051
rect 94945 191023 94979 191051
rect 95007 191023 95041 191051
rect 95069 191023 95103 191051
rect 95131 191023 95179 191051
rect 94869 190989 95179 191023
rect 94869 190961 94917 190989
rect 94945 190961 94979 190989
rect 95007 190961 95041 190989
rect 95069 190961 95103 190989
rect 95131 190961 95179 190989
rect 94869 182175 95179 190961
rect 94869 182147 94917 182175
rect 94945 182147 94979 182175
rect 95007 182147 95041 182175
rect 95069 182147 95103 182175
rect 95131 182147 95179 182175
rect 94869 182113 95179 182147
rect 94869 182085 94917 182113
rect 94945 182085 94979 182113
rect 95007 182085 95041 182113
rect 95069 182085 95103 182113
rect 95131 182085 95179 182113
rect 94869 182051 95179 182085
rect 94869 182023 94917 182051
rect 94945 182023 94979 182051
rect 95007 182023 95041 182051
rect 95069 182023 95103 182051
rect 95131 182023 95179 182051
rect 94869 181989 95179 182023
rect 94869 181961 94917 181989
rect 94945 181961 94979 181989
rect 95007 181961 95041 181989
rect 95069 181961 95103 181989
rect 95131 181961 95179 181989
rect 85024 173175 85184 173192
rect 85024 173147 85059 173175
rect 85087 173147 85121 173175
rect 85149 173147 85184 173175
rect 85024 173113 85184 173147
rect 85024 173085 85059 173113
rect 85087 173085 85121 173113
rect 85149 173085 85184 173113
rect 85024 173051 85184 173085
rect 85024 173023 85059 173051
rect 85087 173023 85121 173051
rect 85149 173023 85184 173051
rect 85024 172989 85184 173023
rect 85024 172961 85059 172989
rect 85087 172961 85121 172989
rect 85149 172961 85184 172989
rect 85024 172944 85184 172961
rect 94869 173175 95179 181961
rect 94869 173147 94917 173175
rect 94945 173147 94979 173175
rect 95007 173147 95041 173175
rect 95069 173147 95103 173175
rect 95131 173147 95179 173175
rect 94869 173113 95179 173147
rect 94869 173085 94917 173113
rect 94945 173085 94979 173113
rect 95007 173085 95041 173113
rect 95069 173085 95103 173113
rect 95131 173085 95179 173113
rect 94869 173051 95179 173085
rect 94869 173023 94917 173051
rect 94945 173023 94979 173051
rect 95007 173023 95041 173051
rect 95069 173023 95103 173051
rect 95131 173023 95179 173051
rect 94869 172989 95179 173023
rect 94869 172961 94917 172989
rect 94945 172961 94979 172989
rect 95007 172961 95041 172989
rect 95069 172961 95103 172989
rect 95131 172961 95179 172989
rect 81369 167147 81417 167175
rect 81445 167147 81479 167175
rect 81507 167147 81541 167175
rect 81569 167147 81603 167175
rect 81631 167147 81679 167175
rect 81369 167113 81679 167147
rect 81369 167085 81417 167113
rect 81445 167085 81479 167113
rect 81507 167085 81541 167113
rect 81569 167085 81603 167113
rect 81631 167085 81679 167113
rect 81369 167051 81679 167085
rect 81369 167023 81417 167051
rect 81445 167023 81479 167051
rect 81507 167023 81541 167051
rect 81569 167023 81603 167051
rect 81631 167023 81679 167051
rect 81369 166989 81679 167023
rect 81369 166961 81417 166989
rect 81445 166961 81479 166989
rect 81507 166961 81541 166989
rect 81569 166961 81603 166989
rect 81631 166961 81679 166989
rect 81369 158175 81679 166961
rect 92704 167175 92864 167192
rect 92704 167147 92739 167175
rect 92767 167147 92801 167175
rect 92829 167147 92864 167175
rect 92704 167113 92864 167147
rect 92704 167085 92739 167113
rect 92767 167085 92801 167113
rect 92829 167085 92864 167113
rect 92704 167051 92864 167085
rect 92704 167023 92739 167051
rect 92767 167023 92801 167051
rect 92829 167023 92864 167051
rect 92704 166989 92864 167023
rect 92704 166961 92739 166989
rect 92767 166961 92801 166989
rect 92829 166961 92864 166989
rect 92704 166944 92864 166961
rect 85024 164175 85184 164192
rect 85024 164147 85059 164175
rect 85087 164147 85121 164175
rect 85149 164147 85184 164175
rect 85024 164113 85184 164147
rect 85024 164085 85059 164113
rect 85087 164085 85121 164113
rect 85149 164085 85184 164113
rect 85024 164051 85184 164085
rect 85024 164023 85059 164051
rect 85087 164023 85121 164051
rect 85149 164023 85184 164051
rect 85024 163989 85184 164023
rect 85024 163961 85059 163989
rect 85087 163961 85121 163989
rect 85149 163961 85184 163989
rect 85024 163944 85184 163961
rect 94869 164175 95179 172961
rect 94869 164147 94917 164175
rect 94945 164147 94979 164175
rect 95007 164147 95041 164175
rect 95069 164147 95103 164175
rect 95131 164147 95179 164175
rect 94869 164113 95179 164147
rect 94869 164085 94917 164113
rect 94945 164085 94979 164113
rect 95007 164085 95041 164113
rect 95069 164085 95103 164113
rect 95131 164085 95179 164113
rect 94869 164051 95179 164085
rect 94869 164023 94917 164051
rect 94945 164023 94979 164051
rect 95007 164023 95041 164051
rect 95069 164023 95103 164051
rect 95131 164023 95179 164051
rect 94869 163989 95179 164023
rect 94869 163961 94917 163989
rect 94945 163961 94979 163989
rect 95007 163961 95041 163989
rect 95069 163961 95103 163989
rect 95131 163961 95179 163989
rect 81369 158147 81417 158175
rect 81445 158147 81479 158175
rect 81507 158147 81541 158175
rect 81569 158147 81603 158175
rect 81631 158147 81679 158175
rect 81369 158113 81679 158147
rect 81369 158085 81417 158113
rect 81445 158085 81479 158113
rect 81507 158085 81541 158113
rect 81569 158085 81603 158113
rect 81631 158085 81679 158113
rect 81369 158051 81679 158085
rect 81369 158023 81417 158051
rect 81445 158023 81479 158051
rect 81507 158023 81541 158051
rect 81569 158023 81603 158051
rect 81631 158023 81679 158051
rect 81369 157989 81679 158023
rect 81369 157961 81417 157989
rect 81445 157961 81479 157989
rect 81507 157961 81541 157989
rect 81569 157961 81603 157989
rect 81631 157961 81679 157989
rect 81369 149175 81679 157961
rect 92704 158175 92864 158192
rect 92704 158147 92739 158175
rect 92767 158147 92801 158175
rect 92829 158147 92864 158175
rect 92704 158113 92864 158147
rect 92704 158085 92739 158113
rect 92767 158085 92801 158113
rect 92829 158085 92864 158113
rect 92704 158051 92864 158085
rect 92704 158023 92739 158051
rect 92767 158023 92801 158051
rect 92829 158023 92864 158051
rect 92704 157989 92864 158023
rect 92704 157961 92739 157989
rect 92767 157961 92801 157989
rect 92829 157961 92864 157989
rect 92704 157944 92864 157961
rect 85024 155175 85184 155192
rect 85024 155147 85059 155175
rect 85087 155147 85121 155175
rect 85149 155147 85184 155175
rect 85024 155113 85184 155147
rect 85024 155085 85059 155113
rect 85087 155085 85121 155113
rect 85149 155085 85184 155113
rect 85024 155051 85184 155085
rect 85024 155023 85059 155051
rect 85087 155023 85121 155051
rect 85149 155023 85184 155051
rect 85024 154989 85184 155023
rect 85024 154961 85059 154989
rect 85087 154961 85121 154989
rect 85149 154961 85184 154989
rect 85024 154944 85184 154961
rect 94869 155175 95179 163961
rect 94869 155147 94917 155175
rect 94945 155147 94979 155175
rect 95007 155147 95041 155175
rect 95069 155147 95103 155175
rect 95131 155147 95179 155175
rect 94869 155113 95179 155147
rect 94869 155085 94917 155113
rect 94945 155085 94979 155113
rect 95007 155085 95041 155113
rect 95069 155085 95103 155113
rect 95131 155085 95179 155113
rect 94869 155051 95179 155085
rect 94869 155023 94917 155051
rect 94945 155023 94979 155051
rect 95007 155023 95041 155051
rect 95069 155023 95103 155051
rect 95131 155023 95179 155051
rect 94869 154989 95179 155023
rect 94869 154961 94917 154989
rect 94945 154961 94979 154989
rect 95007 154961 95041 154989
rect 95069 154961 95103 154989
rect 95131 154961 95179 154989
rect 81369 149147 81417 149175
rect 81445 149147 81479 149175
rect 81507 149147 81541 149175
rect 81569 149147 81603 149175
rect 81631 149147 81679 149175
rect 81369 149113 81679 149147
rect 81369 149085 81417 149113
rect 81445 149085 81479 149113
rect 81507 149085 81541 149113
rect 81569 149085 81603 149113
rect 81631 149085 81679 149113
rect 81369 149051 81679 149085
rect 81369 149023 81417 149051
rect 81445 149023 81479 149051
rect 81507 149023 81541 149051
rect 81569 149023 81603 149051
rect 81631 149023 81679 149051
rect 81369 148989 81679 149023
rect 81369 148961 81417 148989
rect 81445 148961 81479 148989
rect 81507 148961 81541 148989
rect 81569 148961 81603 148989
rect 81631 148961 81679 148989
rect 81369 140175 81679 148961
rect 92704 149175 92864 149192
rect 92704 149147 92739 149175
rect 92767 149147 92801 149175
rect 92829 149147 92864 149175
rect 92704 149113 92864 149147
rect 92704 149085 92739 149113
rect 92767 149085 92801 149113
rect 92829 149085 92864 149113
rect 92704 149051 92864 149085
rect 92704 149023 92739 149051
rect 92767 149023 92801 149051
rect 92829 149023 92864 149051
rect 92704 148989 92864 149023
rect 92704 148961 92739 148989
rect 92767 148961 92801 148989
rect 92829 148961 92864 148989
rect 92704 148944 92864 148961
rect 85024 146175 85184 146192
rect 85024 146147 85059 146175
rect 85087 146147 85121 146175
rect 85149 146147 85184 146175
rect 85024 146113 85184 146147
rect 85024 146085 85059 146113
rect 85087 146085 85121 146113
rect 85149 146085 85184 146113
rect 85024 146051 85184 146085
rect 85024 146023 85059 146051
rect 85087 146023 85121 146051
rect 85149 146023 85184 146051
rect 85024 145989 85184 146023
rect 85024 145961 85059 145989
rect 85087 145961 85121 145989
rect 85149 145961 85184 145989
rect 85024 145944 85184 145961
rect 94869 146175 95179 154961
rect 94869 146147 94917 146175
rect 94945 146147 94979 146175
rect 95007 146147 95041 146175
rect 95069 146147 95103 146175
rect 95131 146147 95179 146175
rect 94869 146113 95179 146147
rect 94869 146085 94917 146113
rect 94945 146085 94979 146113
rect 95007 146085 95041 146113
rect 95069 146085 95103 146113
rect 95131 146085 95179 146113
rect 94869 146051 95179 146085
rect 94869 146023 94917 146051
rect 94945 146023 94979 146051
rect 95007 146023 95041 146051
rect 95069 146023 95103 146051
rect 95131 146023 95179 146051
rect 94869 145989 95179 146023
rect 94869 145961 94917 145989
rect 94945 145961 94979 145989
rect 95007 145961 95041 145989
rect 95069 145961 95103 145989
rect 95131 145961 95179 145989
rect 81369 140147 81417 140175
rect 81445 140147 81479 140175
rect 81507 140147 81541 140175
rect 81569 140147 81603 140175
rect 81631 140147 81679 140175
rect 81369 140113 81679 140147
rect 81369 140085 81417 140113
rect 81445 140085 81479 140113
rect 81507 140085 81541 140113
rect 81569 140085 81603 140113
rect 81631 140085 81679 140113
rect 81369 140051 81679 140085
rect 81369 140023 81417 140051
rect 81445 140023 81479 140051
rect 81507 140023 81541 140051
rect 81569 140023 81603 140051
rect 81631 140023 81679 140051
rect 81369 139989 81679 140023
rect 81369 139961 81417 139989
rect 81445 139961 81479 139989
rect 81507 139961 81541 139989
rect 81569 139961 81603 139989
rect 81631 139961 81679 139989
rect 81369 131175 81679 139961
rect 92704 140175 92864 140192
rect 92704 140147 92739 140175
rect 92767 140147 92801 140175
rect 92829 140147 92864 140175
rect 92704 140113 92864 140147
rect 92704 140085 92739 140113
rect 92767 140085 92801 140113
rect 92829 140085 92864 140113
rect 92704 140051 92864 140085
rect 92704 140023 92739 140051
rect 92767 140023 92801 140051
rect 92829 140023 92864 140051
rect 92704 139989 92864 140023
rect 92704 139961 92739 139989
rect 92767 139961 92801 139989
rect 92829 139961 92864 139989
rect 92704 139944 92864 139961
rect 85024 137175 85184 137192
rect 85024 137147 85059 137175
rect 85087 137147 85121 137175
rect 85149 137147 85184 137175
rect 85024 137113 85184 137147
rect 85024 137085 85059 137113
rect 85087 137085 85121 137113
rect 85149 137085 85184 137113
rect 85024 137051 85184 137085
rect 85024 137023 85059 137051
rect 85087 137023 85121 137051
rect 85149 137023 85184 137051
rect 85024 136989 85184 137023
rect 85024 136961 85059 136989
rect 85087 136961 85121 136989
rect 85149 136961 85184 136989
rect 85024 136944 85184 136961
rect 94869 137175 95179 145961
rect 94869 137147 94917 137175
rect 94945 137147 94979 137175
rect 95007 137147 95041 137175
rect 95069 137147 95103 137175
rect 95131 137147 95179 137175
rect 94869 137113 95179 137147
rect 94869 137085 94917 137113
rect 94945 137085 94979 137113
rect 95007 137085 95041 137113
rect 95069 137085 95103 137113
rect 95131 137085 95179 137113
rect 94869 137051 95179 137085
rect 94869 137023 94917 137051
rect 94945 137023 94979 137051
rect 95007 137023 95041 137051
rect 95069 137023 95103 137051
rect 95131 137023 95179 137051
rect 94869 136989 95179 137023
rect 94869 136961 94917 136989
rect 94945 136961 94979 136989
rect 95007 136961 95041 136989
rect 95069 136961 95103 136989
rect 95131 136961 95179 136989
rect 81369 131147 81417 131175
rect 81445 131147 81479 131175
rect 81507 131147 81541 131175
rect 81569 131147 81603 131175
rect 81631 131147 81679 131175
rect 81369 131113 81679 131147
rect 81369 131085 81417 131113
rect 81445 131085 81479 131113
rect 81507 131085 81541 131113
rect 81569 131085 81603 131113
rect 81631 131085 81679 131113
rect 81369 131051 81679 131085
rect 81369 131023 81417 131051
rect 81445 131023 81479 131051
rect 81507 131023 81541 131051
rect 81569 131023 81603 131051
rect 81631 131023 81679 131051
rect 81369 130989 81679 131023
rect 81369 130961 81417 130989
rect 81445 130961 81479 130989
rect 81507 130961 81541 130989
rect 81569 130961 81603 130989
rect 81631 130961 81679 130989
rect 81369 122175 81679 130961
rect 92704 131175 92864 131192
rect 92704 131147 92739 131175
rect 92767 131147 92801 131175
rect 92829 131147 92864 131175
rect 92704 131113 92864 131147
rect 92704 131085 92739 131113
rect 92767 131085 92801 131113
rect 92829 131085 92864 131113
rect 92704 131051 92864 131085
rect 92704 131023 92739 131051
rect 92767 131023 92801 131051
rect 92829 131023 92864 131051
rect 92704 130989 92864 131023
rect 92704 130961 92739 130989
rect 92767 130961 92801 130989
rect 92829 130961 92864 130989
rect 92704 130944 92864 130961
rect 85024 128175 85184 128192
rect 85024 128147 85059 128175
rect 85087 128147 85121 128175
rect 85149 128147 85184 128175
rect 85024 128113 85184 128147
rect 85024 128085 85059 128113
rect 85087 128085 85121 128113
rect 85149 128085 85184 128113
rect 85024 128051 85184 128085
rect 85024 128023 85059 128051
rect 85087 128023 85121 128051
rect 85149 128023 85184 128051
rect 85024 127989 85184 128023
rect 85024 127961 85059 127989
rect 85087 127961 85121 127989
rect 85149 127961 85184 127989
rect 85024 127944 85184 127961
rect 94869 128175 95179 136961
rect 94869 128147 94917 128175
rect 94945 128147 94979 128175
rect 95007 128147 95041 128175
rect 95069 128147 95103 128175
rect 95131 128147 95179 128175
rect 94869 128113 95179 128147
rect 94869 128085 94917 128113
rect 94945 128085 94979 128113
rect 95007 128085 95041 128113
rect 95069 128085 95103 128113
rect 95131 128085 95179 128113
rect 94869 128051 95179 128085
rect 94869 128023 94917 128051
rect 94945 128023 94979 128051
rect 95007 128023 95041 128051
rect 95069 128023 95103 128051
rect 95131 128023 95179 128051
rect 94869 127989 95179 128023
rect 94869 127961 94917 127989
rect 94945 127961 94979 127989
rect 95007 127961 95041 127989
rect 95069 127961 95103 127989
rect 95131 127961 95179 127989
rect 81369 122147 81417 122175
rect 81445 122147 81479 122175
rect 81507 122147 81541 122175
rect 81569 122147 81603 122175
rect 81631 122147 81679 122175
rect 81369 122113 81679 122147
rect 81369 122085 81417 122113
rect 81445 122085 81479 122113
rect 81507 122085 81541 122113
rect 81569 122085 81603 122113
rect 81631 122085 81679 122113
rect 81369 122051 81679 122085
rect 81369 122023 81417 122051
rect 81445 122023 81479 122051
rect 81507 122023 81541 122051
rect 81569 122023 81603 122051
rect 81631 122023 81679 122051
rect 81369 121989 81679 122023
rect 81369 121961 81417 121989
rect 81445 121961 81479 121989
rect 81507 121961 81541 121989
rect 81569 121961 81603 121989
rect 81631 121961 81679 121989
rect 81369 113175 81679 121961
rect 92704 122175 92864 122192
rect 92704 122147 92739 122175
rect 92767 122147 92801 122175
rect 92829 122147 92864 122175
rect 92704 122113 92864 122147
rect 92704 122085 92739 122113
rect 92767 122085 92801 122113
rect 92829 122085 92864 122113
rect 92704 122051 92864 122085
rect 92704 122023 92739 122051
rect 92767 122023 92801 122051
rect 92829 122023 92864 122051
rect 92704 121989 92864 122023
rect 92704 121961 92739 121989
rect 92767 121961 92801 121989
rect 92829 121961 92864 121989
rect 92704 121944 92864 121961
rect 85024 119175 85184 119192
rect 85024 119147 85059 119175
rect 85087 119147 85121 119175
rect 85149 119147 85184 119175
rect 85024 119113 85184 119147
rect 85024 119085 85059 119113
rect 85087 119085 85121 119113
rect 85149 119085 85184 119113
rect 85024 119051 85184 119085
rect 85024 119023 85059 119051
rect 85087 119023 85121 119051
rect 85149 119023 85184 119051
rect 85024 118989 85184 119023
rect 85024 118961 85059 118989
rect 85087 118961 85121 118989
rect 85149 118961 85184 118989
rect 85024 118944 85184 118961
rect 94869 119175 95179 127961
rect 94869 119147 94917 119175
rect 94945 119147 94979 119175
rect 95007 119147 95041 119175
rect 95069 119147 95103 119175
rect 95131 119147 95179 119175
rect 94869 119113 95179 119147
rect 94869 119085 94917 119113
rect 94945 119085 94979 119113
rect 95007 119085 95041 119113
rect 95069 119085 95103 119113
rect 95131 119085 95179 119113
rect 94869 119051 95179 119085
rect 94869 119023 94917 119051
rect 94945 119023 94979 119051
rect 95007 119023 95041 119051
rect 95069 119023 95103 119051
rect 95131 119023 95179 119051
rect 94869 118989 95179 119023
rect 94869 118961 94917 118989
rect 94945 118961 94979 118989
rect 95007 118961 95041 118989
rect 95069 118961 95103 118989
rect 95131 118961 95179 118989
rect 81369 113147 81417 113175
rect 81445 113147 81479 113175
rect 81507 113147 81541 113175
rect 81569 113147 81603 113175
rect 81631 113147 81679 113175
rect 81369 113113 81679 113147
rect 81369 113085 81417 113113
rect 81445 113085 81479 113113
rect 81507 113085 81541 113113
rect 81569 113085 81603 113113
rect 81631 113085 81679 113113
rect 81369 113051 81679 113085
rect 81369 113023 81417 113051
rect 81445 113023 81479 113051
rect 81507 113023 81541 113051
rect 81569 113023 81603 113051
rect 81631 113023 81679 113051
rect 81369 112989 81679 113023
rect 81369 112961 81417 112989
rect 81445 112961 81479 112989
rect 81507 112961 81541 112989
rect 81569 112961 81603 112989
rect 81631 112961 81679 112989
rect 81369 104175 81679 112961
rect 92704 113175 92864 113192
rect 92704 113147 92739 113175
rect 92767 113147 92801 113175
rect 92829 113147 92864 113175
rect 92704 113113 92864 113147
rect 92704 113085 92739 113113
rect 92767 113085 92801 113113
rect 92829 113085 92864 113113
rect 92704 113051 92864 113085
rect 92704 113023 92739 113051
rect 92767 113023 92801 113051
rect 92829 113023 92864 113051
rect 92704 112989 92864 113023
rect 92704 112961 92739 112989
rect 92767 112961 92801 112989
rect 92829 112961 92864 112989
rect 92704 112944 92864 112961
rect 85024 110175 85184 110192
rect 85024 110147 85059 110175
rect 85087 110147 85121 110175
rect 85149 110147 85184 110175
rect 85024 110113 85184 110147
rect 85024 110085 85059 110113
rect 85087 110085 85121 110113
rect 85149 110085 85184 110113
rect 85024 110051 85184 110085
rect 85024 110023 85059 110051
rect 85087 110023 85121 110051
rect 85149 110023 85184 110051
rect 85024 109989 85184 110023
rect 85024 109961 85059 109989
rect 85087 109961 85121 109989
rect 85149 109961 85184 109989
rect 85024 109944 85184 109961
rect 94869 110175 95179 118961
rect 94869 110147 94917 110175
rect 94945 110147 94979 110175
rect 95007 110147 95041 110175
rect 95069 110147 95103 110175
rect 95131 110147 95179 110175
rect 94869 110113 95179 110147
rect 94869 110085 94917 110113
rect 94945 110085 94979 110113
rect 95007 110085 95041 110113
rect 95069 110085 95103 110113
rect 95131 110085 95179 110113
rect 94869 110051 95179 110085
rect 94869 110023 94917 110051
rect 94945 110023 94979 110051
rect 95007 110023 95041 110051
rect 95069 110023 95103 110051
rect 95131 110023 95179 110051
rect 94869 109989 95179 110023
rect 94869 109961 94917 109989
rect 94945 109961 94979 109989
rect 95007 109961 95041 109989
rect 95069 109961 95103 109989
rect 95131 109961 95179 109989
rect 81369 104147 81417 104175
rect 81445 104147 81479 104175
rect 81507 104147 81541 104175
rect 81569 104147 81603 104175
rect 81631 104147 81679 104175
rect 81369 104113 81679 104147
rect 81369 104085 81417 104113
rect 81445 104085 81479 104113
rect 81507 104085 81541 104113
rect 81569 104085 81603 104113
rect 81631 104085 81679 104113
rect 81369 104051 81679 104085
rect 81369 104023 81417 104051
rect 81445 104023 81479 104051
rect 81507 104023 81541 104051
rect 81569 104023 81603 104051
rect 81631 104023 81679 104051
rect 81369 103989 81679 104023
rect 81369 103961 81417 103989
rect 81445 103961 81479 103989
rect 81507 103961 81541 103989
rect 81569 103961 81603 103989
rect 81631 103961 81679 103989
rect 81369 95175 81679 103961
rect 92704 104175 92864 104192
rect 92704 104147 92739 104175
rect 92767 104147 92801 104175
rect 92829 104147 92864 104175
rect 92704 104113 92864 104147
rect 92704 104085 92739 104113
rect 92767 104085 92801 104113
rect 92829 104085 92864 104113
rect 92704 104051 92864 104085
rect 92704 104023 92739 104051
rect 92767 104023 92801 104051
rect 92829 104023 92864 104051
rect 92704 103989 92864 104023
rect 92704 103961 92739 103989
rect 92767 103961 92801 103989
rect 92829 103961 92864 103989
rect 92704 103944 92864 103961
rect 85024 101175 85184 101192
rect 85024 101147 85059 101175
rect 85087 101147 85121 101175
rect 85149 101147 85184 101175
rect 85024 101113 85184 101147
rect 85024 101085 85059 101113
rect 85087 101085 85121 101113
rect 85149 101085 85184 101113
rect 85024 101051 85184 101085
rect 85024 101023 85059 101051
rect 85087 101023 85121 101051
rect 85149 101023 85184 101051
rect 85024 100989 85184 101023
rect 85024 100961 85059 100989
rect 85087 100961 85121 100989
rect 85149 100961 85184 100989
rect 85024 100944 85184 100961
rect 94869 101175 95179 109961
rect 94869 101147 94917 101175
rect 94945 101147 94979 101175
rect 95007 101147 95041 101175
rect 95069 101147 95103 101175
rect 95131 101147 95179 101175
rect 94869 101113 95179 101147
rect 94869 101085 94917 101113
rect 94945 101085 94979 101113
rect 95007 101085 95041 101113
rect 95069 101085 95103 101113
rect 95131 101085 95179 101113
rect 94869 101051 95179 101085
rect 94869 101023 94917 101051
rect 94945 101023 94979 101051
rect 95007 101023 95041 101051
rect 95069 101023 95103 101051
rect 95131 101023 95179 101051
rect 94869 100989 95179 101023
rect 94869 100961 94917 100989
rect 94945 100961 94979 100989
rect 95007 100961 95041 100989
rect 95069 100961 95103 100989
rect 95131 100961 95179 100989
rect 81369 95147 81417 95175
rect 81445 95147 81479 95175
rect 81507 95147 81541 95175
rect 81569 95147 81603 95175
rect 81631 95147 81679 95175
rect 81369 95113 81679 95147
rect 81369 95085 81417 95113
rect 81445 95085 81479 95113
rect 81507 95085 81541 95113
rect 81569 95085 81603 95113
rect 81631 95085 81679 95113
rect 81369 95051 81679 95085
rect 81369 95023 81417 95051
rect 81445 95023 81479 95051
rect 81507 95023 81541 95051
rect 81569 95023 81603 95051
rect 81631 95023 81679 95051
rect 81369 94989 81679 95023
rect 81369 94961 81417 94989
rect 81445 94961 81479 94989
rect 81507 94961 81541 94989
rect 81569 94961 81603 94989
rect 81631 94961 81679 94989
rect 81369 86175 81679 94961
rect 92704 95175 92864 95192
rect 92704 95147 92739 95175
rect 92767 95147 92801 95175
rect 92829 95147 92864 95175
rect 92704 95113 92864 95147
rect 92704 95085 92739 95113
rect 92767 95085 92801 95113
rect 92829 95085 92864 95113
rect 92704 95051 92864 95085
rect 92704 95023 92739 95051
rect 92767 95023 92801 95051
rect 92829 95023 92864 95051
rect 92704 94989 92864 95023
rect 92704 94961 92739 94989
rect 92767 94961 92801 94989
rect 92829 94961 92864 94989
rect 92704 94944 92864 94961
rect 85024 92175 85184 92192
rect 85024 92147 85059 92175
rect 85087 92147 85121 92175
rect 85149 92147 85184 92175
rect 85024 92113 85184 92147
rect 85024 92085 85059 92113
rect 85087 92085 85121 92113
rect 85149 92085 85184 92113
rect 85024 92051 85184 92085
rect 85024 92023 85059 92051
rect 85087 92023 85121 92051
rect 85149 92023 85184 92051
rect 85024 91989 85184 92023
rect 85024 91961 85059 91989
rect 85087 91961 85121 91989
rect 85149 91961 85184 91989
rect 85024 91944 85184 91961
rect 94869 92175 95179 100961
rect 94869 92147 94917 92175
rect 94945 92147 94979 92175
rect 95007 92147 95041 92175
rect 95069 92147 95103 92175
rect 95131 92147 95179 92175
rect 94869 92113 95179 92147
rect 94869 92085 94917 92113
rect 94945 92085 94979 92113
rect 95007 92085 95041 92113
rect 95069 92085 95103 92113
rect 95131 92085 95179 92113
rect 94869 92051 95179 92085
rect 94869 92023 94917 92051
rect 94945 92023 94979 92051
rect 95007 92023 95041 92051
rect 95069 92023 95103 92051
rect 95131 92023 95179 92051
rect 94869 91989 95179 92023
rect 94869 91961 94917 91989
rect 94945 91961 94979 91989
rect 95007 91961 95041 91989
rect 95069 91961 95103 91989
rect 95131 91961 95179 91989
rect 81369 86147 81417 86175
rect 81445 86147 81479 86175
rect 81507 86147 81541 86175
rect 81569 86147 81603 86175
rect 81631 86147 81679 86175
rect 81369 86113 81679 86147
rect 81369 86085 81417 86113
rect 81445 86085 81479 86113
rect 81507 86085 81541 86113
rect 81569 86085 81603 86113
rect 81631 86085 81679 86113
rect 81369 86051 81679 86085
rect 81369 86023 81417 86051
rect 81445 86023 81479 86051
rect 81507 86023 81541 86051
rect 81569 86023 81603 86051
rect 81631 86023 81679 86051
rect 81369 85989 81679 86023
rect 81369 85961 81417 85989
rect 81445 85961 81479 85989
rect 81507 85961 81541 85989
rect 81569 85961 81603 85989
rect 81631 85961 81679 85989
rect 81369 77175 81679 85961
rect 92704 86175 92864 86192
rect 92704 86147 92739 86175
rect 92767 86147 92801 86175
rect 92829 86147 92864 86175
rect 92704 86113 92864 86147
rect 92704 86085 92739 86113
rect 92767 86085 92801 86113
rect 92829 86085 92864 86113
rect 92704 86051 92864 86085
rect 92704 86023 92739 86051
rect 92767 86023 92801 86051
rect 92829 86023 92864 86051
rect 92704 85989 92864 86023
rect 92704 85961 92739 85989
rect 92767 85961 92801 85989
rect 92829 85961 92864 85989
rect 92704 85944 92864 85961
rect 85024 83175 85184 83192
rect 85024 83147 85059 83175
rect 85087 83147 85121 83175
rect 85149 83147 85184 83175
rect 85024 83113 85184 83147
rect 85024 83085 85059 83113
rect 85087 83085 85121 83113
rect 85149 83085 85184 83113
rect 85024 83051 85184 83085
rect 85024 83023 85059 83051
rect 85087 83023 85121 83051
rect 85149 83023 85184 83051
rect 85024 82989 85184 83023
rect 85024 82961 85059 82989
rect 85087 82961 85121 82989
rect 85149 82961 85184 82989
rect 85024 82944 85184 82961
rect 94869 83175 95179 91961
rect 94869 83147 94917 83175
rect 94945 83147 94979 83175
rect 95007 83147 95041 83175
rect 95069 83147 95103 83175
rect 95131 83147 95179 83175
rect 94869 83113 95179 83147
rect 94869 83085 94917 83113
rect 94945 83085 94979 83113
rect 95007 83085 95041 83113
rect 95069 83085 95103 83113
rect 95131 83085 95179 83113
rect 94869 83051 95179 83085
rect 94869 83023 94917 83051
rect 94945 83023 94979 83051
rect 95007 83023 95041 83051
rect 95069 83023 95103 83051
rect 95131 83023 95179 83051
rect 94869 82989 95179 83023
rect 94869 82961 94917 82989
rect 94945 82961 94979 82989
rect 95007 82961 95041 82989
rect 95069 82961 95103 82989
rect 95131 82961 95179 82989
rect 81369 77147 81417 77175
rect 81445 77147 81479 77175
rect 81507 77147 81541 77175
rect 81569 77147 81603 77175
rect 81631 77147 81679 77175
rect 81369 77113 81679 77147
rect 81369 77085 81417 77113
rect 81445 77085 81479 77113
rect 81507 77085 81541 77113
rect 81569 77085 81603 77113
rect 81631 77085 81679 77113
rect 81369 77051 81679 77085
rect 81369 77023 81417 77051
rect 81445 77023 81479 77051
rect 81507 77023 81541 77051
rect 81569 77023 81603 77051
rect 81631 77023 81679 77051
rect 81369 76989 81679 77023
rect 81369 76961 81417 76989
rect 81445 76961 81479 76989
rect 81507 76961 81541 76989
rect 81569 76961 81603 76989
rect 81631 76961 81679 76989
rect 81369 68175 81679 76961
rect 92704 77175 92864 77192
rect 92704 77147 92739 77175
rect 92767 77147 92801 77175
rect 92829 77147 92864 77175
rect 92704 77113 92864 77147
rect 92704 77085 92739 77113
rect 92767 77085 92801 77113
rect 92829 77085 92864 77113
rect 92704 77051 92864 77085
rect 92704 77023 92739 77051
rect 92767 77023 92801 77051
rect 92829 77023 92864 77051
rect 92704 76989 92864 77023
rect 92704 76961 92739 76989
rect 92767 76961 92801 76989
rect 92829 76961 92864 76989
rect 92704 76944 92864 76961
rect 85024 74175 85184 74192
rect 85024 74147 85059 74175
rect 85087 74147 85121 74175
rect 85149 74147 85184 74175
rect 85024 74113 85184 74147
rect 85024 74085 85059 74113
rect 85087 74085 85121 74113
rect 85149 74085 85184 74113
rect 85024 74051 85184 74085
rect 85024 74023 85059 74051
rect 85087 74023 85121 74051
rect 85149 74023 85184 74051
rect 85024 73989 85184 74023
rect 85024 73961 85059 73989
rect 85087 73961 85121 73989
rect 85149 73961 85184 73989
rect 85024 73944 85184 73961
rect 94869 74175 95179 82961
rect 94869 74147 94917 74175
rect 94945 74147 94979 74175
rect 95007 74147 95041 74175
rect 95069 74147 95103 74175
rect 95131 74147 95179 74175
rect 94869 74113 95179 74147
rect 94869 74085 94917 74113
rect 94945 74085 94979 74113
rect 95007 74085 95041 74113
rect 95069 74085 95103 74113
rect 95131 74085 95179 74113
rect 94869 74051 95179 74085
rect 94869 74023 94917 74051
rect 94945 74023 94979 74051
rect 95007 74023 95041 74051
rect 95069 74023 95103 74051
rect 95131 74023 95179 74051
rect 94869 73989 95179 74023
rect 94869 73961 94917 73989
rect 94945 73961 94979 73989
rect 95007 73961 95041 73989
rect 95069 73961 95103 73989
rect 95131 73961 95179 73989
rect 81369 68147 81417 68175
rect 81445 68147 81479 68175
rect 81507 68147 81541 68175
rect 81569 68147 81603 68175
rect 81631 68147 81679 68175
rect 81369 68113 81679 68147
rect 81369 68085 81417 68113
rect 81445 68085 81479 68113
rect 81507 68085 81541 68113
rect 81569 68085 81603 68113
rect 81631 68085 81679 68113
rect 81369 68051 81679 68085
rect 81369 68023 81417 68051
rect 81445 68023 81479 68051
rect 81507 68023 81541 68051
rect 81569 68023 81603 68051
rect 81631 68023 81679 68051
rect 81369 67989 81679 68023
rect 81369 67961 81417 67989
rect 81445 67961 81479 67989
rect 81507 67961 81541 67989
rect 81569 67961 81603 67989
rect 81631 67961 81679 67989
rect 81369 59175 81679 67961
rect 92704 68175 92864 68192
rect 92704 68147 92739 68175
rect 92767 68147 92801 68175
rect 92829 68147 92864 68175
rect 92704 68113 92864 68147
rect 92704 68085 92739 68113
rect 92767 68085 92801 68113
rect 92829 68085 92864 68113
rect 92704 68051 92864 68085
rect 92704 68023 92739 68051
rect 92767 68023 92801 68051
rect 92829 68023 92864 68051
rect 92704 67989 92864 68023
rect 92704 67961 92739 67989
rect 92767 67961 92801 67989
rect 92829 67961 92864 67989
rect 92704 67944 92864 67961
rect 85024 65175 85184 65192
rect 85024 65147 85059 65175
rect 85087 65147 85121 65175
rect 85149 65147 85184 65175
rect 85024 65113 85184 65147
rect 85024 65085 85059 65113
rect 85087 65085 85121 65113
rect 85149 65085 85184 65113
rect 85024 65051 85184 65085
rect 85024 65023 85059 65051
rect 85087 65023 85121 65051
rect 85149 65023 85184 65051
rect 85024 64989 85184 65023
rect 85024 64961 85059 64989
rect 85087 64961 85121 64989
rect 85149 64961 85184 64989
rect 85024 64944 85184 64961
rect 94869 65175 95179 73961
rect 94869 65147 94917 65175
rect 94945 65147 94979 65175
rect 95007 65147 95041 65175
rect 95069 65147 95103 65175
rect 95131 65147 95179 65175
rect 94869 65113 95179 65147
rect 94869 65085 94917 65113
rect 94945 65085 94979 65113
rect 95007 65085 95041 65113
rect 95069 65085 95103 65113
rect 95131 65085 95179 65113
rect 94869 65051 95179 65085
rect 94869 65023 94917 65051
rect 94945 65023 94979 65051
rect 95007 65023 95041 65051
rect 95069 65023 95103 65051
rect 95131 65023 95179 65051
rect 94869 64989 95179 65023
rect 94869 64961 94917 64989
rect 94945 64961 94979 64989
rect 95007 64961 95041 64989
rect 95069 64961 95103 64989
rect 95131 64961 95179 64989
rect 81369 59147 81417 59175
rect 81445 59147 81479 59175
rect 81507 59147 81541 59175
rect 81569 59147 81603 59175
rect 81631 59147 81679 59175
rect 81369 59113 81679 59147
rect 81369 59085 81417 59113
rect 81445 59085 81479 59113
rect 81507 59085 81541 59113
rect 81569 59085 81603 59113
rect 81631 59085 81679 59113
rect 81369 59051 81679 59085
rect 81369 59023 81417 59051
rect 81445 59023 81479 59051
rect 81507 59023 81541 59051
rect 81569 59023 81603 59051
rect 81631 59023 81679 59051
rect 81369 58989 81679 59023
rect 81369 58961 81417 58989
rect 81445 58961 81479 58989
rect 81507 58961 81541 58989
rect 81569 58961 81603 58989
rect 81631 58961 81679 58989
rect 81369 50175 81679 58961
rect 92704 59175 92864 59192
rect 92704 59147 92739 59175
rect 92767 59147 92801 59175
rect 92829 59147 92864 59175
rect 92704 59113 92864 59147
rect 92704 59085 92739 59113
rect 92767 59085 92801 59113
rect 92829 59085 92864 59113
rect 92704 59051 92864 59085
rect 92704 59023 92739 59051
rect 92767 59023 92801 59051
rect 92829 59023 92864 59051
rect 92704 58989 92864 59023
rect 92704 58961 92739 58989
rect 92767 58961 92801 58989
rect 92829 58961 92864 58989
rect 92704 58944 92864 58961
rect 85024 56175 85184 56192
rect 85024 56147 85059 56175
rect 85087 56147 85121 56175
rect 85149 56147 85184 56175
rect 85024 56113 85184 56147
rect 85024 56085 85059 56113
rect 85087 56085 85121 56113
rect 85149 56085 85184 56113
rect 85024 56051 85184 56085
rect 85024 56023 85059 56051
rect 85087 56023 85121 56051
rect 85149 56023 85184 56051
rect 85024 55989 85184 56023
rect 85024 55961 85059 55989
rect 85087 55961 85121 55989
rect 85149 55961 85184 55989
rect 85024 55944 85184 55961
rect 94869 56175 95179 64961
rect 94869 56147 94917 56175
rect 94945 56147 94979 56175
rect 95007 56147 95041 56175
rect 95069 56147 95103 56175
rect 95131 56147 95179 56175
rect 94869 56113 95179 56147
rect 94869 56085 94917 56113
rect 94945 56085 94979 56113
rect 95007 56085 95041 56113
rect 95069 56085 95103 56113
rect 95131 56085 95179 56113
rect 94869 56051 95179 56085
rect 94869 56023 94917 56051
rect 94945 56023 94979 56051
rect 95007 56023 95041 56051
rect 95069 56023 95103 56051
rect 95131 56023 95179 56051
rect 94869 55989 95179 56023
rect 94869 55961 94917 55989
rect 94945 55961 94979 55989
rect 95007 55961 95041 55989
rect 95069 55961 95103 55989
rect 95131 55961 95179 55989
rect 81369 50147 81417 50175
rect 81445 50147 81479 50175
rect 81507 50147 81541 50175
rect 81569 50147 81603 50175
rect 81631 50147 81679 50175
rect 81369 50113 81679 50147
rect 81369 50085 81417 50113
rect 81445 50085 81479 50113
rect 81507 50085 81541 50113
rect 81569 50085 81603 50113
rect 81631 50085 81679 50113
rect 81369 50051 81679 50085
rect 81369 50023 81417 50051
rect 81445 50023 81479 50051
rect 81507 50023 81541 50051
rect 81569 50023 81603 50051
rect 81631 50023 81679 50051
rect 81369 49989 81679 50023
rect 81369 49961 81417 49989
rect 81445 49961 81479 49989
rect 81507 49961 81541 49989
rect 81569 49961 81603 49989
rect 81631 49961 81679 49989
rect 81369 41175 81679 49961
rect 92704 50175 92864 50192
rect 92704 50147 92739 50175
rect 92767 50147 92801 50175
rect 92829 50147 92864 50175
rect 92704 50113 92864 50147
rect 92704 50085 92739 50113
rect 92767 50085 92801 50113
rect 92829 50085 92864 50113
rect 92704 50051 92864 50085
rect 92704 50023 92739 50051
rect 92767 50023 92801 50051
rect 92829 50023 92864 50051
rect 92704 49989 92864 50023
rect 92704 49961 92739 49989
rect 92767 49961 92801 49989
rect 92829 49961 92864 49989
rect 92704 49944 92864 49961
rect 85024 47175 85184 47192
rect 85024 47147 85059 47175
rect 85087 47147 85121 47175
rect 85149 47147 85184 47175
rect 85024 47113 85184 47147
rect 85024 47085 85059 47113
rect 85087 47085 85121 47113
rect 85149 47085 85184 47113
rect 85024 47051 85184 47085
rect 85024 47023 85059 47051
rect 85087 47023 85121 47051
rect 85149 47023 85184 47051
rect 85024 46989 85184 47023
rect 85024 46961 85059 46989
rect 85087 46961 85121 46989
rect 85149 46961 85184 46989
rect 85024 46944 85184 46961
rect 94869 47175 95179 55961
rect 94869 47147 94917 47175
rect 94945 47147 94979 47175
rect 95007 47147 95041 47175
rect 95069 47147 95103 47175
rect 95131 47147 95179 47175
rect 94869 47113 95179 47147
rect 94869 47085 94917 47113
rect 94945 47085 94979 47113
rect 95007 47085 95041 47113
rect 95069 47085 95103 47113
rect 95131 47085 95179 47113
rect 94869 47051 95179 47085
rect 94869 47023 94917 47051
rect 94945 47023 94979 47051
rect 95007 47023 95041 47051
rect 95069 47023 95103 47051
rect 95131 47023 95179 47051
rect 94869 46989 95179 47023
rect 94869 46961 94917 46989
rect 94945 46961 94979 46989
rect 95007 46961 95041 46989
rect 95069 46961 95103 46989
rect 95131 46961 95179 46989
rect 81369 41147 81417 41175
rect 81445 41147 81479 41175
rect 81507 41147 81541 41175
rect 81569 41147 81603 41175
rect 81631 41147 81679 41175
rect 81369 41113 81679 41147
rect 81369 41085 81417 41113
rect 81445 41085 81479 41113
rect 81507 41085 81541 41113
rect 81569 41085 81603 41113
rect 81631 41085 81679 41113
rect 81369 41051 81679 41085
rect 81369 41023 81417 41051
rect 81445 41023 81479 41051
rect 81507 41023 81541 41051
rect 81569 41023 81603 41051
rect 81631 41023 81679 41051
rect 81369 40989 81679 41023
rect 81369 40961 81417 40989
rect 81445 40961 81479 40989
rect 81507 40961 81541 40989
rect 81569 40961 81603 40989
rect 81631 40961 81679 40989
rect 81369 32175 81679 40961
rect 92704 41175 92864 41192
rect 92704 41147 92739 41175
rect 92767 41147 92801 41175
rect 92829 41147 92864 41175
rect 92704 41113 92864 41147
rect 92704 41085 92739 41113
rect 92767 41085 92801 41113
rect 92829 41085 92864 41113
rect 92704 41051 92864 41085
rect 92704 41023 92739 41051
rect 92767 41023 92801 41051
rect 92829 41023 92864 41051
rect 92704 40989 92864 41023
rect 92704 40961 92739 40989
rect 92767 40961 92801 40989
rect 92829 40961 92864 40989
rect 92704 40944 92864 40961
rect 85024 38175 85184 38192
rect 85024 38147 85059 38175
rect 85087 38147 85121 38175
rect 85149 38147 85184 38175
rect 85024 38113 85184 38147
rect 85024 38085 85059 38113
rect 85087 38085 85121 38113
rect 85149 38085 85184 38113
rect 85024 38051 85184 38085
rect 85024 38023 85059 38051
rect 85087 38023 85121 38051
rect 85149 38023 85184 38051
rect 85024 37989 85184 38023
rect 85024 37961 85059 37989
rect 85087 37961 85121 37989
rect 85149 37961 85184 37989
rect 85024 37944 85184 37961
rect 94869 38175 95179 46961
rect 94869 38147 94917 38175
rect 94945 38147 94979 38175
rect 95007 38147 95041 38175
rect 95069 38147 95103 38175
rect 95131 38147 95179 38175
rect 94869 38113 95179 38147
rect 94869 38085 94917 38113
rect 94945 38085 94979 38113
rect 95007 38085 95041 38113
rect 95069 38085 95103 38113
rect 95131 38085 95179 38113
rect 94869 38051 95179 38085
rect 94869 38023 94917 38051
rect 94945 38023 94979 38051
rect 95007 38023 95041 38051
rect 95069 38023 95103 38051
rect 95131 38023 95179 38051
rect 94869 37989 95179 38023
rect 94869 37961 94917 37989
rect 94945 37961 94979 37989
rect 95007 37961 95041 37989
rect 95069 37961 95103 37989
rect 95131 37961 95179 37989
rect 81369 32147 81417 32175
rect 81445 32147 81479 32175
rect 81507 32147 81541 32175
rect 81569 32147 81603 32175
rect 81631 32147 81679 32175
rect 81369 32113 81679 32147
rect 81369 32085 81417 32113
rect 81445 32085 81479 32113
rect 81507 32085 81541 32113
rect 81569 32085 81603 32113
rect 81631 32085 81679 32113
rect 81369 32051 81679 32085
rect 81369 32023 81417 32051
rect 81445 32023 81479 32051
rect 81507 32023 81541 32051
rect 81569 32023 81603 32051
rect 81631 32023 81679 32051
rect 81369 31989 81679 32023
rect 81369 31961 81417 31989
rect 81445 31961 81479 31989
rect 81507 31961 81541 31989
rect 81569 31961 81603 31989
rect 81631 31961 81679 31989
rect 81369 23175 81679 31961
rect 92704 32175 92864 32192
rect 92704 32147 92739 32175
rect 92767 32147 92801 32175
rect 92829 32147 92864 32175
rect 92704 32113 92864 32147
rect 92704 32085 92739 32113
rect 92767 32085 92801 32113
rect 92829 32085 92864 32113
rect 92704 32051 92864 32085
rect 92704 32023 92739 32051
rect 92767 32023 92801 32051
rect 92829 32023 92864 32051
rect 92704 31989 92864 32023
rect 92704 31961 92739 31989
rect 92767 31961 92801 31989
rect 92829 31961 92864 31989
rect 92704 31944 92864 31961
rect 85024 29175 85184 29192
rect 85024 29147 85059 29175
rect 85087 29147 85121 29175
rect 85149 29147 85184 29175
rect 85024 29113 85184 29147
rect 85024 29085 85059 29113
rect 85087 29085 85121 29113
rect 85149 29085 85184 29113
rect 85024 29051 85184 29085
rect 85024 29023 85059 29051
rect 85087 29023 85121 29051
rect 85149 29023 85184 29051
rect 85024 28989 85184 29023
rect 85024 28961 85059 28989
rect 85087 28961 85121 28989
rect 85149 28961 85184 28989
rect 85024 28944 85184 28961
rect 94869 29175 95179 37961
rect 94869 29147 94917 29175
rect 94945 29147 94979 29175
rect 95007 29147 95041 29175
rect 95069 29147 95103 29175
rect 95131 29147 95179 29175
rect 94869 29113 95179 29147
rect 94869 29085 94917 29113
rect 94945 29085 94979 29113
rect 95007 29085 95041 29113
rect 95069 29085 95103 29113
rect 95131 29085 95179 29113
rect 94869 29051 95179 29085
rect 94869 29023 94917 29051
rect 94945 29023 94979 29051
rect 95007 29023 95041 29051
rect 95069 29023 95103 29051
rect 95131 29023 95179 29051
rect 94869 28989 95179 29023
rect 94869 28961 94917 28989
rect 94945 28961 94979 28989
rect 95007 28961 95041 28989
rect 95069 28961 95103 28989
rect 95131 28961 95179 28989
rect 81369 23147 81417 23175
rect 81445 23147 81479 23175
rect 81507 23147 81541 23175
rect 81569 23147 81603 23175
rect 81631 23147 81679 23175
rect 81369 23113 81679 23147
rect 81369 23085 81417 23113
rect 81445 23085 81479 23113
rect 81507 23085 81541 23113
rect 81569 23085 81603 23113
rect 81631 23085 81679 23113
rect 81369 23051 81679 23085
rect 81369 23023 81417 23051
rect 81445 23023 81479 23051
rect 81507 23023 81541 23051
rect 81569 23023 81603 23051
rect 81631 23023 81679 23051
rect 81369 22989 81679 23023
rect 81369 22961 81417 22989
rect 81445 22961 81479 22989
rect 81507 22961 81541 22989
rect 81569 22961 81603 22989
rect 81631 22961 81679 22989
rect 81369 14175 81679 22961
rect 92704 23175 92864 23192
rect 92704 23147 92739 23175
rect 92767 23147 92801 23175
rect 92829 23147 92864 23175
rect 92704 23113 92864 23147
rect 92704 23085 92739 23113
rect 92767 23085 92801 23113
rect 92829 23085 92864 23113
rect 92704 23051 92864 23085
rect 92704 23023 92739 23051
rect 92767 23023 92801 23051
rect 92829 23023 92864 23051
rect 92704 22989 92864 23023
rect 92704 22961 92739 22989
rect 92767 22961 92801 22989
rect 92829 22961 92864 22989
rect 92704 22944 92864 22961
rect 85024 20175 85184 20192
rect 85024 20147 85059 20175
rect 85087 20147 85121 20175
rect 85149 20147 85184 20175
rect 85024 20113 85184 20147
rect 85024 20085 85059 20113
rect 85087 20085 85121 20113
rect 85149 20085 85184 20113
rect 85024 20051 85184 20085
rect 85024 20023 85059 20051
rect 85087 20023 85121 20051
rect 85149 20023 85184 20051
rect 85024 19989 85184 20023
rect 85024 19961 85059 19989
rect 85087 19961 85121 19989
rect 85149 19961 85184 19989
rect 85024 19944 85184 19961
rect 94869 20175 95179 28961
rect 94869 20147 94917 20175
rect 94945 20147 94979 20175
rect 95007 20147 95041 20175
rect 95069 20147 95103 20175
rect 95131 20147 95179 20175
rect 94869 20113 95179 20147
rect 94869 20085 94917 20113
rect 94945 20085 94979 20113
rect 95007 20085 95041 20113
rect 95069 20085 95103 20113
rect 95131 20085 95179 20113
rect 94869 20051 95179 20085
rect 94869 20023 94917 20051
rect 94945 20023 94979 20051
rect 95007 20023 95041 20051
rect 95069 20023 95103 20051
rect 95131 20023 95179 20051
rect 94869 19989 95179 20023
rect 94869 19961 94917 19989
rect 94945 19961 94979 19989
rect 95007 19961 95041 19989
rect 95069 19961 95103 19989
rect 95131 19961 95179 19989
rect 81369 14147 81417 14175
rect 81445 14147 81479 14175
rect 81507 14147 81541 14175
rect 81569 14147 81603 14175
rect 81631 14147 81679 14175
rect 81369 14113 81679 14147
rect 81369 14085 81417 14113
rect 81445 14085 81479 14113
rect 81507 14085 81541 14113
rect 81569 14085 81603 14113
rect 81631 14085 81679 14113
rect 81369 14051 81679 14085
rect 81369 14023 81417 14051
rect 81445 14023 81479 14051
rect 81507 14023 81541 14051
rect 81569 14023 81603 14051
rect 81631 14023 81679 14051
rect 81369 13989 81679 14023
rect 81369 13961 81417 13989
rect 81445 13961 81479 13989
rect 81507 13961 81541 13989
rect 81569 13961 81603 13989
rect 81631 13961 81679 13989
rect 81369 5175 81679 13961
rect 92704 14175 92864 14192
rect 92704 14147 92739 14175
rect 92767 14147 92801 14175
rect 92829 14147 92864 14175
rect 92704 14113 92864 14147
rect 92704 14085 92739 14113
rect 92767 14085 92801 14113
rect 92829 14085 92864 14113
rect 92704 14051 92864 14085
rect 92704 14023 92739 14051
rect 92767 14023 92801 14051
rect 92829 14023 92864 14051
rect 92704 13989 92864 14023
rect 92704 13961 92739 13989
rect 92767 13961 92801 13989
rect 92829 13961 92864 13989
rect 92704 13944 92864 13961
rect 85024 11175 85184 11192
rect 85024 11147 85059 11175
rect 85087 11147 85121 11175
rect 85149 11147 85184 11175
rect 85024 11113 85184 11147
rect 85024 11085 85059 11113
rect 85087 11085 85121 11113
rect 85149 11085 85184 11113
rect 85024 11051 85184 11085
rect 85024 11023 85059 11051
rect 85087 11023 85121 11051
rect 85149 11023 85184 11051
rect 85024 10989 85184 11023
rect 85024 10961 85059 10989
rect 85087 10961 85121 10989
rect 85149 10961 85184 10989
rect 85024 10944 85184 10961
rect 94869 11175 95179 19961
rect 94869 11147 94917 11175
rect 94945 11147 94979 11175
rect 95007 11147 95041 11175
rect 95069 11147 95103 11175
rect 95131 11147 95179 11175
rect 94869 11113 95179 11147
rect 94869 11085 94917 11113
rect 94945 11085 94979 11113
rect 95007 11085 95041 11113
rect 95069 11085 95103 11113
rect 95131 11085 95179 11113
rect 94869 11051 95179 11085
rect 94869 11023 94917 11051
rect 94945 11023 94979 11051
rect 95007 11023 95041 11051
rect 95069 11023 95103 11051
rect 95131 11023 95179 11051
rect 94869 10989 95179 11023
rect 94869 10961 94917 10989
rect 94945 10961 94979 10989
rect 95007 10961 95041 10989
rect 95069 10961 95103 10989
rect 95131 10961 95179 10989
rect 81369 5147 81417 5175
rect 81445 5147 81479 5175
rect 81507 5147 81541 5175
rect 81569 5147 81603 5175
rect 81631 5147 81679 5175
rect 81369 5113 81679 5147
rect 81369 5085 81417 5113
rect 81445 5085 81479 5113
rect 81507 5085 81541 5113
rect 81569 5085 81603 5113
rect 81631 5085 81679 5113
rect 81369 5051 81679 5085
rect 81369 5023 81417 5051
rect 81445 5023 81479 5051
rect 81507 5023 81541 5051
rect 81569 5023 81603 5051
rect 81631 5023 81679 5051
rect 81369 4989 81679 5023
rect 81369 4961 81417 4989
rect 81445 4961 81479 4989
rect 81507 4961 81541 4989
rect 81569 4961 81603 4989
rect 81631 4961 81679 4989
rect 81369 -560 81679 4961
rect 92704 5175 92864 5192
rect 92704 5147 92739 5175
rect 92767 5147 92801 5175
rect 92829 5147 92864 5175
rect 92704 5113 92864 5147
rect 92704 5085 92739 5113
rect 92767 5085 92801 5113
rect 92829 5085 92864 5113
rect 92704 5051 92864 5085
rect 92704 5023 92739 5051
rect 92767 5023 92801 5051
rect 92829 5023 92864 5051
rect 92704 4989 92864 5023
rect 92704 4961 92739 4989
rect 92767 4961 92801 4989
rect 92829 4961 92864 4989
rect 92704 4944 92864 4961
rect 81369 -588 81417 -560
rect 81445 -588 81479 -560
rect 81507 -588 81541 -560
rect 81569 -588 81603 -560
rect 81631 -588 81679 -560
rect 81369 -622 81679 -588
rect 81369 -650 81417 -622
rect 81445 -650 81479 -622
rect 81507 -650 81541 -622
rect 81569 -650 81603 -622
rect 81631 -650 81679 -622
rect 81369 -684 81679 -650
rect 81369 -712 81417 -684
rect 81445 -712 81479 -684
rect 81507 -712 81541 -684
rect 81569 -712 81603 -684
rect 81631 -712 81679 -684
rect 81369 -746 81679 -712
rect 81369 -774 81417 -746
rect 81445 -774 81479 -746
rect 81507 -774 81541 -746
rect 81569 -774 81603 -746
rect 81631 -774 81679 -746
rect 81369 -822 81679 -774
rect 94869 2175 95179 10961
rect 94869 2147 94917 2175
rect 94945 2147 94979 2175
rect 95007 2147 95041 2175
rect 95069 2147 95103 2175
rect 95131 2147 95179 2175
rect 94869 2113 95179 2147
rect 94869 2085 94917 2113
rect 94945 2085 94979 2113
rect 95007 2085 95041 2113
rect 95069 2085 95103 2113
rect 95131 2085 95179 2113
rect 94869 2051 95179 2085
rect 94869 2023 94917 2051
rect 94945 2023 94979 2051
rect 95007 2023 95041 2051
rect 95069 2023 95103 2051
rect 95131 2023 95179 2051
rect 94869 1989 95179 2023
rect 94869 1961 94917 1989
rect 94945 1961 94979 1989
rect 95007 1961 95041 1989
rect 95069 1961 95103 1989
rect 95131 1961 95179 1989
rect 94869 -80 95179 1961
rect 94869 -108 94917 -80
rect 94945 -108 94979 -80
rect 95007 -108 95041 -80
rect 95069 -108 95103 -80
rect 95131 -108 95179 -80
rect 94869 -142 95179 -108
rect 94869 -170 94917 -142
rect 94945 -170 94979 -142
rect 95007 -170 95041 -142
rect 95069 -170 95103 -142
rect 95131 -170 95179 -142
rect 94869 -204 95179 -170
rect 94869 -232 94917 -204
rect 94945 -232 94979 -204
rect 95007 -232 95041 -204
rect 95069 -232 95103 -204
rect 95131 -232 95179 -204
rect 94869 -266 95179 -232
rect 94869 -294 94917 -266
rect 94945 -294 94979 -266
rect 95007 -294 95041 -266
rect 95069 -294 95103 -266
rect 95131 -294 95179 -266
rect 94869 -822 95179 -294
rect 96729 299086 97039 299134
rect 96729 299058 96777 299086
rect 96805 299058 96839 299086
rect 96867 299058 96901 299086
rect 96929 299058 96963 299086
rect 96991 299058 97039 299086
rect 96729 299024 97039 299058
rect 96729 298996 96777 299024
rect 96805 298996 96839 299024
rect 96867 298996 96901 299024
rect 96929 298996 96963 299024
rect 96991 298996 97039 299024
rect 96729 298962 97039 298996
rect 96729 298934 96777 298962
rect 96805 298934 96839 298962
rect 96867 298934 96901 298962
rect 96929 298934 96963 298962
rect 96991 298934 97039 298962
rect 96729 298900 97039 298934
rect 96729 298872 96777 298900
rect 96805 298872 96839 298900
rect 96867 298872 96901 298900
rect 96929 298872 96963 298900
rect 96991 298872 97039 298900
rect 96729 293175 97039 298872
rect 96729 293147 96777 293175
rect 96805 293147 96839 293175
rect 96867 293147 96901 293175
rect 96929 293147 96963 293175
rect 96991 293147 97039 293175
rect 96729 293113 97039 293147
rect 96729 293085 96777 293113
rect 96805 293085 96839 293113
rect 96867 293085 96901 293113
rect 96929 293085 96963 293113
rect 96991 293085 97039 293113
rect 96729 293051 97039 293085
rect 96729 293023 96777 293051
rect 96805 293023 96839 293051
rect 96867 293023 96901 293051
rect 96929 293023 96963 293051
rect 96991 293023 97039 293051
rect 96729 292989 97039 293023
rect 96729 292961 96777 292989
rect 96805 292961 96839 292989
rect 96867 292961 96901 292989
rect 96929 292961 96963 292989
rect 96991 292961 97039 292989
rect 96729 284175 97039 292961
rect 96729 284147 96777 284175
rect 96805 284147 96839 284175
rect 96867 284147 96901 284175
rect 96929 284147 96963 284175
rect 96991 284147 97039 284175
rect 96729 284113 97039 284147
rect 96729 284085 96777 284113
rect 96805 284085 96839 284113
rect 96867 284085 96901 284113
rect 96929 284085 96963 284113
rect 96991 284085 97039 284113
rect 96729 284051 97039 284085
rect 96729 284023 96777 284051
rect 96805 284023 96839 284051
rect 96867 284023 96901 284051
rect 96929 284023 96963 284051
rect 96991 284023 97039 284051
rect 96729 283989 97039 284023
rect 96729 283961 96777 283989
rect 96805 283961 96839 283989
rect 96867 283961 96901 283989
rect 96929 283961 96963 283989
rect 96991 283961 97039 283989
rect 96729 275175 97039 283961
rect 96729 275147 96777 275175
rect 96805 275147 96839 275175
rect 96867 275147 96901 275175
rect 96929 275147 96963 275175
rect 96991 275147 97039 275175
rect 96729 275113 97039 275147
rect 96729 275085 96777 275113
rect 96805 275085 96839 275113
rect 96867 275085 96901 275113
rect 96929 275085 96963 275113
rect 96991 275085 97039 275113
rect 96729 275051 97039 275085
rect 96729 275023 96777 275051
rect 96805 275023 96839 275051
rect 96867 275023 96901 275051
rect 96929 275023 96963 275051
rect 96991 275023 97039 275051
rect 96729 274989 97039 275023
rect 96729 274961 96777 274989
rect 96805 274961 96839 274989
rect 96867 274961 96901 274989
rect 96929 274961 96963 274989
rect 96991 274961 97039 274989
rect 96729 266175 97039 274961
rect 96729 266147 96777 266175
rect 96805 266147 96839 266175
rect 96867 266147 96901 266175
rect 96929 266147 96963 266175
rect 96991 266147 97039 266175
rect 96729 266113 97039 266147
rect 96729 266085 96777 266113
rect 96805 266085 96839 266113
rect 96867 266085 96901 266113
rect 96929 266085 96963 266113
rect 96991 266085 97039 266113
rect 96729 266051 97039 266085
rect 96729 266023 96777 266051
rect 96805 266023 96839 266051
rect 96867 266023 96901 266051
rect 96929 266023 96963 266051
rect 96991 266023 97039 266051
rect 96729 265989 97039 266023
rect 96729 265961 96777 265989
rect 96805 265961 96839 265989
rect 96867 265961 96901 265989
rect 96929 265961 96963 265989
rect 96991 265961 97039 265989
rect 96729 257175 97039 265961
rect 96729 257147 96777 257175
rect 96805 257147 96839 257175
rect 96867 257147 96901 257175
rect 96929 257147 96963 257175
rect 96991 257147 97039 257175
rect 96729 257113 97039 257147
rect 96729 257085 96777 257113
rect 96805 257085 96839 257113
rect 96867 257085 96901 257113
rect 96929 257085 96963 257113
rect 96991 257085 97039 257113
rect 96729 257051 97039 257085
rect 96729 257023 96777 257051
rect 96805 257023 96839 257051
rect 96867 257023 96901 257051
rect 96929 257023 96963 257051
rect 96991 257023 97039 257051
rect 96729 256989 97039 257023
rect 96729 256961 96777 256989
rect 96805 256961 96839 256989
rect 96867 256961 96901 256989
rect 96929 256961 96963 256989
rect 96991 256961 97039 256989
rect 96729 248175 97039 256961
rect 96729 248147 96777 248175
rect 96805 248147 96839 248175
rect 96867 248147 96901 248175
rect 96929 248147 96963 248175
rect 96991 248147 97039 248175
rect 96729 248113 97039 248147
rect 96729 248085 96777 248113
rect 96805 248085 96839 248113
rect 96867 248085 96901 248113
rect 96929 248085 96963 248113
rect 96991 248085 97039 248113
rect 96729 248051 97039 248085
rect 96729 248023 96777 248051
rect 96805 248023 96839 248051
rect 96867 248023 96901 248051
rect 96929 248023 96963 248051
rect 96991 248023 97039 248051
rect 96729 247989 97039 248023
rect 96729 247961 96777 247989
rect 96805 247961 96839 247989
rect 96867 247961 96901 247989
rect 96929 247961 96963 247989
rect 96991 247961 97039 247989
rect 96729 239175 97039 247961
rect 96729 239147 96777 239175
rect 96805 239147 96839 239175
rect 96867 239147 96901 239175
rect 96929 239147 96963 239175
rect 96991 239147 97039 239175
rect 96729 239113 97039 239147
rect 96729 239085 96777 239113
rect 96805 239085 96839 239113
rect 96867 239085 96901 239113
rect 96929 239085 96963 239113
rect 96991 239085 97039 239113
rect 96729 239051 97039 239085
rect 96729 239023 96777 239051
rect 96805 239023 96839 239051
rect 96867 239023 96901 239051
rect 96929 239023 96963 239051
rect 96991 239023 97039 239051
rect 96729 238989 97039 239023
rect 96729 238961 96777 238989
rect 96805 238961 96839 238989
rect 96867 238961 96901 238989
rect 96929 238961 96963 238989
rect 96991 238961 97039 238989
rect 96729 230175 97039 238961
rect 96729 230147 96777 230175
rect 96805 230147 96839 230175
rect 96867 230147 96901 230175
rect 96929 230147 96963 230175
rect 96991 230147 97039 230175
rect 96729 230113 97039 230147
rect 96729 230085 96777 230113
rect 96805 230085 96839 230113
rect 96867 230085 96901 230113
rect 96929 230085 96963 230113
rect 96991 230085 97039 230113
rect 96729 230051 97039 230085
rect 96729 230023 96777 230051
rect 96805 230023 96839 230051
rect 96867 230023 96901 230051
rect 96929 230023 96963 230051
rect 96991 230023 97039 230051
rect 96729 229989 97039 230023
rect 96729 229961 96777 229989
rect 96805 229961 96839 229989
rect 96867 229961 96901 229989
rect 96929 229961 96963 229989
rect 96991 229961 97039 229989
rect 96729 221175 97039 229961
rect 96729 221147 96777 221175
rect 96805 221147 96839 221175
rect 96867 221147 96901 221175
rect 96929 221147 96963 221175
rect 96991 221147 97039 221175
rect 96729 221113 97039 221147
rect 96729 221085 96777 221113
rect 96805 221085 96839 221113
rect 96867 221085 96901 221113
rect 96929 221085 96963 221113
rect 96991 221085 97039 221113
rect 96729 221051 97039 221085
rect 96729 221023 96777 221051
rect 96805 221023 96839 221051
rect 96867 221023 96901 221051
rect 96929 221023 96963 221051
rect 96991 221023 97039 221051
rect 96729 220989 97039 221023
rect 96729 220961 96777 220989
rect 96805 220961 96839 220989
rect 96867 220961 96901 220989
rect 96929 220961 96963 220989
rect 96991 220961 97039 220989
rect 96729 212175 97039 220961
rect 96729 212147 96777 212175
rect 96805 212147 96839 212175
rect 96867 212147 96901 212175
rect 96929 212147 96963 212175
rect 96991 212147 97039 212175
rect 96729 212113 97039 212147
rect 96729 212085 96777 212113
rect 96805 212085 96839 212113
rect 96867 212085 96901 212113
rect 96929 212085 96963 212113
rect 96991 212085 97039 212113
rect 96729 212051 97039 212085
rect 96729 212023 96777 212051
rect 96805 212023 96839 212051
rect 96867 212023 96901 212051
rect 96929 212023 96963 212051
rect 96991 212023 97039 212051
rect 96729 211989 97039 212023
rect 96729 211961 96777 211989
rect 96805 211961 96839 211989
rect 96867 211961 96901 211989
rect 96929 211961 96963 211989
rect 96991 211961 97039 211989
rect 96729 203175 97039 211961
rect 96729 203147 96777 203175
rect 96805 203147 96839 203175
rect 96867 203147 96901 203175
rect 96929 203147 96963 203175
rect 96991 203147 97039 203175
rect 96729 203113 97039 203147
rect 96729 203085 96777 203113
rect 96805 203085 96839 203113
rect 96867 203085 96901 203113
rect 96929 203085 96963 203113
rect 96991 203085 97039 203113
rect 96729 203051 97039 203085
rect 96729 203023 96777 203051
rect 96805 203023 96839 203051
rect 96867 203023 96901 203051
rect 96929 203023 96963 203051
rect 96991 203023 97039 203051
rect 96729 202989 97039 203023
rect 96729 202961 96777 202989
rect 96805 202961 96839 202989
rect 96867 202961 96901 202989
rect 96929 202961 96963 202989
rect 96991 202961 97039 202989
rect 96729 194175 97039 202961
rect 96729 194147 96777 194175
rect 96805 194147 96839 194175
rect 96867 194147 96901 194175
rect 96929 194147 96963 194175
rect 96991 194147 97039 194175
rect 96729 194113 97039 194147
rect 96729 194085 96777 194113
rect 96805 194085 96839 194113
rect 96867 194085 96901 194113
rect 96929 194085 96963 194113
rect 96991 194085 97039 194113
rect 96729 194051 97039 194085
rect 96729 194023 96777 194051
rect 96805 194023 96839 194051
rect 96867 194023 96901 194051
rect 96929 194023 96963 194051
rect 96991 194023 97039 194051
rect 96729 193989 97039 194023
rect 96729 193961 96777 193989
rect 96805 193961 96839 193989
rect 96867 193961 96901 193989
rect 96929 193961 96963 193989
rect 96991 193961 97039 193989
rect 96729 185175 97039 193961
rect 96729 185147 96777 185175
rect 96805 185147 96839 185175
rect 96867 185147 96901 185175
rect 96929 185147 96963 185175
rect 96991 185147 97039 185175
rect 96729 185113 97039 185147
rect 96729 185085 96777 185113
rect 96805 185085 96839 185113
rect 96867 185085 96901 185113
rect 96929 185085 96963 185113
rect 96991 185085 97039 185113
rect 96729 185051 97039 185085
rect 96729 185023 96777 185051
rect 96805 185023 96839 185051
rect 96867 185023 96901 185051
rect 96929 185023 96963 185051
rect 96991 185023 97039 185051
rect 96729 184989 97039 185023
rect 96729 184961 96777 184989
rect 96805 184961 96839 184989
rect 96867 184961 96901 184989
rect 96929 184961 96963 184989
rect 96991 184961 97039 184989
rect 96729 176175 97039 184961
rect 96729 176147 96777 176175
rect 96805 176147 96839 176175
rect 96867 176147 96901 176175
rect 96929 176147 96963 176175
rect 96991 176147 97039 176175
rect 96729 176113 97039 176147
rect 96729 176085 96777 176113
rect 96805 176085 96839 176113
rect 96867 176085 96901 176113
rect 96929 176085 96963 176113
rect 96991 176085 97039 176113
rect 96729 176051 97039 176085
rect 96729 176023 96777 176051
rect 96805 176023 96839 176051
rect 96867 176023 96901 176051
rect 96929 176023 96963 176051
rect 96991 176023 97039 176051
rect 96729 175989 97039 176023
rect 96729 175961 96777 175989
rect 96805 175961 96839 175989
rect 96867 175961 96901 175989
rect 96929 175961 96963 175989
rect 96991 175961 97039 175989
rect 96729 167175 97039 175961
rect 110229 298606 110539 299134
rect 110229 298578 110277 298606
rect 110305 298578 110339 298606
rect 110367 298578 110401 298606
rect 110429 298578 110463 298606
rect 110491 298578 110539 298606
rect 110229 298544 110539 298578
rect 110229 298516 110277 298544
rect 110305 298516 110339 298544
rect 110367 298516 110401 298544
rect 110429 298516 110463 298544
rect 110491 298516 110539 298544
rect 110229 298482 110539 298516
rect 110229 298454 110277 298482
rect 110305 298454 110339 298482
rect 110367 298454 110401 298482
rect 110429 298454 110463 298482
rect 110491 298454 110539 298482
rect 110229 298420 110539 298454
rect 110229 298392 110277 298420
rect 110305 298392 110339 298420
rect 110367 298392 110401 298420
rect 110429 298392 110463 298420
rect 110491 298392 110539 298420
rect 110229 290175 110539 298392
rect 110229 290147 110277 290175
rect 110305 290147 110339 290175
rect 110367 290147 110401 290175
rect 110429 290147 110463 290175
rect 110491 290147 110539 290175
rect 110229 290113 110539 290147
rect 110229 290085 110277 290113
rect 110305 290085 110339 290113
rect 110367 290085 110401 290113
rect 110429 290085 110463 290113
rect 110491 290085 110539 290113
rect 110229 290051 110539 290085
rect 110229 290023 110277 290051
rect 110305 290023 110339 290051
rect 110367 290023 110401 290051
rect 110429 290023 110463 290051
rect 110491 290023 110539 290051
rect 110229 289989 110539 290023
rect 110229 289961 110277 289989
rect 110305 289961 110339 289989
rect 110367 289961 110401 289989
rect 110429 289961 110463 289989
rect 110491 289961 110539 289989
rect 110229 281175 110539 289961
rect 110229 281147 110277 281175
rect 110305 281147 110339 281175
rect 110367 281147 110401 281175
rect 110429 281147 110463 281175
rect 110491 281147 110539 281175
rect 110229 281113 110539 281147
rect 110229 281085 110277 281113
rect 110305 281085 110339 281113
rect 110367 281085 110401 281113
rect 110429 281085 110463 281113
rect 110491 281085 110539 281113
rect 110229 281051 110539 281085
rect 110229 281023 110277 281051
rect 110305 281023 110339 281051
rect 110367 281023 110401 281051
rect 110429 281023 110463 281051
rect 110491 281023 110539 281051
rect 110229 280989 110539 281023
rect 110229 280961 110277 280989
rect 110305 280961 110339 280989
rect 110367 280961 110401 280989
rect 110429 280961 110463 280989
rect 110491 280961 110539 280989
rect 110229 272175 110539 280961
rect 110229 272147 110277 272175
rect 110305 272147 110339 272175
rect 110367 272147 110401 272175
rect 110429 272147 110463 272175
rect 110491 272147 110539 272175
rect 110229 272113 110539 272147
rect 110229 272085 110277 272113
rect 110305 272085 110339 272113
rect 110367 272085 110401 272113
rect 110429 272085 110463 272113
rect 110491 272085 110539 272113
rect 110229 272051 110539 272085
rect 110229 272023 110277 272051
rect 110305 272023 110339 272051
rect 110367 272023 110401 272051
rect 110429 272023 110463 272051
rect 110491 272023 110539 272051
rect 110229 271989 110539 272023
rect 110229 271961 110277 271989
rect 110305 271961 110339 271989
rect 110367 271961 110401 271989
rect 110429 271961 110463 271989
rect 110491 271961 110539 271989
rect 110229 263175 110539 271961
rect 110229 263147 110277 263175
rect 110305 263147 110339 263175
rect 110367 263147 110401 263175
rect 110429 263147 110463 263175
rect 110491 263147 110539 263175
rect 110229 263113 110539 263147
rect 110229 263085 110277 263113
rect 110305 263085 110339 263113
rect 110367 263085 110401 263113
rect 110429 263085 110463 263113
rect 110491 263085 110539 263113
rect 110229 263051 110539 263085
rect 110229 263023 110277 263051
rect 110305 263023 110339 263051
rect 110367 263023 110401 263051
rect 110429 263023 110463 263051
rect 110491 263023 110539 263051
rect 110229 262989 110539 263023
rect 110229 262961 110277 262989
rect 110305 262961 110339 262989
rect 110367 262961 110401 262989
rect 110429 262961 110463 262989
rect 110491 262961 110539 262989
rect 110229 254175 110539 262961
rect 110229 254147 110277 254175
rect 110305 254147 110339 254175
rect 110367 254147 110401 254175
rect 110429 254147 110463 254175
rect 110491 254147 110539 254175
rect 110229 254113 110539 254147
rect 110229 254085 110277 254113
rect 110305 254085 110339 254113
rect 110367 254085 110401 254113
rect 110429 254085 110463 254113
rect 110491 254085 110539 254113
rect 110229 254051 110539 254085
rect 110229 254023 110277 254051
rect 110305 254023 110339 254051
rect 110367 254023 110401 254051
rect 110429 254023 110463 254051
rect 110491 254023 110539 254051
rect 110229 253989 110539 254023
rect 110229 253961 110277 253989
rect 110305 253961 110339 253989
rect 110367 253961 110401 253989
rect 110429 253961 110463 253989
rect 110491 253961 110539 253989
rect 110229 245175 110539 253961
rect 110229 245147 110277 245175
rect 110305 245147 110339 245175
rect 110367 245147 110401 245175
rect 110429 245147 110463 245175
rect 110491 245147 110539 245175
rect 110229 245113 110539 245147
rect 110229 245085 110277 245113
rect 110305 245085 110339 245113
rect 110367 245085 110401 245113
rect 110429 245085 110463 245113
rect 110491 245085 110539 245113
rect 110229 245051 110539 245085
rect 110229 245023 110277 245051
rect 110305 245023 110339 245051
rect 110367 245023 110401 245051
rect 110429 245023 110463 245051
rect 110491 245023 110539 245051
rect 110229 244989 110539 245023
rect 110229 244961 110277 244989
rect 110305 244961 110339 244989
rect 110367 244961 110401 244989
rect 110429 244961 110463 244989
rect 110491 244961 110539 244989
rect 110229 236175 110539 244961
rect 110229 236147 110277 236175
rect 110305 236147 110339 236175
rect 110367 236147 110401 236175
rect 110429 236147 110463 236175
rect 110491 236147 110539 236175
rect 110229 236113 110539 236147
rect 110229 236085 110277 236113
rect 110305 236085 110339 236113
rect 110367 236085 110401 236113
rect 110429 236085 110463 236113
rect 110491 236085 110539 236113
rect 110229 236051 110539 236085
rect 110229 236023 110277 236051
rect 110305 236023 110339 236051
rect 110367 236023 110401 236051
rect 110429 236023 110463 236051
rect 110491 236023 110539 236051
rect 110229 235989 110539 236023
rect 110229 235961 110277 235989
rect 110305 235961 110339 235989
rect 110367 235961 110401 235989
rect 110429 235961 110463 235989
rect 110491 235961 110539 235989
rect 110229 227175 110539 235961
rect 110229 227147 110277 227175
rect 110305 227147 110339 227175
rect 110367 227147 110401 227175
rect 110429 227147 110463 227175
rect 110491 227147 110539 227175
rect 110229 227113 110539 227147
rect 110229 227085 110277 227113
rect 110305 227085 110339 227113
rect 110367 227085 110401 227113
rect 110429 227085 110463 227113
rect 110491 227085 110539 227113
rect 110229 227051 110539 227085
rect 110229 227023 110277 227051
rect 110305 227023 110339 227051
rect 110367 227023 110401 227051
rect 110429 227023 110463 227051
rect 110491 227023 110539 227051
rect 110229 226989 110539 227023
rect 110229 226961 110277 226989
rect 110305 226961 110339 226989
rect 110367 226961 110401 226989
rect 110429 226961 110463 226989
rect 110491 226961 110539 226989
rect 110229 218175 110539 226961
rect 110229 218147 110277 218175
rect 110305 218147 110339 218175
rect 110367 218147 110401 218175
rect 110429 218147 110463 218175
rect 110491 218147 110539 218175
rect 110229 218113 110539 218147
rect 110229 218085 110277 218113
rect 110305 218085 110339 218113
rect 110367 218085 110401 218113
rect 110429 218085 110463 218113
rect 110491 218085 110539 218113
rect 110229 218051 110539 218085
rect 110229 218023 110277 218051
rect 110305 218023 110339 218051
rect 110367 218023 110401 218051
rect 110429 218023 110463 218051
rect 110491 218023 110539 218051
rect 110229 217989 110539 218023
rect 110229 217961 110277 217989
rect 110305 217961 110339 217989
rect 110367 217961 110401 217989
rect 110429 217961 110463 217989
rect 110491 217961 110539 217989
rect 110229 209175 110539 217961
rect 110229 209147 110277 209175
rect 110305 209147 110339 209175
rect 110367 209147 110401 209175
rect 110429 209147 110463 209175
rect 110491 209147 110539 209175
rect 110229 209113 110539 209147
rect 110229 209085 110277 209113
rect 110305 209085 110339 209113
rect 110367 209085 110401 209113
rect 110429 209085 110463 209113
rect 110491 209085 110539 209113
rect 110229 209051 110539 209085
rect 110229 209023 110277 209051
rect 110305 209023 110339 209051
rect 110367 209023 110401 209051
rect 110429 209023 110463 209051
rect 110491 209023 110539 209051
rect 110229 208989 110539 209023
rect 110229 208961 110277 208989
rect 110305 208961 110339 208989
rect 110367 208961 110401 208989
rect 110429 208961 110463 208989
rect 110491 208961 110539 208989
rect 110229 200175 110539 208961
rect 110229 200147 110277 200175
rect 110305 200147 110339 200175
rect 110367 200147 110401 200175
rect 110429 200147 110463 200175
rect 110491 200147 110539 200175
rect 110229 200113 110539 200147
rect 110229 200085 110277 200113
rect 110305 200085 110339 200113
rect 110367 200085 110401 200113
rect 110429 200085 110463 200113
rect 110491 200085 110539 200113
rect 110229 200051 110539 200085
rect 110229 200023 110277 200051
rect 110305 200023 110339 200051
rect 110367 200023 110401 200051
rect 110429 200023 110463 200051
rect 110491 200023 110539 200051
rect 110229 199989 110539 200023
rect 110229 199961 110277 199989
rect 110305 199961 110339 199989
rect 110367 199961 110401 199989
rect 110429 199961 110463 199989
rect 110491 199961 110539 199989
rect 110229 191175 110539 199961
rect 110229 191147 110277 191175
rect 110305 191147 110339 191175
rect 110367 191147 110401 191175
rect 110429 191147 110463 191175
rect 110491 191147 110539 191175
rect 110229 191113 110539 191147
rect 110229 191085 110277 191113
rect 110305 191085 110339 191113
rect 110367 191085 110401 191113
rect 110429 191085 110463 191113
rect 110491 191085 110539 191113
rect 110229 191051 110539 191085
rect 110229 191023 110277 191051
rect 110305 191023 110339 191051
rect 110367 191023 110401 191051
rect 110429 191023 110463 191051
rect 110491 191023 110539 191051
rect 110229 190989 110539 191023
rect 110229 190961 110277 190989
rect 110305 190961 110339 190989
rect 110367 190961 110401 190989
rect 110429 190961 110463 190989
rect 110491 190961 110539 190989
rect 110229 182175 110539 190961
rect 110229 182147 110277 182175
rect 110305 182147 110339 182175
rect 110367 182147 110401 182175
rect 110429 182147 110463 182175
rect 110491 182147 110539 182175
rect 110229 182113 110539 182147
rect 110229 182085 110277 182113
rect 110305 182085 110339 182113
rect 110367 182085 110401 182113
rect 110429 182085 110463 182113
rect 110491 182085 110539 182113
rect 110229 182051 110539 182085
rect 110229 182023 110277 182051
rect 110305 182023 110339 182051
rect 110367 182023 110401 182051
rect 110429 182023 110463 182051
rect 110491 182023 110539 182051
rect 110229 181989 110539 182023
rect 110229 181961 110277 181989
rect 110305 181961 110339 181989
rect 110367 181961 110401 181989
rect 110429 181961 110463 181989
rect 110491 181961 110539 181989
rect 100384 173175 100544 173192
rect 100384 173147 100419 173175
rect 100447 173147 100481 173175
rect 100509 173147 100544 173175
rect 100384 173113 100544 173147
rect 100384 173085 100419 173113
rect 100447 173085 100481 173113
rect 100509 173085 100544 173113
rect 100384 173051 100544 173085
rect 100384 173023 100419 173051
rect 100447 173023 100481 173051
rect 100509 173023 100544 173051
rect 100384 172989 100544 173023
rect 100384 172961 100419 172989
rect 100447 172961 100481 172989
rect 100509 172961 100544 172989
rect 100384 172944 100544 172961
rect 110229 173175 110539 181961
rect 110229 173147 110277 173175
rect 110305 173147 110339 173175
rect 110367 173147 110401 173175
rect 110429 173147 110463 173175
rect 110491 173147 110539 173175
rect 110229 173113 110539 173147
rect 110229 173085 110277 173113
rect 110305 173085 110339 173113
rect 110367 173085 110401 173113
rect 110429 173085 110463 173113
rect 110491 173085 110539 173113
rect 110229 173051 110539 173085
rect 110229 173023 110277 173051
rect 110305 173023 110339 173051
rect 110367 173023 110401 173051
rect 110429 173023 110463 173051
rect 110491 173023 110539 173051
rect 110229 172989 110539 173023
rect 110229 172961 110277 172989
rect 110305 172961 110339 172989
rect 110367 172961 110401 172989
rect 110429 172961 110463 172989
rect 110491 172961 110539 172989
rect 96729 167147 96777 167175
rect 96805 167147 96839 167175
rect 96867 167147 96901 167175
rect 96929 167147 96963 167175
rect 96991 167147 97039 167175
rect 96729 167113 97039 167147
rect 96729 167085 96777 167113
rect 96805 167085 96839 167113
rect 96867 167085 96901 167113
rect 96929 167085 96963 167113
rect 96991 167085 97039 167113
rect 96729 167051 97039 167085
rect 96729 167023 96777 167051
rect 96805 167023 96839 167051
rect 96867 167023 96901 167051
rect 96929 167023 96963 167051
rect 96991 167023 97039 167051
rect 96729 166989 97039 167023
rect 96729 166961 96777 166989
rect 96805 166961 96839 166989
rect 96867 166961 96901 166989
rect 96929 166961 96963 166989
rect 96991 166961 97039 166989
rect 96729 158175 97039 166961
rect 108064 167175 108224 167192
rect 108064 167147 108099 167175
rect 108127 167147 108161 167175
rect 108189 167147 108224 167175
rect 108064 167113 108224 167147
rect 108064 167085 108099 167113
rect 108127 167085 108161 167113
rect 108189 167085 108224 167113
rect 108064 167051 108224 167085
rect 108064 167023 108099 167051
rect 108127 167023 108161 167051
rect 108189 167023 108224 167051
rect 108064 166989 108224 167023
rect 108064 166961 108099 166989
rect 108127 166961 108161 166989
rect 108189 166961 108224 166989
rect 108064 166944 108224 166961
rect 100384 164175 100544 164192
rect 100384 164147 100419 164175
rect 100447 164147 100481 164175
rect 100509 164147 100544 164175
rect 100384 164113 100544 164147
rect 100384 164085 100419 164113
rect 100447 164085 100481 164113
rect 100509 164085 100544 164113
rect 100384 164051 100544 164085
rect 100384 164023 100419 164051
rect 100447 164023 100481 164051
rect 100509 164023 100544 164051
rect 100384 163989 100544 164023
rect 100384 163961 100419 163989
rect 100447 163961 100481 163989
rect 100509 163961 100544 163989
rect 100384 163944 100544 163961
rect 110229 164175 110539 172961
rect 110229 164147 110277 164175
rect 110305 164147 110339 164175
rect 110367 164147 110401 164175
rect 110429 164147 110463 164175
rect 110491 164147 110539 164175
rect 110229 164113 110539 164147
rect 110229 164085 110277 164113
rect 110305 164085 110339 164113
rect 110367 164085 110401 164113
rect 110429 164085 110463 164113
rect 110491 164085 110539 164113
rect 110229 164051 110539 164085
rect 110229 164023 110277 164051
rect 110305 164023 110339 164051
rect 110367 164023 110401 164051
rect 110429 164023 110463 164051
rect 110491 164023 110539 164051
rect 110229 163989 110539 164023
rect 110229 163961 110277 163989
rect 110305 163961 110339 163989
rect 110367 163961 110401 163989
rect 110429 163961 110463 163989
rect 110491 163961 110539 163989
rect 96729 158147 96777 158175
rect 96805 158147 96839 158175
rect 96867 158147 96901 158175
rect 96929 158147 96963 158175
rect 96991 158147 97039 158175
rect 96729 158113 97039 158147
rect 96729 158085 96777 158113
rect 96805 158085 96839 158113
rect 96867 158085 96901 158113
rect 96929 158085 96963 158113
rect 96991 158085 97039 158113
rect 96729 158051 97039 158085
rect 96729 158023 96777 158051
rect 96805 158023 96839 158051
rect 96867 158023 96901 158051
rect 96929 158023 96963 158051
rect 96991 158023 97039 158051
rect 96729 157989 97039 158023
rect 96729 157961 96777 157989
rect 96805 157961 96839 157989
rect 96867 157961 96901 157989
rect 96929 157961 96963 157989
rect 96991 157961 97039 157989
rect 96729 149175 97039 157961
rect 108064 158175 108224 158192
rect 108064 158147 108099 158175
rect 108127 158147 108161 158175
rect 108189 158147 108224 158175
rect 108064 158113 108224 158147
rect 108064 158085 108099 158113
rect 108127 158085 108161 158113
rect 108189 158085 108224 158113
rect 108064 158051 108224 158085
rect 108064 158023 108099 158051
rect 108127 158023 108161 158051
rect 108189 158023 108224 158051
rect 108064 157989 108224 158023
rect 108064 157961 108099 157989
rect 108127 157961 108161 157989
rect 108189 157961 108224 157989
rect 108064 157944 108224 157961
rect 100384 155175 100544 155192
rect 100384 155147 100419 155175
rect 100447 155147 100481 155175
rect 100509 155147 100544 155175
rect 100384 155113 100544 155147
rect 100384 155085 100419 155113
rect 100447 155085 100481 155113
rect 100509 155085 100544 155113
rect 100384 155051 100544 155085
rect 100384 155023 100419 155051
rect 100447 155023 100481 155051
rect 100509 155023 100544 155051
rect 100384 154989 100544 155023
rect 100384 154961 100419 154989
rect 100447 154961 100481 154989
rect 100509 154961 100544 154989
rect 100384 154944 100544 154961
rect 110229 155175 110539 163961
rect 110229 155147 110277 155175
rect 110305 155147 110339 155175
rect 110367 155147 110401 155175
rect 110429 155147 110463 155175
rect 110491 155147 110539 155175
rect 110229 155113 110539 155147
rect 110229 155085 110277 155113
rect 110305 155085 110339 155113
rect 110367 155085 110401 155113
rect 110429 155085 110463 155113
rect 110491 155085 110539 155113
rect 110229 155051 110539 155085
rect 110229 155023 110277 155051
rect 110305 155023 110339 155051
rect 110367 155023 110401 155051
rect 110429 155023 110463 155051
rect 110491 155023 110539 155051
rect 110229 154989 110539 155023
rect 110229 154961 110277 154989
rect 110305 154961 110339 154989
rect 110367 154961 110401 154989
rect 110429 154961 110463 154989
rect 110491 154961 110539 154989
rect 96729 149147 96777 149175
rect 96805 149147 96839 149175
rect 96867 149147 96901 149175
rect 96929 149147 96963 149175
rect 96991 149147 97039 149175
rect 96729 149113 97039 149147
rect 96729 149085 96777 149113
rect 96805 149085 96839 149113
rect 96867 149085 96901 149113
rect 96929 149085 96963 149113
rect 96991 149085 97039 149113
rect 96729 149051 97039 149085
rect 96729 149023 96777 149051
rect 96805 149023 96839 149051
rect 96867 149023 96901 149051
rect 96929 149023 96963 149051
rect 96991 149023 97039 149051
rect 96729 148989 97039 149023
rect 96729 148961 96777 148989
rect 96805 148961 96839 148989
rect 96867 148961 96901 148989
rect 96929 148961 96963 148989
rect 96991 148961 97039 148989
rect 96729 140175 97039 148961
rect 108064 149175 108224 149192
rect 108064 149147 108099 149175
rect 108127 149147 108161 149175
rect 108189 149147 108224 149175
rect 108064 149113 108224 149147
rect 108064 149085 108099 149113
rect 108127 149085 108161 149113
rect 108189 149085 108224 149113
rect 108064 149051 108224 149085
rect 108064 149023 108099 149051
rect 108127 149023 108161 149051
rect 108189 149023 108224 149051
rect 108064 148989 108224 149023
rect 108064 148961 108099 148989
rect 108127 148961 108161 148989
rect 108189 148961 108224 148989
rect 108064 148944 108224 148961
rect 100384 146175 100544 146192
rect 100384 146147 100419 146175
rect 100447 146147 100481 146175
rect 100509 146147 100544 146175
rect 100384 146113 100544 146147
rect 100384 146085 100419 146113
rect 100447 146085 100481 146113
rect 100509 146085 100544 146113
rect 100384 146051 100544 146085
rect 100384 146023 100419 146051
rect 100447 146023 100481 146051
rect 100509 146023 100544 146051
rect 100384 145989 100544 146023
rect 100384 145961 100419 145989
rect 100447 145961 100481 145989
rect 100509 145961 100544 145989
rect 100384 145944 100544 145961
rect 110229 146175 110539 154961
rect 110229 146147 110277 146175
rect 110305 146147 110339 146175
rect 110367 146147 110401 146175
rect 110429 146147 110463 146175
rect 110491 146147 110539 146175
rect 110229 146113 110539 146147
rect 110229 146085 110277 146113
rect 110305 146085 110339 146113
rect 110367 146085 110401 146113
rect 110429 146085 110463 146113
rect 110491 146085 110539 146113
rect 110229 146051 110539 146085
rect 110229 146023 110277 146051
rect 110305 146023 110339 146051
rect 110367 146023 110401 146051
rect 110429 146023 110463 146051
rect 110491 146023 110539 146051
rect 110229 145989 110539 146023
rect 110229 145961 110277 145989
rect 110305 145961 110339 145989
rect 110367 145961 110401 145989
rect 110429 145961 110463 145989
rect 110491 145961 110539 145989
rect 96729 140147 96777 140175
rect 96805 140147 96839 140175
rect 96867 140147 96901 140175
rect 96929 140147 96963 140175
rect 96991 140147 97039 140175
rect 96729 140113 97039 140147
rect 96729 140085 96777 140113
rect 96805 140085 96839 140113
rect 96867 140085 96901 140113
rect 96929 140085 96963 140113
rect 96991 140085 97039 140113
rect 96729 140051 97039 140085
rect 96729 140023 96777 140051
rect 96805 140023 96839 140051
rect 96867 140023 96901 140051
rect 96929 140023 96963 140051
rect 96991 140023 97039 140051
rect 96729 139989 97039 140023
rect 96729 139961 96777 139989
rect 96805 139961 96839 139989
rect 96867 139961 96901 139989
rect 96929 139961 96963 139989
rect 96991 139961 97039 139989
rect 96729 131175 97039 139961
rect 108064 140175 108224 140192
rect 108064 140147 108099 140175
rect 108127 140147 108161 140175
rect 108189 140147 108224 140175
rect 108064 140113 108224 140147
rect 108064 140085 108099 140113
rect 108127 140085 108161 140113
rect 108189 140085 108224 140113
rect 108064 140051 108224 140085
rect 108064 140023 108099 140051
rect 108127 140023 108161 140051
rect 108189 140023 108224 140051
rect 108064 139989 108224 140023
rect 108064 139961 108099 139989
rect 108127 139961 108161 139989
rect 108189 139961 108224 139989
rect 108064 139944 108224 139961
rect 100384 137175 100544 137192
rect 100384 137147 100419 137175
rect 100447 137147 100481 137175
rect 100509 137147 100544 137175
rect 100384 137113 100544 137147
rect 100384 137085 100419 137113
rect 100447 137085 100481 137113
rect 100509 137085 100544 137113
rect 100384 137051 100544 137085
rect 100384 137023 100419 137051
rect 100447 137023 100481 137051
rect 100509 137023 100544 137051
rect 100384 136989 100544 137023
rect 100384 136961 100419 136989
rect 100447 136961 100481 136989
rect 100509 136961 100544 136989
rect 100384 136944 100544 136961
rect 110229 137175 110539 145961
rect 110229 137147 110277 137175
rect 110305 137147 110339 137175
rect 110367 137147 110401 137175
rect 110429 137147 110463 137175
rect 110491 137147 110539 137175
rect 110229 137113 110539 137147
rect 110229 137085 110277 137113
rect 110305 137085 110339 137113
rect 110367 137085 110401 137113
rect 110429 137085 110463 137113
rect 110491 137085 110539 137113
rect 110229 137051 110539 137085
rect 110229 137023 110277 137051
rect 110305 137023 110339 137051
rect 110367 137023 110401 137051
rect 110429 137023 110463 137051
rect 110491 137023 110539 137051
rect 110229 136989 110539 137023
rect 110229 136961 110277 136989
rect 110305 136961 110339 136989
rect 110367 136961 110401 136989
rect 110429 136961 110463 136989
rect 110491 136961 110539 136989
rect 96729 131147 96777 131175
rect 96805 131147 96839 131175
rect 96867 131147 96901 131175
rect 96929 131147 96963 131175
rect 96991 131147 97039 131175
rect 96729 131113 97039 131147
rect 96729 131085 96777 131113
rect 96805 131085 96839 131113
rect 96867 131085 96901 131113
rect 96929 131085 96963 131113
rect 96991 131085 97039 131113
rect 96729 131051 97039 131085
rect 96729 131023 96777 131051
rect 96805 131023 96839 131051
rect 96867 131023 96901 131051
rect 96929 131023 96963 131051
rect 96991 131023 97039 131051
rect 96729 130989 97039 131023
rect 96729 130961 96777 130989
rect 96805 130961 96839 130989
rect 96867 130961 96901 130989
rect 96929 130961 96963 130989
rect 96991 130961 97039 130989
rect 96729 122175 97039 130961
rect 108064 131175 108224 131192
rect 108064 131147 108099 131175
rect 108127 131147 108161 131175
rect 108189 131147 108224 131175
rect 108064 131113 108224 131147
rect 108064 131085 108099 131113
rect 108127 131085 108161 131113
rect 108189 131085 108224 131113
rect 108064 131051 108224 131085
rect 108064 131023 108099 131051
rect 108127 131023 108161 131051
rect 108189 131023 108224 131051
rect 108064 130989 108224 131023
rect 108064 130961 108099 130989
rect 108127 130961 108161 130989
rect 108189 130961 108224 130989
rect 108064 130944 108224 130961
rect 100384 128175 100544 128192
rect 100384 128147 100419 128175
rect 100447 128147 100481 128175
rect 100509 128147 100544 128175
rect 100384 128113 100544 128147
rect 100384 128085 100419 128113
rect 100447 128085 100481 128113
rect 100509 128085 100544 128113
rect 100384 128051 100544 128085
rect 100384 128023 100419 128051
rect 100447 128023 100481 128051
rect 100509 128023 100544 128051
rect 100384 127989 100544 128023
rect 100384 127961 100419 127989
rect 100447 127961 100481 127989
rect 100509 127961 100544 127989
rect 100384 127944 100544 127961
rect 110229 128175 110539 136961
rect 110229 128147 110277 128175
rect 110305 128147 110339 128175
rect 110367 128147 110401 128175
rect 110429 128147 110463 128175
rect 110491 128147 110539 128175
rect 110229 128113 110539 128147
rect 110229 128085 110277 128113
rect 110305 128085 110339 128113
rect 110367 128085 110401 128113
rect 110429 128085 110463 128113
rect 110491 128085 110539 128113
rect 110229 128051 110539 128085
rect 110229 128023 110277 128051
rect 110305 128023 110339 128051
rect 110367 128023 110401 128051
rect 110429 128023 110463 128051
rect 110491 128023 110539 128051
rect 110229 127989 110539 128023
rect 110229 127961 110277 127989
rect 110305 127961 110339 127989
rect 110367 127961 110401 127989
rect 110429 127961 110463 127989
rect 110491 127961 110539 127989
rect 96729 122147 96777 122175
rect 96805 122147 96839 122175
rect 96867 122147 96901 122175
rect 96929 122147 96963 122175
rect 96991 122147 97039 122175
rect 96729 122113 97039 122147
rect 96729 122085 96777 122113
rect 96805 122085 96839 122113
rect 96867 122085 96901 122113
rect 96929 122085 96963 122113
rect 96991 122085 97039 122113
rect 96729 122051 97039 122085
rect 96729 122023 96777 122051
rect 96805 122023 96839 122051
rect 96867 122023 96901 122051
rect 96929 122023 96963 122051
rect 96991 122023 97039 122051
rect 96729 121989 97039 122023
rect 96729 121961 96777 121989
rect 96805 121961 96839 121989
rect 96867 121961 96901 121989
rect 96929 121961 96963 121989
rect 96991 121961 97039 121989
rect 96729 113175 97039 121961
rect 108064 122175 108224 122192
rect 108064 122147 108099 122175
rect 108127 122147 108161 122175
rect 108189 122147 108224 122175
rect 108064 122113 108224 122147
rect 108064 122085 108099 122113
rect 108127 122085 108161 122113
rect 108189 122085 108224 122113
rect 108064 122051 108224 122085
rect 108064 122023 108099 122051
rect 108127 122023 108161 122051
rect 108189 122023 108224 122051
rect 108064 121989 108224 122023
rect 108064 121961 108099 121989
rect 108127 121961 108161 121989
rect 108189 121961 108224 121989
rect 108064 121944 108224 121961
rect 100384 119175 100544 119192
rect 100384 119147 100419 119175
rect 100447 119147 100481 119175
rect 100509 119147 100544 119175
rect 100384 119113 100544 119147
rect 100384 119085 100419 119113
rect 100447 119085 100481 119113
rect 100509 119085 100544 119113
rect 100384 119051 100544 119085
rect 100384 119023 100419 119051
rect 100447 119023 100481 119051
rect 100509 119023 100544 119051
rect 100384 118989 100544 119023
rect 100384 118961 100419 118989
rect 100447 118961 100481 118989
rect 100509 118961 100544 118989
rect 100384 118944 100544 118961
rect 110229 119175 110539 127961
rect 110229 119147 110277 119175
rect 110305 119147 110339 119175
rect 110367 119147 110401 119175
rect 110429 119147 110463 119175
rect 110491 119147 110539 119175
rect 110229 119113 110539 119147
rect 110229 119085 110277 119113
rect 110305 119085 110339 119113
rect 110367 119085 110401 119113
rect 110429 119085 110463 119113
rect 110491 119085 110539 119113
rect 110229 119051 110539 119085
rect 110229 119023 110277 119051
rect 110305 119023 110339 119051
rect 110367 119023 110401 119051
rect 110429 119023 110463 119051
rect 110491 119023 110539 119051
rect 110229 118989 110539 119023
rect 110229 118961 110277 118989
rect 110305 118961 110339 118989
rect 110367 118961 110401 118989
rect 110429 118961 110463 118989
rect 110491 118961 110539 118989
rect 96729 113147 96777 113175
rect 96805 113147 96839 113175
rect 96867 113147 96901 113175
rect 96929 113147 96963 113175
rect 96991 113147 97039 113175
rect 96729 113113 97039 113147
rect 96729 113085 96777 113113
rect 96805 113085 96839 113113
rect 96867 113085 96901 113113
rect 96929 113085 96963 113113
rect 96991 113085 97039 113113
rect 96729 113051 97039 113085
rect 96729 113023 96777 113051
rect 96805 113023 96839 113051
rect 96867 113023 96901 113051
rect 96929 113023 96963 113051
rect 96991 113023 97039 113051
rect 96729 112989 97039 113023
rect 96729 112961 96777 112989
rect 96805 112961 96839 112989
rect 96867 112961 96901 112989
rect 96929 112961 96963 112989
rect 96991 112961 97039 112989
rect 96729 104175 97039 112961
rect 108064 113175 108224 113192
rect 108064 113147 108099 113175
rect 108127 113147 108161 113175
rect 108189 113147 108224 113175
rect 108064 113113 108224 113147
rect 108064 113085 108099 113113
rect 108127 113085 108161 113113
rect 108189 113085 108224 113113
rect 108064 113051 108224 113085
rect 108064 113023 108099 113051
rect 108127 113023 108161 113051
rect 108189 113023 108224 113051
rect 108064 112989 108224 113023
rect 108064 112961 108099 112989
rect 108127 112961 108161 112989
rect 108189 112961 108224 112989
rect 108064 112944 108224 112961
rect 100384 110175 100544 110192
rect 100384 110147 100419 110175
rect 100447 110147 100481 110175
rect 100509 110147 100544 110175
rect 100384 110113 100544 110147
rect 100384 110085 100419 110113
rect 100447 110085 100481 110113
rect 100509 110085 100544 110113
rect 100384 110051 100544 110085
rect 100384 110023 100419 110051
rect 100447 110023 100481 110051
rect 100509 110023 100544 110051
rect 100384 109989 100544 110023
rect 100384 109961 100419 109989
rect 100447 109961 100481 109989
rect 100509 109961 100544 109989
rect 100384 109944 100544 109961
rect 110229 110175 110539 118961
rect 110229 110147 110277 110175
rect 110305 110147 110339 110175
rect 110367 110147 110401 110175
rect 110429 110147 110463 110175
rect 110491 110147 110539 110175
rect 110229 110113 110539 110147
rect 110229 110085 110277 110113
rect 110305 110085 110339 110113
rect 110367 110085 110401 110113
rect 110429 110085 110463 110113
rect 110491 110085 110539 110113
rect 110229 110051 110539 110085
rect 110229 110023 110277 110051
rect 110305 110023 110339 110051
rect 110367 110023 110401 110051
rect 110429 110023 110463 110051
rect 110491 110023 110539 110051
rect 110229 109989 110539 110023
rect 110229 109961 110277 109989
rect 110305 109961 110339 109989
rect 110367 109961 110401 109989
rect 110429 109961 110463 109989
rect 110491 109961 110539 109989
rect 96729 104147 96777 104175
rect 96805 104147 96839 104175
rect 96867 104147 96901 104175
rect 96929 104147 96963 104175
rect 96991 104147 97039 104175
rect 96729 104113 97039 104147
rect 96729 104085 96777 104113
rect 96805 104085 96839 104113
rect 96867 104085 96901 104113
rect 96929 104085 96963 104113
rect 96991 104085 97039 104113
rect 96729 104051 97039 104085
rect 96729 104023 96777 104051
rect 96805 104023 96839 104051
rect 96867 104023 96901 104051
rect 96929 104023 96963 104051
rect 96991 104023 97039 104051
rect 96729 103989 97039 104023
rect 96729 103961 96777 103989
rect 96805 103961 96839 103989
rect 96867 103961 96901 103989
rect 96929 103961 96963 103989
rect 96991 103961 97039 103989
rect 96729 95175 97039 103961
rect 108064 104175 108224 104192
rect 108064 104147 108099 104175
rect 108127 104147 108161 104175
rect 108189 104147 108224 104175
rect 108064 104113 108224 104147
rect 108064 104085 108099 104113
rect 108127 104085 108161 104113
rect 108189 104085 108224 104113
rect 108064 104051 108224 104085
rect 108064 104023 108099 104051
rect 108127 104023 108161 104051
rect 108189 104023 108224 104051
rect 108064 103989 108224 104023
rect 108064 103961 108099 103989
rect 108127 103961 108161 103989
rect 108189 103961 108224 103989
rect 108064 103944 108224 103961
rect 100384 101175 100544 101192
rect 100384 101147 100419 101175
rect 100447 101147 100481 101175
rect 100509 101147 100544 101175
rect 100384 101113 100544 101147
rect 100384 101085 100419 101113
rect 100447 101085 100481 101113
rect 100509 101085 100544 101113
rect 100384 101051 100544 101085
rect 100384 101023 100419 101051
rect 100447 101023 100481 101051
rect 100509 101023 100544 101051
rect 100384 100989 100544 101023
rect 100384 100961 100419 100989
rect 100447 100961 100481 100989
rect 100509 100961 100544 100989
rect 100384 100944 100544 100961
rect 110229 101175 110539 109961
rect 110229 101147 110277 101175
rect 110305 101147 110339 101175
rect 110367 101147 110401 101175
rect 110429 101147 110463 101175
rect 110491 101147 110539 101175
rect 110229 101113 110539 101147
rect 110229 101085 110277 101113
rect 110305 101085 110339 101113
rect 110367 101085 110401 101113
rect 110429 101085 110463 101113
rect 110491 101085 110539 101113
rect 110229 101051 110539 101085
rect 110229 101023 110277 101051
rect 110305 101023 110339 101051
rect 110367 101023 110401 101051
rect 110429 101023 110463 101051
rect 110491 101023 110539 101051
rect 110229 100989 110539 101023
rect 110229 100961 110277 100989
rect 110305 100961 110339 100989
rect 110367 100961 110401 100989
rect 110429 100961 110463 100989
rect 110491 100961 110539 100989
rect 96729 95147 96777 95175
rect 96805 95147 96839 95175
rect 96867 95147 96901 95175
rect 96929 95147 96963 95175
rect 96991 95147 97039 95175
rect 96729 95113 97039 95147
rect 96729 95085 96777 95113
rect 96805 95085 96839 95113
rect 96867 95085 96901 95113
rect 96929 95085 96963 95113
rect 96991 95085 97039 95113
rect 96729 95051 97039 95085
rect 96729 95023 96777 95051
rect 96805 95023 96839 95051
rect 96867 95023 96901 95051
rect 96929 95023 96963 95051
rect 96991 95023 97039 95051
rect 96729 94989 97039 95023
rect 96729 94961 96777 94989
rect 96805 94961 96839 94989
rect 96867 94961 96901 94989
rect 96929 94961 96963 94989
rect 96991 94961 97039 94989
rect 96729 86175 97039 94961
rect 108064 95175 108224 95192
rect 108064 95147 108099 95175
rect 108127 95147 108161 95175
rect 108189 95147 108224 95175
rect 108064 95113 108224 95147
rect 108064 95085 108099 95113
rect 108127 95085 108161 95113
rect 108189 95085 108224 95113
rect 108064 95051 108224 95085
rect 108064 95023 108099 95051
rect 108127 95023 108161 95051
rect 108189 95023 108224 95051
rect 108064 94989 108224 95023
rect 108064 94961 108099 94989
rect 108127 94961 108161 94989
rect 108189 94961 108224 94989
rect 108064 94944 108224 94961
rect 100384 92175 100544 92192
rect 100384 92147 100419 92175
rect 100447 92147 100481 92175
rect 100509 92147 100544 92175
rect 100384 92113 100544 92147
rect 100384 92085 100419 92113
rect 100447 92085 100481 92113
rect 100509 92085 100544 92113
rect 100384 92051 100544 92085
rect 100384 92023 100419 92051
rect 100447 92023 100481 92051
rect 100509 92023 100544 92051
rect 100384 91989 100544 92023
rect 100384 91961 100419 91989
rect 100447 91961 100481 91989
rect 100509 91961 100544 91989
rect 100384 91944 100544 91961
rect 110229 92175 110539 100961
rect 110229 92147 110277 92175
rect 110305 92147 110339 92175
rect 110367 92147 110401 92175
rect 110429 92147 110463 92175
rect 110491 92147 110539 92175
rect 110229 92113 110539 92147
rect 110229 92085 110277 92113
rect 110305 92085 110339 92113
rect 110367 92085 110401 92113
rect 110429 92085 110463 92113
rect 110491 92085 110539 92113
rect 110229 92051 110539 92085
rect 110229 92023 110277 92051
rect 110305 92023 110339 92051
rect 110367 92023 110401 92051
rect 110429 92023 110463 92051
rect 110491 92023 110539 92051
rect 110229 91989 110539 92023
rect 110229 91961 110277 91989
rect 110305 91961 110339 91989
rect 110367 91961 110401 91989
rect 110429 91961 110463 91989
rect 110491 91961 110539 91989
rect 96729 86147 96777 86175
rect 96805 86147 96839 86175
rect 96867 86147 96901 86175
rect 96929 86147 96963 86175
rect 96991 86147 97039 86175
rect 96729 86113 97039 86147
rect 96729 86085 96777 86113
rect 96805 86085 96839 86113
rect 96867 86085 96901 86113
rect 96929 86085 96963 86113
rect 96991 86085 97039 86113
rect 96729 86051 97039 86085
rect 96729 86023 96777 86051
rect 96805 86023 96839 86051
rect 96867 86023 96901 86051
rect 96929 86023 96963 86051
rect 96991 86023 97039 86051
rect 96729 85989 97039 86023
rect 96729 85961 96777 85989
rect 96805 85961 96839 85989
rect 96867 85961 96901 85989
rect 96929 85961 96963 85989
rect 96991 85961 97039 85989
rect 96729 77175 97039 85961
rect 108064 86175 108224 86192
rect 108064 86147 108099 86175
rect 108127 86147 108161 86175
rect 108189 86147 108224 86175
rect 108064 86113 108224 86147
rect 108064 86085 108099 86113
rect 108127 86085 108161 86113
rect 108189 86085 108224 86113
rect 108064 86051 108224 86085
rect 108064 86023 108099 86051
rect 108127 86023 108161 86051
rect 108189 86023 108224 86051
rect 108064 85989 108224 86023
rect 108064 85961 108099 85989
rect 108127 85961 108161 85989
rect 108189 85961 108224 85989
rect 108064 85944 108224 85961
rect 100384 83175 100544 83192
rect 100384 83147 100419 83175
rect 100447 83147 100481 83175
rect 100509 83147 100544 83175
rect 100384 83113 100544 83147
rect 100384 83085 100419 83113
rect 100447 83085 100481 83113
rect 100509 83085 100544 83113
rect 100384 83051 100544 83085
rect 100384 83023 100419 83051
rect 100447 83023 100481 83051
rect 100509 83023 100544 83051
rect 100384 82989 100544 83023
rect 100384 82961 100419 82989
rect 100447 82961 100481 82989
rect 100509 82961 100544 82989
rect 100384 82944 100544 82961
rect 110229 83175 110539 91961
rect 110229 83147 110277 83175
rect 110305 83147 110339 83175
rect 110367 83147 110401 83175
rect 110429 83147 110463 83175
rect 110491 83147 110539 83175
rect 110229 83113 110539 83147
rect 110229 83085 110277 83113
rect 110305 83085 110339 83113
rect 110367 83085 110401 83113
rect 110429 83085 110463 83113
rect 110491 83085 110539 83113
rect 110229 83051 110539 83085
rect 110229 83023 110277 83051
rect 110305 83023 110339 83051
rect 110367 83023 110401 83051
rect 110429 83023 110463 83051
rect 110491 83023 110539 83051
rect 110229 82989 110539 83023
rect 110229 82961 110277 82989
rect 110305 82961 110339 82989
rect 110367 82961 110401 82989
rect 110429 82961 110463 82989
rect 110491 82961 110539 82989
rect 96729 77147 96777 77175
rect 96805 77147 96839 77175
rect 96867 77147 96901 77175
rect 96929 77147 96963 77175
rect 96991 77147 97039 77175
rect 96729 77113 97039 77147
rect 96729 77085 96777 77113
rect 96805 77085 96839 77113
rect 96867 77085 96901 77113
rect 96929 77085 96963 77113
rect 96991 77085 97039 77113
rect 96729 77051 97039 77085
rect 96729 77023 96777 77051
rect 96805 77023 96839 77051
rect 96867 77023 96901 77051
rect 96929 77023 96963 77051
rect 96991 77023 97039 77051
rect 96729 76989 97039 77023
rect 96729 76961 96777 76989
rect 96805 76961 96839 76989
rect 96867 76961 96901 76989
rect 96929 76961 96963 76989
rect 96991 76961 97039 76989
rect 96729 68175 97039 76961
rect 108064 77175 108224 77192
rect 108064 77147 108099 77175
rect 108127 77147 108161 77175
rect 108189 77147 108224 77175
rect 108064 77113 108224 77147
rect 108064 77085 108099 77113
rect 108127 77085 108161 77113
rect 108189 77085 108224 77113
rect 108064 77051 108224 77085
rect 108064 77023 108099 77051
rect 108127 77023 108161 77051
rect 108189 77023 108224 77051
rect 108064 76989 108224 77023
rect 108064 76961 108099 76989
rect 108127 76961 108161 76989
rect 108189 76961 108224 76989
rect 108064 76944 108224 76961
rect 100384 74175 100544 74192
rect 100384 74147 100419 74175
rect 100447 74147 100481 74175
rect 100509 74147 100544 74175
rect 100384 74113 100544 74147
rect 100384 74085 100419 74113
rect 100447 74085 100481 74113
rect 100509 74085 100544 74113
rect 100384 74051 100544 74085
rect 100384 74023 100419 74051
rect 100447 74023 100481 74051
rect 100509 74023 100544 74051
rect 100384 73989 100544 74023
rect 100384 73961 100419 73989
rect 100447 73961 100481 73989
rect 100509 73961 100544 73989
rect 100384 73944 100544 73961
rect 110229 74175 110539 82961
rect 110229 74147 110277 74175
rect 110305 74147 110339 74175
rect 110367 74147 110401 74175
rect 110429 74147 110463 74175
rect 110491 74147 110539 74175
rect 110229 74113 110539 74147
rect 110229 74085 110277 74113
rect 110305 74085 110339 74113
rect 110367 74085 110401 74113
rect 110429 74085 110463 74113
rect 110491 74085 110539 74113
rect 110229 74051 110539 74085
rect 110229 74023 110277 74051
rect 110305 74023 110339 74051
rect 110367 74023 110401 74051
rect 110429 74023 110463 74051
rect 110491 74023 110539 74051
rect 110229 73989 110539 74023
rect 110229 73961 110277 73989
rect 110305 73961 110339 73989
rect 110367 73961 110401 73989
rect 110429 73961 110463 73989
rect 110491 73961 110539 73989
rect 96729 68147 96777 68175
rect 96805 68147 96839 68175
rect 96867 68147 96901 68175
rect 96929 68147 96963 68175
rect 96991 68147 97039 68175
rect 96729 68113 97039 68147
rect 96729 68085 96777 68113
rect 96805 68085 96839 68113
rect 96867 68085 96901 68113
rect 96929 68085 96963 68113
rect 96991 68085 97039 68113
rect 96729 68051 97039 68085
rect 96729 68023 96777 68051
rect 96805 68023 96839 68051
rect 96867 68023 96901 68051
rect 96929 68023 96963 68051
rect 96991 68023 97039 68051
rect 96729 67989 97039 68023
rect 96729 67961 96777 67989
rect 96805 67961 96839 67989
rect 96867 67961 96901 67989
rect 96929 67961 96963 67989
rect 96991 67961 97039 67989
rect 96729 59175 97039 67961
rect 108064 68175 108224 68192
rect 108064 68147 108099 68175
rect 108127 68147 108161 68175
rect 108189 68147 108224 68175
rect 108064 68113 108224 68147
rect 108064 68085 108099 68113
rect 108127 68085 108161 68113
rect 108189 68085 108224 68113
rect 108064 68051 108224 68085
rect 108064 68023 108099 68051
rect 108127 68023 108161 68051
rect 108189 68023 108224 68051
rect 108064 67989 108224 68023
rect 108064 67961 108099 67989
rect 108127 67961 108161 67989
rect 108189 67961 108224 67989
rect 108064 67944 108224 67961
rect 100384 65175 100544 65192
rect 100384 65147 100419 65175
rect 100447 65147 100481 65175
rect 100509 65147 100544 65175
rect 100384 65113 100544 65147
rect 100384 65085 100419 65113
rect 100447 65085 100481 65113
rect 100509 65085 100544 65113
rect 100384 65051 100544 65085
rect 100384 65023 100419 65051
rect 100447 65023 100481 65051
rect 100509 65023 100544 65051
rect 100384 64989 100544 65023
rect 100384 64961 100419 64989
rect 100447 64961 100481 64989
rect 100509 64961 100544 64989
rect 100384 64944 100544 64961
rect 110229 65175 110539 73961
rect 110229 65147 110277 65175
rect 110305 65147 110339 65175
rect 110367 65147 110401 65175
rect 110429 65147 110463 65175
rect 110491 65147 110539 65175
rect 110229 65113 110539 65147
rect 110229 65085 110277 65113
rect 110305 65085 110339 65113
rect 110367 65085 110401 65113
rect 110429 65085 110463 65113
rect 110491 65085 110539 65113
rect 110229 65051 110539 65085
rect 110229 65023 110277 65051
rect 110305 65023 110339 65051
rect 110367 65023 110401 65051
rect 110429 65023 110463 65051
rect 110491 65023 110539 65051
rect 110229 64989 110539 65023
rect 110229 64961 110277 64989
rect 110305 64961 110339 64989
rect 110367 64961 110401 64989
rect 110429 64961 110463 64989
rect 110491 64961 110539 64989
rect 96729 59147 96777 59175
rect 96805 59147 96839 59175
rect 96867 59147 96901 59175
rect 96929 59147 96963 59175
rect 96991 59147 97039 59175
rect 96729 59113 97039 59147
rect 96729 59085 96777 59113
rect 96805 59085 96839 59113
rect 96867 59085 96901 59113
rect 96929 59085 96963 59113
rect 96991 59085 97039 59113
rect 96729 59051 97039 59085
rect 96729 59023 96777 59051
rect 96805 59023 96839 59051
rect 96867 59023 96901 59051
rect 96929 59023 96963 59051
rect 96991 59023 97039 59051
rect 96729 58989 97039 59023
rect 96729 58961 96777 58989
rect 96805 58961 96839 58989
rect 96867 58961 96901 58989
rect 96929 58961 96963 58989
rect 96991 58961 97039 58989
rect 96729 50175 97039 58961
rect 108064 59175 108224 59192
rect 108064 59147 108099 59175
rect 108127 59147 108161 59175
rect 108189 59147 108224 59175
rect 108064 59113 108224 59147
rect 108064 59085 108099 59113
rect 108127 59085 108161 59113
rect 108189 59085 108224 59113
rect 108064 59051 108224 59085
rect 108064 59023 108099 59051
rect 108127 59023 108161 59051
rect 108189 59023 108224 59051
rect 108064 58989 108224 59023
rect 108064 58961 108099 58989
rect 108127 58961 108161 58989
rect 108189 58961 108224 58989
rect 108064 58944 108224 58961
rect 100384 56175 100544 56192
rect 100384 56147 100419 56175
rect 100447 56147 100481 56175
rect 100509 56147 100544 56175
rect 100384 56113 100544 56147
rect 100384 56085 100419 56113
rect 100447 56085 100481 56113
rect 100509 56085 100544 56113
rect 100384 56051 100544 56085
rect 100384 56023 100419 56051
rect 100447 56023 100481 56051
rect 100509 56023 100544 56051
rect 100384 55989 100544 56023
rect 100384 55961 100419 55989
rect 100447 55961 100481 55989
rect 100509 55961 100544 55989
rect 100384 55944 100544 55961
rect 110229 56175 110539 64961
rect 110229 56147 110277 56175
rect 110305 56147 110339 56175
rect 110367 56147 110401 56175
rect 110429 56147 110463 56175
rect 110491 56147 110539 56175
rect 110229 56113 110539 56147
rect 110229 56085 110277 56113
rect 110305 56085 110339 56113
rect 110367 56085 110401 56113
rect 110429 56085 110463 56113
rect 110491 56085 110539 56113
rect 110229 56051 110539 56085
rect 110229 56023 110277 56051
rect 110305 56023 110339 56051
rect 110367 56023 110401 56051
rect 110429 56023 110463 56051
rect 110491 56023 110539 56051
rect 110229 55989 110539 56023
rect 110229 55961 110277 55989
rect 110305 55961 110339 55989
rect 110367 55961 110401 55989
rect 110429 55961 110463 55989
rect 110491 55961 110539 55989
rect 96729 50147 96777 50175
rect 96805 50147 96839 50175
rect 96867 50147 96901 50175
rect 96929 50147 96963 50175
rect 96991 50147 97039 50175
rect 96729 50113 97039 50147
rect 96729 50085 96777 50113
rect 96805 50085 96839 50113
rect 96867 50085 96901 50113
rect 96929 50085 96963 50113
rect 96991 50085 97039 50113
rect 96729 50051 97039 50085
rect 96729 50023 96777 50051
rect 96805 50023 96839 50051
rect 96867 50023 96901 50051
rect 96929 50023 96963 50051
rect 96991 50023 97039 50051
rect 96729 49989 97039 50023
rect 96729 49961 96777 49989
rect 96805 49961 96839 49989
rect 96867 49961 96901 49989
rect 96929 49961 96963 49989
rect 96991 49961 97039 49989
rect 96729 41175 97039 49961
rect 108064 50175 108224 50192
rect 108064 50147 108099 50175
rect 108127 50147 108161 50175
rect 108189 50147 108224 50175
rect 108064 50113 108224 50147
rect 108064 50085 108099 50113
rect 108127 50085 108161 50113
rect 108189 50085 108224 50113
rect 108064 50051 108224 50085
rect 108064 50023 108099 50051
rect 108127 50023 108161 50051
rect 108189 50023 108224 50051
rect 108064 49989 108224 50023
rect 108064 49961 108099 49989
rect 108127 49961 108161 49989
rect 108189 49961 108224 49989
rect 108064 49944 108224 49961
rect 100384 47175 100544 47192
rect 100384 47147 100419 47175
rect 100447 47147 100481 47175
rect 100509 47147 100544 47175
rect 100384 47113 100544 47147
rect 100384 47085 100419 47113
rect 100447 47085 100481 47113
rect 100509 47085 100544 47113
rect 100384 47051 100544 47085
rect 100384 47023 100419 47051
rect 100447 47023 100481 47051
rect 100509 47023 100544 47051
rect 100384 46989 100544 47023
rect 100384 46961 100419 46989
rect 100447 46961 100481 46989
rect 100509 46961 100544 46989
rect 100384 46944 100544 46961
rect 110229 47175 110539 55961
rect 110229 47147 110277 47175
rect 110305 47147 110339 47175
rect 110367 47147 110401 47175
rect 110429 47147 110463 47175
rect 110491 47147 110539 47175
rect 110229 47113 110539 47147
rect 110229 47085 110277 47113
rect 110305 47085 110339 47113
rect 110367 47085 110401 47113
rect 110429 47085 110463 47113
rect 110491 47085 110539 47113
rect 110229 47051 110539 47085
rect 110229 47023 110277 47051
rect 110305 47023 110339 47051
rect 110367 47023 110401 47051
rect 110429 47023 110463 47051
rect 110491 47023 110539 47051
rect 110229 46989 110539 47023
rect 110229 46961 110277 46989
rect 110305 46961 110339 46989
rect 110367 46961 110401 46989
rect 110429 46961 110463 46989
rect 110491 46961 110539 46989
rect 96729 41147 96777 41175
rect 96805 41147 96839 41175
rect 96867 41147 96901 41175
rect 96929 41147 96963 41175
rect 96991 41147 97039 41175
rect 96729 41113 97039 41147
rect 96729 41085 96777 41113
rect 96805 41085 96839 41113
rect 96867 41085 96901 41113
rect 96929 41085 96963 41113
rect 96991 41085 97039 41113
rect 96729 41051 97039 41085
rect 96729 41023 96777 41051
rect 96805 41023 96839 41051
rect 96867 41023 96901 41051
rect 96929 41023 96963 41051
rect 96991 41023 97039 41051
rect 96729 40989 97039 41023
rect 96729 40961 96777 40989
rect 96805 40961 96839 40989
rect 96867 40961 96901 40989
rect 96929 40961 96963 40989
rect 96991 40961 97039 40989
rect 96729 32175 97039 40961
rect 108064 41175 108224 41192
rect 108064 41147 108099 41175
rect 108127 41147 108161 41175
rect 108189 41147 108224 41175
rect 108064 41113 108224 41147
rect 108064 41085 108099 41113
rect 108127 41085 108161 41113
rect 108189 41085 108224 41113
rect 108064 41051 108224 41085
rect 108064 41023 108099 41051
rect 108127 41023 108161 41051
rect 108189 41023 108224 41051
rect 108064 40989 108224 41023
rect 108064 40961 108099 40989
rect 108127 40961 108161 40989
rect 108189 40961 108224 40989
rect 108064 40944 108224 40961
rect 100384 38175 100544 38192
rect 100384 38147 100419 38175
rect 100447 38147 100481 38175
rect 100509 38147 100544 38175
rect 100384 38113 100544 38147
rect 100384 38085 100419 38113
rect 100447 38085 100481 38113
rect 100509 38085 100544 38113
rect 100384 38051 100544 38085
rect 100384 38023 100419 38051
rect 100447 38023 100481 38051
rect 100509 38023 100544 38051
rect 100384 37989 100544 38023
rect 100384 37961 100419 37989
rect 100447 37961 100481 37989
rect 100509 37961 100544 37989
rect 100384 37944 100544 37961
rect 110229 38175 110539 46961
rect 110229 38147 110277 38175
rect 110305 38147 110339 38175
rect 110367 38147 110401 38175
rect 110429 38147 110463 38175
rect 110491 38147 110539 38175
rect 110229 38113 110539 38147
rect 110229 38085 110277 38113
rect 110305 38085 110339 38113
rect 110367 38085 110401 38113
rect 110429 38085 110463 38113
rect 110491 38085 110539 38113
rect 110229 38051 110539 38085
rect 110229 38023 110277 38051
rect 110305 38023 110339 38051
rect 110367 38023 110401 38051
rect 110429 38023 110463 38051
rect 110491 38023 110539 38051
rect 110229 37989 110539 38023
rect 110229 37961 110277 37989
rect 110305 37961 110339 37989
rect 110367 37961 110401 37989
rect 110429 37961 110463 37989
rect 110491 37961 110539 37989
rect 96729 32147 96777 32175
rect 96805 32147 96839 32175
rect 96867 32147 96901 32175
rect 96929 32147 96963 32175
rect 96991 32147 97039 32175
rect 96729 32113 97039 32147
rect 96729 32085 96777 32113
rect 96805 32085 96839 32113
rect 96867 32085 96901 32113
rect 96929 32085 96963 32113
rect 96991 32085 97039 32113
rect 96729 32051 97039 32085
rect 96729 32023 96777 32051
rect 96805 32023 96839 32051
rect 96867 32023 96901 32051
rect 96929 32023 96963 32051
rect 96991 32023 97039 32051
rect 96729 31989 97039 32023
rect 96729 31961 96777 31989
rect 96805 31961 96839 31989
rect 96867 31961 96901 31989
rect 96929 31961 96963 31989
rect 96991 31961 97039 31989
rect 96729 23175 97039 31961
rect 108064 32175 108224 32192
rect 108064 32147 108099 32175
rect 108127 32147 108161 32175
rect 108189 32147 108224 32175
rect 108064 32113 108224 32147
rect 108064 32085 108099 32113
rect 108127 32085 108161 32113
rect 108189 32085 108224 32113
rect 108064 32051 108224 32085
rect 108064 32023 108099 32051
rect 108127 32023 108161 32051
rect 108189 32023 108224 32051
rect 108064 31989 108224 32023
rect 108064 31961 108099 31989
rect 108127 31961 108161 31989
rect 108189 31961 108224 31989
rect 108064 31944 108224 31961
rect 100384 29175 100544 29192
rect 100384 29147 100419 29175
rect 100447 29147 100481 29175
rect 100509 29147 100544 29175
rect 100384 29113 100544 29147
rect 100384 29085 100419 29113
rect 100447 29085 100481 29113
rect 100509 29085 100544 29113
rect 100384 29051 100544 29085
rect 100384 29023 100419 29051
rect 100447 29023 100481 29051
rect 100509 29023 100544 29051
rect 100384 28989 100544 29023
rect 100384 28961 100419 28989
rect 100447 28961 100481 28989
rect 100509 28961 100544 28989
rect 100384 28944 100544 28961
rect 110229 29175 110539 37961
rect 110229 29147 110277 29175
rect 110305 29147 110339 29175
rect 110367 29147 110401 29175
rect 110429 29147 110463 29175
rect 110491 29147 110539 29175
rect 110229 29113 110539 29147
rect 110229 29085 110277 29113
rect 110305 29085 110339 29113
rect 110367 29085 110401 29113
rect 110429 29085 110463 29113
rect 110491 29085 110539 29113
rect 110229 29051 110539 29085
rect 110229 29023 110277 29051
rect 110305 29023 110339 29051
rect 110367 29023 110401 29051
rect 110429 29023 110463 29051
rect 110491 29023 110539 29051
rect 110229 28989 110539 29023
rect 110229 28961 110277 28989
rect 110305 28961 110339 28989
rect 110367 28961 110401 28989
rect 110429 28961 110463 28989
rect 110491 28961 110539 28989
rect 96729 23147 96777 23175
rect 96805 23147 96839 23175
rect 96867 23147 96901 23175
rect 96929 23147 96963 23175
rect 96991 23147 97039 23175
rect 96729 23113 97039 23147
rect 96729 23085 96777 23113
rect 96805 23085 96839 23113
rect 96867 23085 96901 23113
rect 96929 23085 96963 23113
rect 96991 23085 97039 23113
rect 96729 23051 97039 23085
rect 96729 23023 96777 23051
rect 96805 23023 96839 23051
rect 96867 23023 96901 23051
rect 96929 23023 96963 23051
rect 96991 23023 97039 23051
rect 96729 22989 97039 23023
rect 96729 22961 96777 22989
rect 96805 22961 96839 22989
rect 96867 22961 96901 22989
rect 96929 22961 96963 22989
rect 96991 22961 97039 22989
rect 96729 14175 97039 22961
rect 108064 23175 108224 23192
rect 108064 23147 108099 23175
rect 108127 23147 108161 23175
rect 108189 23147 108224 23175
rect 108064 23113 108224 23147
rect 108064 23085 108099 23113
rect 108127 23085 108161 23113
rect 108189 23085 108224 23113
rect 108064 23051 108224 23085
rect 108064 23023 108099 23051
rect 108127 23023 108161 23051
rect 108189 23023 108224 23051
rect 108064 22989 108224 23023
rect 108064 22961 108099 22989
rect 108127 22961 108161 22989
rect 108189 22961 108224 22989
rect 108064 22944 108224 22961
rect 100384 20175 100544 20192
rect 100384 20147 100419 20175
rect 100447 20147 100481 20175
rect 100509 20147 100544 20175
rect 100384 20113 100544 20147
rect 100384 20085 100419 20113
rect 100447 20085 100481 20113
rect 100509 20085 100544 20113
rect 100384 20051 100544 20085
rect 100384 20023 100419 20051
rect 100447 20023 100481 20051
rect 100509 20023 100544 20051
rect 100384 19989 100544 20023
rect 100384 19961 100419 19989
rect 100447 19961 100481 19989
rect 100509 19961 100544 19989
rect 100384 19944 100544 19961
rect 110229 20175 110539 28961
rect 110229 20147 110277 20175
rect 110305 20147 110339 20175
rect 110367 20147 110401 20175
rect 110429 20147 110463 20175
rect 110491 20147 110539 20175
rect 110229 20113 110539 20147
rect 110229 20085 110277 20113
rect 110305 20085 110339 20113
rect 110367 20085 110401 20113
rect 110429 20085 110463 20113
rect 110491 20085 110539 20113
rect 110229 20051 110539 20085
rect 110229 20023 110277 20051
rect 110305 20023 110339 20051
rect 110367 20023 110401 20051
rect 110429 20023 110463 20051
rect 110491 20023 110539 20051
rect 110229 19989 110539 20023
rect 110229 19961 110277 19989
rect 110305 19961 110339 19989
rect 110367 19961 110401 19989
rect 110429 19961 110463 19989
rect 110491 19961 110539 19989
rect 96729 14147 96777 14175
rect 96805 14147 96839 14175
rect 96867 14147 96901 14175
rect 96929 14147 96963 14175
rect 96991 14147 97039 14175
rect 96729 14113 97039 14147
rect 96729 14085 96777 14113
rect 96805 14085 96839 14113
rect 96867 14085 96901 14113
rect 96929 14085 96963 14113
rect 96991 14085 97039 14113
rect 96729 14051 97039 14085
rect 96729 14023 96777 14051
rect 96805 14023 96839 14051
rect 96867 14023 96901 14051
rect 96929 14023 96963 14051
rect 96991 14023 97039 14051
rect 96729 13989 97039 14023
rect 96729 13961 96777 13989
rect 96805 13961 96839 13989
rect 96867 13961 96901 13989
rect 96929 13961 96963 13989
rect 96991 13961 97039 13989
rect 96729 5175 97039 13961
rect 108064 14175 108224 14192
rect 108064 14147 108099 14175
rect 108127 14147 108161 14175
rect 108189 14147 108224 14175
rect 108064 14113 108224 14147
rect 108064 14085 108099 14113
rect 108127 14085 108161 14113
rect 108189 14085 108224 14113
rect 108064 14051 108224 14085
rect 108064 14023 108099 14051
rect 108127 14023 108161 14051
rect 108189 14023 108224 14051
rect 108064 13989 108224 14023
rect 108064 13961 108099 13989
rect 108127 13961 108161 13989
rect 108189 13961 108224 13989
rect 108064 13944 108224 13961
rect 100384 11175 100544 11192
rect 100384 11147 100419 11175
rect 100447 11147 100481 11175
rect 100509 11147 100544 11175
rect 100384 11113 100544 11147
rect 100384 11085 100419 11113
rect 100447 11085 100481 11113
rect 100509 11085 100544 11113
rect 100384 11051 100544 11085
rect 100384 11023 100419 11051
rect 100447 11023 100481 11051
rect 100509 11023 100544 11051
rect 100384 10989 100544 11023
rect 100384 10961 100419 10989
rect 100447 10961 100481 10989
rect 100509 10961 100544 10989
rect 100384 10944 100544 10961
rect 110229 11175 110539 19961
rect 110229 11147 110277 11175
rect 110305 11147 110339 11175
rect 110367 11147 110401 11175
rect 110429 11147 110463 11175
rect 110491 11147 110539 11175
rect 110229 11113 110539 11147
rect 110229 11085 110277 11113
rect 110305 11085 110339 11113
rect 110367 11085 110401 11113
rect 110429 11085 110463 11113
rect 110491 11085 110539 11113
rect 110229 11051 110539 11085
rect 110229 11023 110277 11051
rect 110305 11023 110339 11051
rect 110367 11023 110401 11051
rect 110429 11023 110463 11051
rect 110491 11023 110539 11051
rect 110229 10989 110539 11023
rect 110229 10961 110277 10989
rect 110305 10961 110339 10989
rect 110367 10961 110401 10989
rect 110429 10961 110463 10989
rect 110491 10961 110539 10989
rect 96729 5147 96777 5175
rect 96805 5147 96839 5175
rect 96867 5147 96901 5175
rect 96929 5147 96963 5175
rect 96991 5147 97039 5175
rect 96729 5113 97039 5147
rect 96729 5085 96777 5113
rect 96805 5085 96839 5113
rect 96867 5085 96901 5113
rect 96929 5085 96963 5113
rect 96991 5085 97039 5113
rect 96729 5051 97039 5085
rect 96729 5023 96777 5051
rect 96805 5023 96839 5051
rect 96867 5023 96901 5051
rect 96929 5023 96963 5051
rect 96991 5023 97039 5051
rect 96729 4989 97039 5023
rect 96729 4961 96777 4989
rect 96805 4961 96839 4989
rect 96867 4961 96901 4989
rect 96929 4961 96963 4989
rect 96991 4961 97039 4989
rect 96729 -560 97039 4961
rect 108064 5175 108224 5192
rect 108064 5147 108099 5175
rect 108127 5147 108161 5175
rect 108189 5147 108224 5175
rect 108064 5113 108224 5147
rect 108064 5085 108099 5113
rect 108127 5085 108161 5113
rect 108189 5085 108224 5113
rect 108064 5051 108224 5085
rect 108064 5023 108099 5051
rect 108127 5023 108161 5051
rect 108189 5023 108224 5051
rect 108064 4989 108224 5023
rect 108064 4961 108099 4989
rect 108127 4961 108161 4989
rect 108189 4961 108224 4989
rect 108064 4944 108224 4961
rect 96729 -588 96777 -560
rect 96805 -588 96839 -560
rect 96867 -588 96901 -560
rect 96929 -588 96963 -560
rect 96991 -588 97039 -560
rect 96729 -622 97039 -588
rect 96729 -650 96777 -622
rect 96805 -650 96839 -622
rect 96867 -650 96901 -622
rect 96929 -650 96963 -622
rect 96991 -650 97039 -622
rect 96729 -684 97039 -650
rect 96729 -712 96777 -684
rect 96805 -712 96839 -684
rect 96867 -712 96901 -684
rect 96929 -712 96963 -684
rect 96991 -712 97039 -684
rect 96729 -746 97039 -712
rect 96729 -774 96777 -746
rect 96805 -774 96839 -746
rect 96867 -774 96901 -746
rect 96929 -774 96963 -746
rect 96991 -774 97039 -746
rect 96729 -822 97039 -774
rect 110229 2175 110539 10961
rect 110229 2147 110277 2175
rect 110305 2147 110339 2175
rect 110367 2147 110401 2175
rect 110429 2147 110463 2175
rect 110491 2147 110539 2175
rect 110229 2113 110539 2147
rect 110229 2085 110277 2113
rect 110305 2085 110339 2113
rect 110367 2085 110401 2113
rect 110429 2085 110463 2113
rect 110491 2085 110539 2113
rect 110229 2051 110539 2085
rect 110229 2023 110277 2051
rect 110305 2023 110339 2051
rect 110367 2023 110401 2051
rect 110429 2023 110463 2051
rect 110491 2023 110539 2051
rect 110229 1989 110539 2023
rect 110229 1961 110277 1989
rect 110305 1961 110339 1989
rect 110367 1961 110401 1989
rect 110429 1961 110463 1989
rect 110491 1961 110539 1989
rect 110229 -80 110539 1961
rect 110229 -108 110277 -80
rect 110305 -108 110339 -80
rect 110367 -108 110401 -80
rect 110429 -108 110463 -80
rect 110491 -108 110539 -80
rect 110229 -142 110539 -108
rect 110229 -170 110277 -142
rect 110305 -170 110339 -142
rect 110367 -170 110401 -142
rect 110429 -170 110463 -142
rect 110491 -170 110539 -142
rect 110229 -204 110539 -170
rect 110229 -232 110277 -204
rect 110305 -232 110339 -204
rect 110367 -232 110401 -204
rect 110429 -232 110463 -204
rect 110491 -232 110539 -204
rect 110229 -266 110539 -232
rect 110229 -294 110277 -266
rect 110305 -294 110339 -266
rect 110367 -294 110401 -266
rect 110429 -294 110463 -266
rect 110491 -294 110539 -266
rect 110229 -822 110539 -294
rect 112089 299086 112399 299134
rect 112089 299058 112137 299086
rect 112165 299058 112199 299086
rect 112227 299058 112261 299086
rect 112289 299058 112323 299086
rect 112351 299058 112399 299086
rect 112089 299024 112399 299058
rect 112089 298996 112137 299024
rect 112165 298996 112199 299024
rect 112227 298996 112261 299024
rect 112289 298996 112323 299024
rect 112351 298996 112399 299024
rect 112089 298962 112399 298996
rect 112089 298934 112137 298962
rect 112165 298934 112199 298962
rect 112227 298934 112261 298962
rect 112289 298934 112323 298962
rect 112351 298934 112399 298962
rect 112089 298900 112399 298934
rect 112089 298872 112137 298900
rect 112165 298872 112199 298900
rect 112227 298872 112261 298900
rect 112289 298872 112323 298900
rect 112351 298872 112399 298900
rect 112089 293175 112399 298872
rect 112089 293147 112137 293175
rect 112165 293147 112199 293175
rect 112227 293147 112261 293175
rect 112289 293147 112323 293175
rect 112351 293147 112399 293175
rect 112089 293113 112399 293147
rect 112089 293085 112137 293113
rect 112165 293085 112199 293113
rect 112227 293085 112261 293113
rect 112289 293085 112323 293113
rect 112351 293085 112399 293113
rect 112089 293051 112399 293085
rect 112089 293023 112137 293051
rect 112165 293023 112199 293051
rect 112227 293023 112261 293051
rect 112289 293023 112323 293051
rect 112351 293023 112399 293051
rect 112089 292989 112399 293023
rect 112089 292961 112137 292989
rect 112165 292961 112199 292989
rect 112227 292961 112261 292989
rect 112289 292961 112323 292989
rect 112351 292961 112399 292989
rect 112089 284175 112399 292961
rect 112089 284147 112137 284175
rect 112165 284147 112199 284175
rect 112227 284147 112261 284175
rect 112289 284147 112323 284175
rect 112351 284147 112399 284175
rect 112089 284113 112399 284147
rect 112089 284085 112137 284113
rect 112165 284085 112199 284113
rect 112227 284085 112261 284113
rect 112289 284085 112323 284113
rect 112351 284085 112399 284113
rect 112089 284051 112399 284085
rect 112089 284023 112137 284051
rect 112165 284023 112199 284051
rect 112227 284023 112261 284051
rect 112289 284023 112323 284051
rect 112351 284023 112399 284051
rect 112089 283989 112399 284023
rect 112089 283961 112137 283989
rect 112165 283961 112199 283989
rect 112227 283961 112261 283989
rect 112289 283961 112323 283989
rect 112351 283961 112399 283989
rect 112089 275175 112399 283961
rect 112089 275147 112137 275175
rect 112165 275147 112199 275175
rect 112227 275147 112261 275175
rect 112289 275147 112323 275175
rect 112351 275147 112399 275175
rect 112089 275113 112399 275147
rect 112089 275085 112137 275113
rect 112165 275085 112199 275113
rect 112227 275085 112261 275113
rect 112289 275085 112323 275113
rect 112351 275085 112399 275113
rect 112089 275051 112399 275085
rect 112089 275023 112137 275051
rect 112165 275023 112199 275051
rect 112227 275023 112261 275051
rect 112289 275023 112323 275051
rect 112351 275023 112399 275051
rect 112089 274989 112399 275023
rect 112089 274961 112137 274989
rect 112165 274961 112199 274989
rect 112227 274961 112261 274989
rect 112289 274961 112323 274989
rect 112351 274961 112399 274989
rect 112089 266175 112399 274961
rect 112089 266147 112137 266175
rect 112165 266147 112199 266175
rect 112227 266147 112261 266175
rect 112289 266147 112323 266175
rect 112351 266147 112399 266175
rect 112089 266113 112399 266147
rect 112089 266085 112137 266113
rect 112165 266085 112199 266113
rect 112227 266085 112261 266113
rect 112289 266085 112323 266113
rect 112351 266085 112399 266113
rect 112089 266051 112399 266085
rect 112089 266023 112137 266051
rect 112165 266023 112199 266051
rect 112227 266023 112261 266051
rect 112289 266023 112323 266051
rect 112351 266023 112399 266051
rect 112089 265989 112399 266023
rect 112089 265961 112137 265989
rect 112165 265961 112199 265989
rect 112227 265961 112261 265989
rect 112289 265961 112323 265989
rect 112351 265961 112399 265989
rect 112089 257175 112399 265961
rect 112089 257147 112137 257175
rect 112165 257147 112199 257175
rect 112227 257147 112261 257175
rect 112289 257147 112323 257175
rect 112351 257147 112399 257175
rect 112089 257113 112399 257147
rect 112089 257085 112137 257113
rect 112165 257085 112199 257113
rect 112227 257085 112261 257113
rect 112289 257085 112323 257113
rect 112351 257085 112399 257113
rect 112089 257051 112399 257085
rect 112089 257023 112137 257051
rect 112165 257023 112199 257051
rect 112227 257023 112261 257051
rect 112289 257023 112323 257051
rect 112351 257023 112399 257051
rect 112089 256989 112399 257023
rect 112089 256961 112137 256989
rect 112165 256961 112199 256989
rect 112227 256961 112261 256989
rect 112289 256961 112323 256989
rect 112351 256961 112399 256989
rect 112089 248175 112399 256961
rect 112089 248147 112137 248175
rect 112165 248147 112199 248175
rect 112227 248147 112261 248175
rect 112289 248147 112323 248175
rect 112351 248147 112399 248175
rect 112089 248113 112399 248147
rect 112089 248085 112137 248113
rect 112165 248085 112199 248113
rect 112227 248085 112261 248113
rect 112289 248085 112323 248113
rect 112351 248085 112399 248113
rect 112089 248051 112399 248085
rect 112089 248023 112137 248051
rect 112165 248023 112199 248051
rect 112227 248023 112261 248051
rect 112289 248023 112323 248051
rect 112351 248023 112399 248051
rect 112089 247989 112399 248023
rect 112089 247961 112137 247989
rect 112165 247961 112199 247989
rect 112227 247961 112261 247989
rect 112289 247961 112323 247989
rect 112351 247961 112399 247989
rect 112089 239175 112399 247961
rect 112089 239147 112137 239175
rect 112165 239147 112199 239175
rect 112227 239147 112261 239175
rect 112289 239147 112323 239175
rect 112351 239147 112399 239175
rect 112089 239113 112399 239147
rect 112089 239085 112137 239113
rect 112165 239085 112199 239113
rect 112227 239085 112261 239113
rect 112289 239085 112323 239113
rect 112351 239085 112399 239113
rect 112089 239051 112399 239085
rect 112089 239023 112137 239051
rect 112165 239023 112199 239051
rect 112227 239023 112261 239051
rect 112289 239023 112323 239051
rect 112351 239023 112399 239051
rect 112089 238989 112399 239023
rect 112089 238961 112137 238989
rect 112165 238961 112199 238989
rect 112227 238961 112261 238989
rect 112289 238961 112323 238989
rect 112351 238961 112399 238989
rect 112089 230175 112399 238961
rect 112089 230147 112137 230175
rect 112165 230147 112199 230175
rect 112227 230147 112261 230175
rect 112289 230147 112323 230175
rect 112351 230147 112399 230175
rect 112089 230113 112399 230147
rect 112089 230085 112137 230113
rect 112165 230085 112199 230113
rect 112227 230085 112261 230113
rect 112289 230085 112323 230113
rect 112351 230085 112399 230113
rect 112089 230051 112399 230085
rect 112089 230023 112137 230051
rect 112165 230023 112199 230051
rect 112227 230023 112261 230051
rect 112289 230023 112323 230051
rect 112351 230023 112399 230051
rect 112089 229989 112399 230023
rect 112089 229961 112137 229989
rect 112165 229961 112199 229989
rect 112227 229961 112261 229989
rect 112289 229961 112323 229989
rect 112351 229961 112399 229989
rect 112089 221175 112399 229961
rect 112089 221147 112137 221175
rect 112165 221147 112199 221175
rect 112227 221147 112261 221175
rect 112289 221147 112323 221175
rect 112351 221147 112399 221175
rect 112089 221113 112399 221147
rect 112089 221085 112137 221113
rect 112165 221085 112199 221113
rect 112227 221085 112261 221113
rect 112289 221085 112323 221113
rect 112351 221085 112399 221113
rect 112089 221051 112399 221085
rect 112089 221023 112137 221051
rect 112165 221023 112199 221051
rect 112227 221023 112261 221051
rect 112289 221023 112323 221051
rect 112351 221023 112399 221051
rect 112089 220989 112399 221023
rect 112089 220961 112137 220989
rect 112165 220961 112199 220989
rect 112227 220961 112261 220989
rect 112289 220961 112323 220989
rect 112351 220961 112399 220989
rect 112089 212175 112399 220961
rect 112089 212147 112137 212175
rect 112165 212147 112199 212175
rect 112227 212147 112261 212175
rect 112289 212147 112323 212175
rect 112351 212147 112399 212175
rect 112089 212113 112399 212147
rect 112089 212085 112137 212113
rect 112165 212085 112199 212113
rect 112227 212085 112261 212113
rect 112289 212085 112323 212113
rect 112351 212085 112399 212113
rect 112089 212051 112399 212085
rect 112089 212023 112137 212051
rect 112165 212023 112199 212051
rect 112227 212023 112261 212051
rect 112289 212023 112323 212051
rect 112351 212023 112399 212051
rect 112089 211989 112399 212023
rect 112089 211961 112137 211989
rect 112165 211961 112199 211989
rect 112227 211961 112261 211989
rect 112289 211961 112323 211989
rect 112351 211961 112399 211989
rect 112089 203175 112399 211961
rect 112089 203147 112137 203175
rect 112165 203147 112199 203175
rect 112227 203147 112261 203175
rect 112289 203147 112323 203175
rect 112351 203147 112399 203175
rect 112089 203113 112399 203147
rect 112089 203085 112137 203113
rect 112165 203085 112199 203113
rect 112227 203085 112261 203113
rect 112289 203085 112323 203113
rect 112351 203085 112399 203113
rect 112089 203051 112399 203085
rect 112089 203023 112137 203051
rect 112165 203023 112199 203051
rect 112227 203023 112261 203051
rect 112289 203023 112323 203051
rect 112351 203023 112399 203051
rect 112089 202989 112399 203023
rect 112089 202961 112137 202989
rect 112165 202961 112199 202989
rect 112227 202961 112261 202989
rect 112289 202961 112323 202989
rect 112351 202961 112399 202989
rect 112089 194175 112399 202961
rect 112089 194147 112137 194175
rect 112165 194147 112199 194175
rect 112227 194147 112261 194175
rect 112289 194147 112323 194175
rect 112351 194147 112399 194175
rect 112089 194113 112399 194147
rect 112089 194085 112137 194113
rect 112165 194085 112199 194113
rect 112227 194085 112261 194113
rect 112289 194085 112323 194113
rect 112351 194085 112399 194113
rect 112089 194051 112399 194085
rect 112089 194023 112137 194051
rect 112165 194023 112199 194051
rect 112227 194023 112261 194051
rect 112289 194023 112323 194051
rect 112351 194023 112399 194051
rect 112089 193989 112399 194023
rect 112089 193961 112137 193989
rect 112165 193961 112199 193989
rect 112227 193961 112261 193989
rect 112289 193961 112323 193989
rect 112351 193961 112399 193989
rect 112089 185175 112399 193961
rect 112089 185147 112137 185175
rect 112165 185147 112199 185175
rect 112227 185147 112261 185175
rect 112289 185147 112323 185175
rect 112351 185147 112399 185175
rect 112089 185113 112399 185147
rect 112089 185085 112137 185113
rect 112165 185085 112199 185113
rect 112227 185085 112261 185113
rect 112289 185085 112323 185113
rect 112351 185085 112399 185113
rect 112089 185051 112399 185085
rect 112089 185023 112137 185051
rect 112165 185023 112199 185051
rect 112227 185023 112261 185051
rect 112289 185023 112323 185051
rect 112351 185023 112399 185051
rect 112089 184989 112399 185023
rect 112089 184961 112137 184989
rect 112165 184961 112199 184989
rect 112227 184961 112261 184989
rect 112289 184961 112323 184989
rect 112351 184961 112399 184989
rect 112089 176175 112399 184961
rect 112089 176147 112137 176175
rect 112165 176147 112199 176175
rect 112227 176147 112261 176175
rect 112289 176147 112323 176175
rect 112351 176147 112399 176175
rect 112089 176113 112399 176147
rect 112089 176085 112137 176113
rect 112165 176085 112199 176113
rect 112227 176085 112261 176113
rect 112289 176085 112323 176113
rect 112351 176085 112399 176113
rect 112089 176051 112399 176085
rect 112089 176023 112137 176051
rect 112165 176023 112199 176051
rect 112227 176023 112261 176051
rect 112289 176023 112323 176051
rect 112351 176023 112399 176051
rect 112089 175989 112399 176023
rect 112089 175961 112137 175989
rect 112165 175961 112199 175989
rect 112227 175961 112261 175989
rect 112289 175961 112323 175989
rect 112351 175961 112399 175989
rect 112089 167175 112399 175961
rect 125589 298606 125899 299134
rect 125589 298578 125637 298606
rect 125665 298578 125699 298606
rect 125727 298578 125761 298606
rect 125789 298578 125823 298606
rect 125851 298578 125899 298606
rect 125589 298544 125899 298578
rect 125589 298516 125637 298544
rect 125665 298516 125699 298544
rect 125727 298516 125761 298544
rect 125789 298516 125823 298544
rect 125851 298516 125899 298544
rect 125589 298482 125899 298516
rect 125589 298454 125637 298482
rect 125665 298454 125699 298482
rect 125727 298454 125761 298482
rect 125789 298454 125823 298482
rect 125851 298454 125899 298482
rect 125589 298420 125899 298454
rect 125589 298392 125637 298420
rect 125665 298392 125699 298420
rect 125727 298392 125761 298420
rect 125789 298392 125823 298420
rect 125851 298392 125899 298420
rect 125589 290175 125899 298392
rect 125589 290147 125637 290175
rect 125665 290147 125699 290175
rect 125727 290147 125761 290175
rect 125789 290147 125823 290175
rect 125851 290147 125899 290175
rect 125589 290113 125899 290147
rect 125589 290085 125637 290113
rect 125665 290085 125699 290113
rect 125727 290085 125761 290113
rect 125789 290085 125823 290113
rect 125851 290085 125899 290113
rect 125589 290051 125899 290085
rect 125589 290023 125637 290051
rect 125665 290023 125699 290051
rect 125727 290023 125761 290051
rect 125789 290023 125823 290051
rect 125851 290023 125899 290051
rect 125589 289989 125899 290023
rect 125589 289961 125637 289989
rect 125665 289961 125699 289989
rect 125727 289961 125761 289989
rect 125789 289961 125823 289989
rect 125851 289961 125899 289989
rect 125589 281175 125899 289961
rect 125589 281147 125637 281175
rect 125665 281147 125699 281175
rect 125727 281147 125761 281175
rect 125789 281147 125823 281175
rect 125851 281147 125899 281175
rect 125589 281113 125899 281147
rect 125589 281085 125637 281113
rect 125665 281085 125699 281113
rect 125727 281085 125761 281113
rect 125789 281085 125823 281113
rect 125851 281085 125899 281113
rect 125589 281051 125899 281085
rect 125589 281023 125637 281051
rect 125665 281023 125699 281051
rect 125727 281023 125761 281051
rect 125789 281023 125823 281051
rect 125851 281023 125899 281051
rect 125589 280989 125899 281023
rect 125589 280961 125637 280989
rect 125665 280961 125699 280989
rect 125727 280961 125761 280989
rect 125789 280961 125823 280989
rect 125851 280961 125899 280989
rect 125589 272175 125899 280961
rect 125589 272147 125637 272175
rect 125665 272147 125699 272175
rect 125727 272147 125761 272175
rect 125789 272147 125823 272175
rect 125851 272147 125899 272175
rect 125589 272113 125899 272147
rect 125589 272085 125637 272113
rect 125665 272085 125699 272113
rect 125727 272085 125761 272113
rect 125789 272085 125823 272113
rect 125851 272085 125899 272113
rect 125589 272051 125899 272085
rect 125589 272023 125637 272051
rect 125665 272023 125699 272051
rect 125727 272023 125761 272051
rect 125789 272023 125823 272051
rect 125851 272023 125899 272051
rect 125589 271989 125899 272023
rect 125589 271961 125637 271989
rect 125665 271961 125699 271989
rect 125727 271961 125761 271989
rect 125789 271961 125823 271989
rect 125851 271961 125899 271989
rect 125589 263175 125899 271961
rect 125589 263147 125637 263175
rect 125665 263147 125699 263175
rect 125727 263147 125761 263175
rect 125789 263147 125823 263175
rect 125851 263147 125899 263175
rect 125589 263113 125899 263147
rect 125589 263085 125637 263113
rect 125665 263085 125699 263113
rect 125727 263085 125761 263113
rect 125789 263085 125823 263113
rect 125851 263085 125899 263113
rect 125589 263051 125899 263085
rect 125589 263023 125637 263051
rect 125665 263023 125699 263051
rect 125727 263023 125761 263051
rect 125789 263023 125823 263051
rect 125851 263023 125899 263051
rect 125589 262989 125899 263023
rect 125589 262961 125637 262989
rect 125665 262961 125699 262989
rect 125727 262961 125761 262989
rect 125789 262961 125823 262989
rect 125851 262961 125899 262989
rect 125589 254175 125899 262961
rect 125589 254147 125637 254175
rect 125665 254147 125699 254175
rect 125727 254147 125761 254175
rect 125789 254147 125823 254175
rect 125851 254147 125899 254175
rect 125589 254113 125899 254147
rect 125589 254085 125637 254113
rect 125665 254085 125699 254113
rect 125727 254085 125761 254113
rect 125789 254085 125823 254113
rect 125851 254085 125899 254113
rect 125589 254051 125899 254085
rect 125589 254023 125637 254051
rect 125665 254023 125699 254051
rect 125727 254023 125761 254051
rect 125789 254023 125823 254051
rect 125851 254023 125899 254051
rect 125589 253989 125899 254023
rect 125589 253961 125637 253989
rect 125665 253961 125699 253989
rect 125727 253961 125761 253989
rect 125789 253961 125823 253989
rect 125851 253961 125899 253989
rect 125589 245175 125899 253961
rect 125589 245147 125637 245175
rect 125665 245147 125699 245175
rect 125727 245147 125761 245175
rect 125789 245147 125823 245175
rect 125851 245147 125899 245175
rect 125589 245113 125899 245147
rect 125589 245085 125637 245113
rect 125665 245085 125699 245113
rect 125727 245085 125761 245113
rect 125789 245085 125823 245113
rect 125851 245085 125899 245113
rect 125589 245051 125899 245085
rect 125589 245023 125637 245051
rect 125665 245023 125699 245051
rect 125727 245023 125761 245051
rect 125789 245023 125823 245051
rect 125851 245023 125899 245051
rect 125589 244989 125899 245023
rect 125589 244961 125637 244989
rect 125665 244961 125699 244989
rect 125727 244961 125761 244989
rect 125789 244961 125823 244989
rect 125851 244961 125899 244989
rect 125589 236175 125899 244961
rect 125589 236147 125637 236175
rect 125665 236147 125699 236175
rect 125727 236147 125761 236175
rect 125789 236147 125823 236175
rect 125851 236147 125899 236175
rect 125589 236113 125899 236147
rect 125589 236085 125637 236113
rect 125665 236085 125699 236113
rect 125727 236085 125761 236113
rect 125789 236085 125823 236113
rect 125851 236085 125899 236113
rect 125589 236051 125899 236085
rect 125589 236023 125637 236051
rect 125665 236023 125699 236051
rect 125727 236023 125761 236051
rect 125789 236023 125823 236051
rect 125851 236023 125899 236051
rect 125589 235989 125899 236023
rect 125589 235961 125637 235989
rect 125665 235961 125699 235989
rect 125727 235961 125761 235989
rect 125789 235961 125823 235989
rect 125851 235961 125899 235989
rect 125589 227175 125899 235961
rect 125589 227147 125637 227175
rect 125665 227147 125699 227175
rect 125727 227147 125761 227175
rect 125789 227147 125823 227175
rect 125851 227147 125899 227175
rect 125589 227113 125899 227147
rect 125589 227085 125637 227113
rect 125665 227085 125699 227113
rect 125727 227085 125761 227113
rect 125789 227085 125823 227113
rect 125851 227085 125899 227113
rect 125589 227051 125899 227085
rect 125589 227023 125637 227051
rect 125665 227023 125699 227051
rect 125727 227023 125761 227051
rect 125789 227023 125823 227051
rect 125851 227023 125899 227051
rect 125589 226989 125899 227023
rect 125589 226961 125637 226989
rect 125665 226961 125699 226989
rect 125727 226961 125761 226989
rect 125789 226961 125823 226989
rect 125851 226961 125899 226989
rect 125589 218175 125899 226961
rect 125589 218147 125637 218175
rect 125665 218147 125699 218175
rect 125727 218147 125761 218175
rect 125789 218147 125823 218175
rect 125851 218147 125899 218175
rect 125589 218113 125899 218147
rect 125589 218085 125637 218113
rect 125665 218085 125699 218113
rect 125727 218085 125761 218113
rect 125789 218085 125823 218113
rect 125851 218085 125899 218113
rect 125589 218051 125899 218085
rect 125589 218023 125637 218051
rect 125665 218023 125699 218051
rect 125727 218023 125761 218051
rect 125789 218023 125823 218051
rect 125851 218023 125899 218051
rect 125589 217989 125899 218023
rect 125589 217961 125637 217989
rect 125665 217961 125699 217989
rect 125727 217961 125761 217989
rect 125789 217961 125823 217989
rect 125851 217961 125899 217989
rect 125589 209175 125899 217961
rect 125589 209147 125637 209175
rect 125665 209147 125699 209175
rect 125727 209147 125761 209175
rect 125789 209147 125823 209175
rect 125851 209147 125899 209175
rect 125589 209113 125899 209147
rect 125589 209085 125637 209113
rect 125665 209085 125699 209113
rect 125727 209085 125761 209113
rect 125789 209085 125823 209113
rect 125851 209085 125899 209113
rect 125589 209051 125899 209085
rect 125589 209023 125637 209051
rect 125665 209023 125699 209051
rect 125727 209023 125761 209051
rect 125789 209023 125823 209051
rect 125851 209023 125899 209051
rect 125589 208989 125899 209023
rect 125589 208961 125637 208989
rect 125665 208961 125699 208989
rect 125727 208961 125761 208989
rect 125789 208961 125823 208989
rect 125851 208961 125899 208989
rect 125589 200175 125899 208961
rect 125589 200147 125637 200175
rect 125665 200147 125699 200175
rect 125727 200147 125761 200175
rect 125789 200147 125823 200175
rect 125851 200147 125899 200175
rect 125589 200113 125899 200147
rect 125589 200085 125637 200113
rect 125665 200085 125699 200113
rect 125727 200085 125761 200113
rect 125789 200085 125823 200113
rect 125851 200085 125899 200113
rect 125589 200051 125899 200085
rect 125589 200023 125637 200051
rect 125665 200023 125699 200051
rect 125727 200023 125761 200051
rect 125789 200023 125823 200051
rect 125851 200023 125899 200051
rect 125589 199989 125899 200023
rect 125589 199961 125637 199989
rect 125665 199961 125699 199989
rect 125727 199961 125761 199989
rect 125789 199961 125823 199989
rect 125851 199961 125899 199989
rect 125589 191175 125899 199961
rect 125589 191147 125637 191175
rect 125665 191147 125699 191175
rect 125727 191147 125761 191175
rect 125789 191147 125823 191175
rect 125851 191147 125899 191175
rect 125589 191113 125899 191147
rect 125589 191085 125637 191113
rect 125665 191085 125699 191113
rect 125727 191085 125761 191113
rect 125789 191085 125823 191113
rect 125851 191085 125899 191113
rect 125589 191051 125899 191085
rect 125589 191023 125637 191051
rect 125665 191023 125699 191051
rect 125727 191023 125761 191051
rect 125789 191023 125823 191051
rect 125851 191023 125899 191051
rect 125589 190989 125899 191023
rect 125589 190961 125637 190989
rect 125665 190961 125699 190989
rect 125727 190961 125761 190989
rect 125789 190961 125823 190989
rect 125851 190961 125899 190989
rect 125589 182175 125899 190961
rect 125589 182147 125637 182175
rect 125665 182147 125699 182175
rect 125727 182147 125761 182175
rect 125789 182147 125823 182175
rect 125851 182147 125899 182175
rect 125589 182113 125899 182147
rect 125589 182085 125637 182113
rect 125665 182085 125699 182113
rect 125727 182085 125761 182113
rect 125789 182085 125823 182113
rect 125851 182085 125899 182113
rect 125589 182051 125899 182085
rect 125589 182023 125637 182051
rect 125665 182023 125699 182051
rect 125727 182023 125761 182051
rect 125789 182023 125823 182051
rect 125851 182023 125899 182051
rect 125589 181989 125899 182023
rect 125589 181961 125637 181989
rect 125665 181961 125699 181989
rect 125727 181961 125761 181989
rect 125789 181961 125823 181989
rect 125851 181961 125899 181989
rect 115744 173175 115904 173192
rect 115744 173147 115779 173175
rect 115807 173147 115841 173175
rect 115869 173147 115904 173175
rect 115744 173113 115904 173147
rect 115744 173085 115779 173113
rect 115807 173085 115841 173113
rect 115869 173085 115904 173113
rect 115744 173051 115904 173085
rect 115744 173023 115779 173051
rect 115807 173023 115841 173051
rect 115869 173023 115904 173051
rect 115744 172989 115904 173023
rect 115744 172961 115779 172989
rect 115807 172961 115841 172989
rect 115869 172961 115904 172989
rect 115744 172944 115904 172961
rect 125589 173175 125899 181961
rect 125589 173147 125637 173175
rect 125665 173147 125699 173175
rect 125727 173147 125761 173175
rect 125789 173147 125823 173175
rect 125851 173147 125899 173175
rect 125589 173113 125899 173147
rect 125589 173085 125637 173113
rect 125665 173085 125699 173113
rect 125727 173085 125761 173113
rect 125789 173085 125823 173113
rect 125851 173085 125899 173113
rect 125589 173051 125899 173085
rect 125589 173023 125637 173051
rect 125665 173023 125699 173051
rect 125727 173023 125761 173051
rect 125789 173023 125823 173051
rect 125851 173023 125899 173051
rect 125589 172989 125899 173023
rect 125589 172961 125637 172989
rect 125665 172961 125699 172989
rect 125727 172961 125761 172989
rect 125789 172961 125823 172989
rect 125851 172961 125899 172989
rect 112089 167147 112137 167175
rect 112165 167147 112199 167175
rect 112227 167147 112261 167175
rect 112289 167147 112323 167175
rect 112351 167147 112399 167175
rect 112089 167113 112399 167147
rect 112089 167085 112137 167113
rect 112165 167085 112199 167113
rect 112227 167085 112261 167113
rect 112289 167085 112323 167113
rect 112351 167085 112399 167113
rect 112089 167051 112399 167085
rect 112089 167023 112137 167051
rect 112165 167023 112199 167051
rect 112227 167023 112261 167051
rect 112289 167023 112323 167051
rect 112351 167023 112399 167051
rect 112089 166989 112399 167023
rect 112089 166961 112137 166989
rect 112165 166961 112199 166989
rect 112227 166961 112261 166989
rect 112289 166961 112323 166989
rect 112351 166961 112399 166989
rect 112089 158175 112399 166961
rect 123424 167175 123584 167192
rect 123424 167147 123459 167175
rect 123487 167147 123521 167175
rect 123549 167147 123584 167175
rect 123424 167113 123584 167147
rect 123424 167085 123459 167113
rect 123487 167085 123521 167113
rect 123549 167085 123584 167113
rect 123424 167051 123584 167085
rect 123424 167023 123459 167051
rect 123487 167023 123521 167051
rect 123549 167023 123584 167051
rect 123424 166989 123584 167023
rect 123424 166961 123459 166989
rect 123487 166961 123521 166989
rect 123549 166961 123584 166989
rect 123424 166944 123584 166961
rect 115744 164175 115904 164192
rect 115744 164147 115779 164175
rect 115807 164147 115841 164175
rect 115869 164147 115904 164175
rect 115744 164113 115904 164147
rect 115744 164085 115779 164113
rect 115807 164085 115841 164113
rect 115869 164085 115904 164113
rect 115744 164051 115904 164085
rect 115744 164023 115779 164051
rect 115807 164023 115841 164051
rect 115869 164023 115904 164051
rect 115744 163989 115904 164023
rect 115744 163961 115779 163989
rect 115807 163961 115841 163989
rect 115869 163961 115904 163989
rect 115744 163944 115904 163961
rect 125589 164175 125899 172961
rect 125589 164147 125637 164175
rect 125665 164147 125699 164175
rect 125727 164147 125761 164175
rect 125789 164147 125823 164175
rect 125851 164147 125899 164175
rect 125589 164113 125899 164147
rect 125589 164085 125637 164113
rect 125665 164085 125699 164113
rect 125727 164085 125761 164113
rect 125789 164085 125823 164113
rect 125851 164085 125899 164113
rect 125589 164051 125899 164085
rect 125589 164023 125637 164051
rect 125665 164023 125699 164051
rect 125727 164023 125761 164051
rect 125789 164023 125823 164051
rect 125851 164023 125899 164051
rect 125589 163989 125899 164023
rect 125589 163961 125637 163989
rect 125665 163961 125699 163989
rect 125727 163961 125761 163989
rect 125789 163961 125823 163989
rect 125851 163961 125899 163989
rect 112089 158147 112137 158175
rect 112165 158147 112199 158175
rect 112227 158147 112261 158175
rect 112289 158147 112323 158175
rect 112351 158147 112399 158175
rect 112089 158113 112399 158147
rect 112089 158085 112137 158113
rect 112165 158085 112199 158113
rect 112227 158085 112261 158113
rect 112289 158085 112323 158113
rect 112351 158085 112399 158113
rect 112089 158051 112399 158085
rect 112089 158023 112137 158051
rect 112165 158023 112199 158051
rect 112227 158023 112261 158051
rect 112289 158023 112323 158051
rect 112351 158023 112399 158051
rect 112089 157989 112399 158023
rect 112089 157961 112137 157989
rect 112165 157961 112199 157989
rect 112227 157961 112261 157989
rect 112289 157961 112323 157989
rect 112351 157961 112399 157989
rect 112089 149175 112399 157961
rect 123424 158175 123584 158192
rect 123424 158147 123459 158175
rect 123487 158147 123521 158175
rect 123549 158147 123584 158175
rect 123424 158113 123584 158147
rect 123424 158085 123459 158113
rect 123487 158085 123521 158113
rect 123549 158085 123584 158113
rect 123424 158051 123584 158085
rect 123424 158023 123459 158051
rect 123487 158023 123521 158051
rect 123549 158023 123584 158051
rect 123424 157989 123584 158023
rect 123424 157961 123459 157989
rect 123487 157961 123521 157989
rect 123549 157961 123584 157989
rect 123424 157944 123584 157961
rect 115744 155175 115904 155192
rect 115744 155147 115779 155175
rect 115807 155147 115841 155175
rect 115869 155147 115904 155175
rect 115744 155113 115904 155147
rect 115744 155085 115779 155113
rect 115807 155085 115841 155113
rect 115869 155085 115904 155113
rect 115744 155051 115904 155085
rect 115744 155023 115779 155051
rect 115807 155023 115841 155051
rect 115869 155023 115904 155051
rect 115744 154989 115904 155023
rect 115744 154961 115779 154989
rect 115807 154961 115841 154989
rect 115869 154961 115904 154989
rect 115744 154944 115904 154961
rect 125589 155175 125899 163961
rect 125589 155147 125637 155175
rect 125665 155147 125699 155175
rect 125727 155147 125761 155175
rect 125789 155147 125823 155175
rect 125851 155147 125899 155175
rect 125589 155113 125899 155147
rect 125589 155085 125637 155113
rect 125665 155085 125699 155113
rect 125727 155085 125761 155113
rect 125789 155085 125823 155113
rect 125851 155085 125899 155113
rect 125589 155051 125899 155085
rect 125589 155023 125637 155051
rect 125665 155023 125699 155051
rect 125727 155023 125761 155051
rect 125789 155023 125823 155051
rect 125851 155023 125899 155051
rect 125589 154989 125899 155023
rect 125589 154961 125637 154989
rect 125665 154961 125699 154989
rect 125727 154961 125761 154989
rect 125789 154961 125823 154989
rect 125851 154961 125899 154989
rect 112089 149147 112137 149175
rect 112165 149147 112199 149175
rect 112227 149147 112261 149175
rect 112289 149147 112323 149175
rect 112351 149147 112399 149175
rect 112089 149113 112399 149147
rect 112089 149085 112137 149113
rect 112165 149085 112199 149113
rect 112227 149085 112261 149113
rect 112289 149085 112323 149113
rect 112351 149085 112399 149113
rect 112089 149051 112399 149085
rect 112089 149023 112137 149051
rect 112165 149023 112199 149051
rect 112227 149023 112261 149051
rect 112289 149023 112323 149051
rect 112351 149023 112399 149051
rect 112089 148989 112399 149023
rect 112089 148961 112137 148989
rect 112165 148961 112199 148989
rect 112227 148961 112261 148989
rect 112289 148961 112323 148989
rect 112351 148961 112399 148989
rect 112089 140175 112399 148961
rect 123424 149175 123584 149192
rect 123424 149147 123459 149175
rect 123487 149147 123521 149175
rect 123549 149147 123584 149175
rect 123424 149113 123584 149147
rect 123424 149085 123459 149113
rect 123487 149085 123521 149113
rect 123549 149085 123584 149113
rect 123424 149051 123584 149085
rect 123424 149023 123459 149051
rect 123487 149023 123521 149051
rect 123549 149023 123584 149051
rect 123424 148989 123584 149023
rect 123424 148961 123459 148989
rect 123487 148961 123521 148989
rect 123549 148961 123584 148989
rect 123424 148944 123584 148961
rect 115744 146175 115904 146192
rect 115744 146147 115779 146175
rect 115807 146147 115841 146175
rect 115869 146147 115904 146175
rect 115744 146113 115904 146147
rect 115744 146085 115779 146113
rect 115807 146085 115841 146113
rect 115869 146085 115904 146113
rect 115744 146051 115904 146085
rect 115744 146023 115779 146051
rect 115807 146023 115841 146051
rect 115869 146023 115904 146051
rect 115744 145989 115904 146023
rect 115744 145961 115779 145989
rect 115807 145961 115841 145989
rect 115869 145961 115904 145989
rect 115744 145944 115904 145961
rect 125589 146175 125899 154961
rect 125589 146147 125637 146175
rect 125665 146147 125699 146175
rect 125727 146147 125761 146175
rect 125789 146147 125823 146175
rect 125851 146147 125899 146175
rect 125589 146113 125899 146147
rect 125589 146085 125637 146113
rect 125665 146085 125699 146113
rect 125727 146085 125761 146113
rect 125789 146085 125823 146113
rect 125851 146085 125899 146113
rect 125589 146051 125899 146085
rect 125589 146023 125637 146051
rect 125665 146023 125699 146051
rect 125727 146023 125761 146051
rect 125789 146023 125823 146051
rect 125851 146023 125899 146051
rect 125589 145989 125899 146023
rect 125589 145961 125637 145989
rect 125665 145961 125699 145989
rect 125727 145961 125761 145989
rect 125789 145961 125823 145989
rect 125851 145961 125899 145989
rect 112089 140147 112137 140175
rect 112165 140147 112199 140175
rect 112227 140147 112261 140175
rect 112289 140147 112323 140175
rect 112351 140147 112399 140175
rect 112089 140113 112399 140147
rect 112089 140085 112137 140113
rect 112165 140085 112199 140113
rect 112227 140085 112261 140113
rect 112289 140085 112323 140113
rect 112351 140085 112399 140113
rect 112089 140051 112399 140085
rect 112089 140023 112137 140051
rect 112165 140023 112199 140051
rect 112227 140023 112261 140051
rect 112289 140023 112323 140051
rect 112351 140023 112399 140051
rect 112089 139989 112399 140023
rect 112089 139961 112137 139989
rect 112165 139961 112199 139989
rect 112227 139961 112261 139989
rect 112289 139961 112323 139989
rect 112351 139961 112399 139989
rect 112089 131175 112399 139961
rect 123424 140175 123584 140192
rect 123424 140147 123459 140175
rect 123487 140147 123521 140175
rect 123549 140147 123584 140175
rect 123424 140113 123584 140147
rect 123424 140085 123459 140113
rect 123487 140085 123521 140113
rect 123549 140085 123584 140113
rect 123424 140051 123584 140085
rect 123424 140023 123459 140051
rect 123487 140023 123521 140051
rect 123549 140023 123584 140051
rect 123424 139989 123584 140023
rect 123424 139961 123459 139989
rect 123487 139961 123521 139989
rect 123549 139961 123584 139989
rect 123424 139944 123584 139961
rect 115744 137175 115904 137192
rect 115744 137147 115779 137175
rect 115807 137147 115841 137175
rect 115869 137147 115904 137175
rect 115744 137113 115904 137147
rect 115744 137085 115779 137113
rect 115807 137085 115841 137113
rect 115869 137085 115904 137113
rect 115744 137051 115904 137085
rect 115744 137023 115779 137051
rect 115807 137023 115841 137051
rect 115869 137023 115904 137051
rect 115744 136989 115904 137023
rect 115744 136961 115779 136989
rect 115807 136961 115841 136989
rect 115869 136961 115904 136989
rect 115744 136944 115904 136961
rect 125589 137175 125899 145961
rect 125589 137147 125637 137175
rect 125665 137147 125699 137175
rect 125727 137147 125761 137175
rect 125789 137147 125823 137175
rect 125851 137147 125899 137175
rect 125589 137113 125899 137147
rect 125589 137085 125637 137113
rect 125665 137085 125699 137113
rect 125727 137085 125761 137113
rect 125789 137085 125823 137113
rect 125851 137085 125899 137113
rect 125589 137051 125899 137085
rect 125589 137023 125637 137051
rect 125665 137023 125699 137051
rect 125727 137023 125761 137051
rect 125789 137023 125823 137051
rect 125851 137023 125899 137051
rect 125589 136989 125899 137023
rect 125589 136961 125637 136989
rect 125665 136961 125699 136989
rect 125727 136961 125761 136989
rect 125789 136961 125823 136989
rect 125851 136961 125899 136989
rect 112089 131147 112137 131175
rect 112165 131147 112199 131175
rect 112227 131147 112261 131175
rect 112289 131147 112323 131175
rect 112351 131147 112399 131175
rect 112089 131113 112399 131147
rect 112089 131085 112137 131113
rect 112165 131085 112199 131113
rect 112227 131085 112261 131113
rect 112289 131085 112323 131113
rect 112351 131085 112399 131113
rect 112089 131051 112399 131085
rect 112089 131023 112137 131051
rect 112165 131023 112199 131051
rect 112227 131023 112261 131051
rect 112289 131023 112323 131051
rect 112351 131023 112399 131051
rect 112089 130989 112399 131023
rect 112089 130961 112137 130989
rect 112165 130961 112199 130989
rect 112227 130961 112261 130989
rect 112289 130961 112323 130989
rect 112351 130961 112399 130989
rect 112089 122175 112399 130961
rect 123424 131175 123584 131192
rect 123424 131147 123459 131175
rect 123487 131147 123521 131175
rect 123549 131147 123584 131175
rect 123424 131113 123584 131147
rect 123424 131085 123459 131113
rect 123487 131085 123521 131113
rect 123549 131085 123584 131113
rect 123424 131051 123584 131085
rect 123424 131023 123459 131051
rect 123487 131023 123521 131051
rect 123549 131023 123584 131051
rect 123424 130989 123584 131023
rect 123424 130961 123459 130989
rect 123487 130961 123521 130989
rect 123549 130961 123584 130989
rect 123424 130944 123584 130961
rect 115744 128175 115904 128192
rect 115744 128147 115779 128175
rect 115807 128147 115841 128175
rect 115869 128147 115904 128175
rect 115744 128113 115904 128147
rect 115744 128085 115779 128113
rect 115807 128085 115841 128113
rect 115869 128085 115904 128113
rect 115744 128051 115904 128085
rect 115744 128023 115779 128051
rect 115807 128023 115841 128051
rect 115869 128023 115904 128051
rect 115744 127989 115904 128023
rect 115744 127961 115779 127989
rect 115807 127961 115841 127989
rect 115869 127961 115904 127989
rect 115744 127944 115904 127961
rect 125589 128175 125899 136961
rect 125589 128147 125637 128175
rect 125665 128147 125699 128175
rect 125727 128147 125761 128175
rect 125789 128147 125823 128175
rect 125851 128147 125899 128175
rect 125589 128113 125899 128147
rect 125589 128085 125637 128113
rect 125665 128085 125699 128113
rect 125727 128085 125761 128113
rect 125789 128085 125823 128113
rect 125851 128085 125899 128113
rect 125589 128051 125899 128085
rect 125589 128023 125637 128051
rect 125665 128023 125699 128051
rect 125727 128023 125761 128051
rect 125789 128023 125823 128051
rect 125851 128023 125899 128051
rect 125589 127989 125899 128023
rect 125589 127961 125637 127989
rect 125665 127961 125699 127989
rect 125727 127961 125761 127989
rect 125789 127961 125823 127989
rect 125851 127961 125899 127989
rect 112089 122147 112137 122175
rect 112165 122147 112199 122175
rect 112227 122147 112261 122175
rect 112289 122147 112323 122175
rect 112351 122147 112399 122175
rect 112089 122113 112399 122147
rect 112089 122085 112137 122113
rect 112165 122085 112199 122113
rect 112227 122085 112261 122113
rect 112289 122085 112323 122113
rect 112351 122085 112399 122113
rect 112089 122051 112399 122085
rect 112089 122023 112137 122051
rect 112165 122023 112199 122051
rect 112227 122023 112261 122051
rect 112289 122023 112323 122051
rect 112351 122023 112399 122051
rect 112089 121989 112399 122023
rect 112089 121961 112137 121989
rect 112165 121961 112199 121989
rect 112227 121961 112261 121989
rect 112289 121961 112323 121989
rect 112351 121961 112399 121989
rect 112089 113175 112399 121961
rect 123424 122175 123584 122192
rect 123424 122147 123459 122175
rect 123487 122147 123521 122175
rect 123549 122147 123584 122175
rect 123424 122113 123584 122147
rect 123424 122085 123459 122113
rect 123487 122085 123521 122113
rect 123549 122085 123584 122113
rect 123424 122051 123584 122085
rect 123424 122023 123459 122051
rect 123487 122023 123521 122051
rect 123549 122023 123584 122051
rect 123424 121989 123584 122023
rect 123424 121961 123459 121989
rect 123487 121961 123521 121989
rect 123549 121961 123584 121989
rect 123424 121944 123584 121961
rect 115744 119175 115904 119192
rect 115744 119147 115779 119175
rect 115807 119147 115841 119175
rect 115869 119147 115904 119175
rect 115744 119113 115904 119147
rect 115744 119085 115779 119113
rect 115807 119085 115841 119113
rect 115869 119085 115904 119113
rect 115744 119051 115904 119085
rect 115744 119023 115779 119051
rect 115807 119023 115841 119051
rect 115869 119023 115904 119051
rect 115744 118989 115904 119023
rect 115744 118961 115779 118989
rect 115807 118961 115841 118989
rect 115869 118961 115904 118989
rect 115744 118944 115904 118961
rect 125589 119175 125899 127961
rect 125589 119147 125637 119175
rect 125665 119147 125699 119175
rect 125727 119147 125761 119175
rect 125789 119147 125823 119175
rect 125851 119147 125899 119175
rect 125589 119113 125899 119147
rect 125589 119085 125637 119113
rect 125665 119085 125699 119113
rect 125727 119085 125761 119113
rect 125789 119085 125823 119113
rect 125851 119085 125899 119113
rect 125589 119051 125899 119085
rect 125589 119023 125637 119051
rect 125665 119023 125699 119051
rect 125727 119023 125761 119051
rect 125789 119023 125823 119051
rect 125851 119023 125899 119051
rect 125589 118989 125899 119023
rect 125589 118961 125637 118989
rect 125665 118961 125699 118989
rect 125727 118961 125761 118989
rect 125789 118961 125823 118989
rect 125851 118961 125899 118989
rect 112089 113147 112137 113175
rect 112165 113147 112199 113175
rect 112227 113147 112261 113175
rect 112289 113147 112323 113175
rect 112351 113147 112399 113175
rect 112089 113113 112399 113147
rect 112089 113085 112137 113113
rect 112165 113085 112199 113113
rect 112227 113085 112261 113113
rect 112289 113085 112323 113113
rect 112351 113085 112399 113113
rect 112089 113051 112399 113085
rect 112089 113023 112137 113051
rect 112165 113023 112199 113051
rect 112227 113023 112261 113051
rect 112289 113023 112323 113051
rect 112351 113023 112399 113051
rect 112089 112989 112399 113023
rect 112089 112961 112137 112989
rect 112165 112961 112199 112989
rect 112227 112961 112261 112989
rect 112289 112961 112323 112989
rect 112351 112961 112399 112989
rect 112089 104175 112399 112961
rect 123424 113175 123584 113192
rect 123424 113147 123459 113175
rect 123487 113147 123521 113175
rect 123549 113147 123584 113175
rect 123424 113113 123584 113147
rect 123424 113085 123459 113113
rect 123487 113085 123521 113113
rect 123549 113085 123584 113113
rect 123424 113051 123584 113085
rect 123424 113023 123459 113051
rect 123487 113023 123521 113051
rect 123549 113023 123584 113051
rect 123424 112989 123584 113023
rect 123424 112961 123459 112989
rect 123487 112961 123521 112989
rect 123549 112961 123584 112989
rect 123424 112944 123584 112961
rect 115744 110175 115904 110192
rect 115744 110147 115779 110175
rect 115807 110147 115841 110175
rect 115869 110147 115904 110175
rect 115744 110113 115904 110147
rect 115744 110085 115779 110113
rect 115807 110085 115841 110113
rect 115869 110085 115904 110113
rect 115744 110051 115904 110085
rect 115744 110023 115779 110051
rect 115807 110023 115841 110051
rect 115869 110023 115904 110051
rect 115744 109989 115904 110023
rect 115744 109961 115779 109989
rect 115807 109961 115841 109989
rect 115869 109961 115904 109989
rect 115744 109944 115904 109961
rect 125589 110175 125899 118961
rect 125589 110147 125637 110175
rect 125665 110147 125699 110175
rect 125727 110147 125761 110175
rect 125789 110147 125823 110175
rect 125851 110147 125899 110175
rect 125589 110113 125899 110147
rect 125589 110085 125637 110113
rect 125665 110085 125699 110113
rect 125727 110085 125761 110113
rect 125789 110085 125823 110113
rect 125851 110085 125899 110113
rect 125589 110051 125899 110085
rect 125589 110023 125637 110051
rect 125665 110023 125699 110051
rect 125727 110023 125761 110051
rect 125789 110023 125823 110051
rect 125851 110023 125899 110051
rect 125589 109989 125899 110023
rect 125589 109961 125637 109989
rect 125665 109961 125699 109989
rect 125727 109961 125761 109989
rect 125789 109961 125823 109989
rect 125851 109961 125899 109989
rect 112089 104147 112137 104175
rect 112165 104147 112199 104175
rect 112227 104147 112261 104175
rect 112289 104147 112323 104175
rect 112351 104147 112399 104175
rect 112089 104113 112399 104147
rect 112089 104085 112137 104113
rect 112165 104085 112199 104113
rect 112227 104085 112261 104113
rect 112289 104085 112323 104113
rect 112351 104085 112399 104113
rect 112089 104051 112399 104085
rect 112089 104023 112137 104051
rect 112165 104023 112199 104051
rect 112227 104023 112261 104051
rect 112289 104023 112323 104051
rect 112351 104023 112399 104051
rect 112089 103989 112399 104023
rect 112089 103961 112137 103989
rect 112165 103961 112199 103989
rect 112227 103961 112261 103989
rect 112289 103961 112323 103989
rect 112351 103961 112399 103989
rect 112089 95175 112399 103961
rect 123424 104175 123584 104192
rect 123424 104147 123459 104175
rect 123487 104147 123521 104175
rect 123549 104147 123584 104175
rect 123424 104113 123584 104147
rect 123424 104085 123459 104113
rect 123487 104085 123521 104113
rect 123549 104085 123584 104113
rect 123424 104051 123584 104085
rect 123424 104023 123459 104051
rect 123487 104023 123521 104051
rect 123549 104023 123584 104051
rect 123424 103989 123584 104023
rect 123424 103961 123459 103989
rect 123487 103961 123521 103989
rect 123549 103961 123584 103989
rect 123424 103944 123584 103961
rect 115744 101175 115904 101192
rect 115744 101147 115779 101175
rect 115807 101147 115841 101175
rect 115869 101147 115904 101175
rect 115744 101113 115904 101147
rect 115744 101085 115779 101113
rect 115807 101085 115841 101113
rect 115869 101085 115904 101113
rect 115744 101051 115904 101085
rect 115744 101023 115779 101051
rect 115807 101023 115841 101051
rect 115869 101023 115904 101051
rect 115744 100989 115904 101023
rect 115744 100961 115779 100989
rect 115807 100961 115841 100989
rect 115869 100961 115904 100989
rect 115744 100944 115904 100961
rect 125589 101175 125899 109961
rect 125589 101147 125637 101175
rect 125665 101147 125699 101175
rect 125727 101147 125761 101175
rect 125789 101147 125823 101175
rect 125851 101147 125899 101175
rect 125589 101113 125899 101147
rect 125589 101085 125637 101113
rect 125665 101085 125699 101113
rect 125727 101085 125761 101113
rect 125789 101085 125823 101113
rect 125851 101085 125899 101113
rect 125589 101051 125899 101085
rect 125589 101023 125637 101051
rect 125665 101023 125699 101051
rect 125727 101023 125761 101051
rect 125789 101023 125823 101051
rect 125851 101023 125899 101051
rect 125589 100989 125899 101023
rect 125589 100961 125637 100989
rect 125665 100961 125699 100989
rect 125727 100961 125761 100989
rect 125789 100961 125823 100989
rect 125851 100961 125899 100989
rect 112089 95147 112137 95175
rect 112165 95147 112199 95175
rect 112227 95147 112261 95175
rect 112289 95147 112323 95175
rect 112351 95147 112399 95175
rect 112089 95113 112399 95147
rect 112089 95085 112137 95113
rect 112165 95085 112199 95113
rect 112227 95085 112261 95113
rect 112289 95085 112323 95113
rect 112351 95085 112399 95113
rect 112089 95051 112399 95085
rect 112089 95023 112137 95051
rect 112165 95023 112199 95051
rect 112227 95023 112261 95051
rect 112289 95023 112323 95051
rect 112351 95023 112399 95051
rect 112089 94989 112399 95023
rect 112089 94961 112137 94989
rect 112165 94961 112199 94989
rect 112227 94961 112261 94989
rect 112289 94961 112323 94989
rect 112351 94961 112399 94989
rect 112089 86175 112399 94961
rect 123424 95175 123584 95192
rect 123424 95147 123459 95175
rect 123487 95147 123521 95175
rect 123549 95147 123584 95175
rect 123424 95113 123584 95147
rect 123424 95085 123459 95113
rect 123487 95085 123521 95113
rect 123549 95085 123584 95113
rect 123424 95051 123584 95085
rect 123424 95023 123459 95051
rect 123487 95023 123521 95051
rect 123549 95023 123584 95051
rect 123424 94989 123584 95023
rect 123424 94961 123459 94989
rect 123487 94961 123521 94989
rect 123549 94961 123584 94989
rect 123424 94944 123584 94961
rect 115744 92175 115904 92192
rect 115744 92147 115779 92175
rect 115807 92147 115841 92175
rect 115869 92147 115904 92175
rect 115744 92113 115904 92147
rect 115744 92085 115779 92113
rect 115807 92085 115841 92113
rect 115869 92085 115904 92113
rect 115744 92051 115904 92085
rect 115744 92023 115779 92051
rect 115807 92023 115841 92051
rect 115869 92023 115904 92051
rect 115744 91989 115904 92023
rect 115744 91961 115779 91989
rect 115807 91961 115841 91989
rect 115869 91961 115904 91989
rect 115744 91944 115904 91961
rect 125589 92175 125899 100961
rect 125589 92147 125637 92175
rect 125665 92147 125699 92175
rect 125727 92147 125761 92175
rect 125789 92147 125823 92175
rect 125851 92147 125899 92175
rect 125589 92113 125899 92147
rect 125589 92085 125637 92113
rect 125665 92085 125699 92113
rect 125727 92085 125761 92113
rect 125789 92085 125823 92113
rect 125851 92085 125899 92113
rect 125589 92051 125899 92085
rect 125589 92023 125637 92051
rect 125665 92023 125699 92051
rect 125727 92023 125761 92051
rect 125789 92023 125823 92051
rect 125851 92023 125899 92051
rect 125589 91989 125899 92023
rect 125589 91961 125637 91989
rect 125665 91961 125699 91989
rect 125727 91961 125761 91989
rect 125789 91961 125823 91989
rect 125851 91961 125899 91989
rect 112089 86147 112137 86175
rect 112165 86147 112199 86175
rect 112227 86147 112261 86175
rect 112289 86147 112323 86175
rect 112351 86147 112399 86175
rect 112089 86113 112399 86147
rect 112089 86085 112137 86113
rect 112165 86085 112199 86113
rect 112227 86085 112261 86113
rect 112289 86085 112323 86113
rect 112351 86085 112399 86113
rect 112089 86051 112399 86085
rect 112089 86023 112137 86051
rect 112165 86023 112199 86051
rect 112227 86023 112261 86051
rect 112289 86023 112323 86051
rect 112351 86023 112399 86051
rect 112089 85989 112399 86023
rect 112089 85961 112137 85989
rect 112165 85961 112199 85989
rect 112227 85961 112261 85989
rect 112289 85961 112323 85989
rect 112351 85961 112399 85989
rect 112089 77175 112399 85961
rect 123424 86175 123584 86192
rect 123424 86147 123459 86175
rect 123487 86147 123521 86175
rect 123549 86147 123584 86175
rect 123424 86113 123584 86147
rect 123424 86085 123459 86113
rect 123487 86085 123521 86113
rect 123549 86085 123584 86113
rect 123424 86051 123584 86085
rect 123424 86023 123459 86051
rect 123487 86023 123521 86051
rect 123549 86023 123584 86051
rect 123424 85989 123584 86023
rect 123424 85961 123459 85989
rect 123487 85961 123521 85989
rect 123549 85961 123584 85989
rect 123424 85944 123584 85961
rect 115744 83175 115904 83192
rect 115744 83147 115779 83175
rect 115807 83147 115841 83175
rect 115869 83147 115904 83175
rect 115744 83113 115904 83147
rect 115744 83085 115779 83113
rect 115807 83085 115841 83113
rect 115869 83085 115904 83113
rect 115744 83051 115904 83085
rect 115744 83023 115779 83051
rect 115807 83023 115841 83051
rect 115869 83023 115904 83051
rect 115744 82989 115904 83023
rect 115744 82961 115779 82989
rect 115807 82961 115841 82989
rect 115869 82961 115904 82989
rect 115744 82944 115904 82961
rect 125589 83175 125899 91961
rect 125589 83147 125637 83175
rect 125665 83147 125699 83175
rect 125727 83147 125761 83175
rect 125789 83147 125823 83175
rect 125851 83147 125899 83175
rect 125589 83113 125899 83147
rect 125589 83085 125637 83113
rect 125665 83085 125699 83113
rect 125727 83085 125761 83113
rect 125789 83085 125823 83113
rect 125851 83085 125899 83113
rect 125589 83051 125899 83085
rect 125589 83023 125637 83051
rect 125665 83023 125699 83051
rect 125727 83023 125761 83051
rect 125789 83023 125823 83051
rect 125851 83023 125899 83051
rect 125589 82989 125899 83023
rect 125589 82961 125637 82989
rect 125665 82961 125699 82989
rect 125727 82961 125761 82989
rect 125789 82961 125823 82989
rect 125851 82961 125899 82989
rect 112089 77147 112137 77175
rect 112165 77147 112199 77175
rect 112227 77147 112261 77175
rect 112289 77147 112323 77175
rect 112351 77147 112399 77175
rect 112089 77113 112399 77147
rect 112089 77085 112137 77113
rect 112165 77085 112199 77113
rect 112227 77085 112261 77113
rect 112289 77085 112323 77113
rect 112351 77085 112399 77113
rect 112089 77051 112399 77085
rect 112089 77023 112137 77051
rect 112165 77023 112199 77051
rect 112227 77023 112261 77051
rect 112289 77023 112323 77051
rect 112351 77023 112399 77051
rect 112089 76989 112399 77023
rect 112089 76961 112137 76989
rect 112165 76961 112199 76989
rect 112227 76961 112261 76989
rect 112289 76961 112323 76989
rect 112351 76961 112399 76989
rect 112089 68175 112399 76961
rect 123424 77175 123584 77192
rect 123424 77147 123459 77175
rect 123487 77147 123521 77175
rect 123549 77147 123584 77175
rect 123424 77113 123584 77147
rect 123424 77085 123459 77113
rect 123487 77085 123521 77113
rect 123549 77085 123584 77113
rect 123424 77051 123584 77085
rect 123424 77023 123459 77051
rect 123487 77023 123521 77051
rect 123549 77023 123584 77051
rect 123424 76989 123584 77023
rect 123424 76961 123459 76989
rect 123487 76961 123521 76989
rect 123549 76961 123584 76989
rect 123424 76944 123584 76961
rect 115744 74175 115904 74192
rect 115744 74147 115779 74175
rect 115807 74147 115841 74175
rect 115869 74147 115904 74175
rect 115744 74113 115904 74147
rect 115744 74085 115779 74113
rect 115807 74085 115841 74113
rect 115869 74085 115904 74113
rect 115744 74051 115904 74085
rect 115744 74023 115779 74051
rect 115807 74023 115841 74051
rect 115869 74023 115904 74051
rect 115744 73989 115904 74023
rect 115744 73961 115779 73989
rect 115807 73961 115841 73989
rect 115869 73961 115904 73989
rect 115744 73944 115904 73961
rect 125589 74175 125899 82961
rect 125589 74147 125637 74175
rect 125665 74147 125699 74175
rect 125727 74147 125761 74175
rect 125789 74147 125823 74175
rect 125851 74147 125899 74175
rect 125589 74113 125899 74147
rect 125589 74085 125637 74113
rect 125665 74085 125699 74113
rect 125727 74085 125761 74113
rect 125789 74085 125823 74113
rect 125851 74085 125899 74113
rect 125589 74051 125899 74085
rect 125589 74023 125637 74051
rect 125665 74023 125699 74051
rect 125727 74023 125761 74051
rect 125789 74023 125823 74051
rect 125851 74023 125899 74051
rect 125589 73989 125899 74023
rect 125589 73961 125637 73989
rect 125665 73961 125699 73989
rect 125727 73961 125761 73989
rect 125789 73961 125823 73989
rect 125851 73961 125899 73989
rect 112089 68147 112137 68175
rect 112165 68147 112199 68175
rect 112227 68147 112261 68175
rect 112289 68147 112323 68175
rect 112351 68147 112399 68175
rect 112089 68113 112399 68147
rect 112089 68085 112137 68113
rect 112165 68085 112199 68113
rect 112227 68085 112261 68113
rect 112289 68085 112323 68113
rect 112351 68085 112399 68113
rect 112089 68051 112399 68085
rect 112089 68023 112137 68051
rect 112165 68023 112199 68051
rect 112227 68023 112261 68051
rect 112289 68023 112323 68051
rect 112351 68023 112399 68051
rect 112089 67989 112399 68023
rect 112089 67961 112137 67989
rect 112165 67961 112199 67989
rect 112227 67961 112261 67989
rect 112289 67961 112323 67989
rect 112351 67961 112399 67989
rect 112089 59175 112399 67961
rect 123424 68175 123584 68192
rect 123424 68147 123459 68175
rect 123487 68147 123521 68175
rect 123549 68147 123584 68175
rect 123424 68113 123584 68147
rect 123424 68085 123459 68113
rect 123487 68085 123521 68113
rect 123549 68085 123584 68113
rect 123424 68051 123584 68085
rect 123424 68023 123459 68051
rect 123487 68023 123521 68051
rect 123549 68023 123584 68051
rect 123424 67989 123584 68023
rect 123424 67961 123459 67989
rect 123487 67961 123521 67989
rect 123549 67961 123584 67989
rect 123424 67944 123584 67961
rect 115744 65175 115904 65192
rect 115744 65147 115779 65175
rect 115807 65147 115841 65175
rect 115869 65147 115904 65175
rect 115744 65113 115904 65147
rect 115744 65085 115779 65113
rect 115807 65085 115841 65113
rect 115869 65085 115904 65113
rect 115744 65051 115904 65085
rect 115744 65023 115779 65051
rect 115807 65023 115841 65051
rect 115869 65023 115904 65051
rect 115744 64989 115904 65023
rect 115744 64961 115779 64989
rect 115807 64961 115841 64989
rect 115869 64961 115904 64989
rect 115744 64944 115904 64961
rect 125589 65175 125899 73961
rect 125589 65147 125637 65175
rect 125665 65147 125699 65175
rect 125727 65147 125761 65175
rect 125789 65147 125823 65175
rect 125851 65147 125899 65175
rect 125589 65113 125899 65147
rect 125589 65085 125637 65113
rect 125665 65085 125699 65113
rect 125727 65085 125761 65113
rect 125789 65085 125823 65113
rect 125851 65085 125899 65113
rect 125589 65051 125899 65085
rect 125589 65023 125637 65051
rect 125665 65023 125699 65051
rect 125727 65023 125761 65051
rect 125789 65023 125823 65051
rect 125851 65023 125899 65051
rect 125589 64989 125899 65023
rect 125589 64961 125637 64989
rect 125665 64961 125699 64989
rect 125727 64961 125761 64989
rect 125789 64961 125823 64989
rect 125851 64961 125899 64989
rect 112089 59147 112137 59175
rect 112165 59147 112199 59175
rect 112227 59147 112261 59175
rect 112289 59147 112323 59175
rect 112351 59147 112399 59175
rect 112089 59113 112399 59147
rect 112089 59085 112137 59113
rect 112165 59085 112199 59113
rect 112227 59085 112261 59113
rect 112289 59085 112323 59113
rect 112351 59085 112399 59113
rect 112089 59051 112399 59085
rect 112089 59023 112137 59051
rect 112165 59023 112199 59051
rect 112227 59023 112261 59051
rect 112289 59023 112323 59051
rect 112351 59023 112399 59051
rect 112089 58989 112399 59023
rect 112089 58961 112137 58989
rect 112165 58961 112199 58989
rect 112227 58961 112261 58989
rect 112289 58961 112323 58989
rect 112351 58961 112399 58989
rect 112089 50175 112399 58961
rect 123424 59175 123584 59192
rect 123424 59147 123459 59175
rect 123487 59147 123521 59175
rect 123549 59147 123584 59175
rect 123424 59113 123584 59147
rect 123424 59085 123459 59113
rect 123487 59085 123521 59113
rect 123549 59085 123584 59113
rect 123424 59051 123584 59085
rect 123424 59023 123459 59051
rect 123487 59023 123521 59051
rect 123549 59023 123584 59051
rect 123424 58989 123584 59023
rect 123424 58961 123459 58989
rect 123487 58961 123521 58989
rect 123549 58961 123584 58989
rect 123424 58944 123584 58961
rect 115744 56175 115904 56192
rect 115744 56147 115779 56175
rect 115807 56147 115841 56175
rect 115869 56147 115904 56175
rect 115744 56113 115904 56147
rect 115744 56085 115779 56113
rect 115807 56085 115841 56113
rect 115869 56085 115904 56113
rect 115744 56051 115904 56085
rect 115744 56023 115779 56051
rect 115807 56023 115841 56051
rect 115869 56023 115904 56051
rect 115744 55989 115904 56023
rect 115744 55961 115779 55989
rect 115807 55961 115841 55989
rect 115869 55961 115904 55989
rect 115744 55944 115904 55961
rect 125589 56175 125899 64961
rect 125589 56147 125637 56175
rect 125665 56147 125699 56175
rect 125727 56147 125761 56175
rect 125789 56147 125823 56175
rect 125851 56147 125899 56175
rect 125589 56113 125899 56147
rect 125589 56085 125637 56113
rect 125665 56085 125699 56113
rect 125727 56085 125761 56113
rect 125789 56085 125823 56113
rect 125851 56085 125899 56113
rect 125589 56051 125899 56085
rect 125589 56023 125637 56051
rect 125665 56023 125699 56051
rect 125727 56023 125761 56051
rect 125789 56023 125823 56051
rect 125851 56023 125899 56051
rect 125589 55989 125899 56023
rect 125589 55961 125637 55989
rect 125665 55961 125699 55989
rect 125727 55961 125761 55989
rect 125789 55961 125823 55989
rect 125851 55961 125899 55989
rect 112089 50147 112137 50175
rect 112165 50147 112199 50175
rect 112227 50147 112261 50175
rect 112289 50147 112323 50175
rect 112351 50147 112399 50175
rect 112089 50113 112399 50147
rect 112089 50085 112137 50113
rect 112165 50085 112199 50113
rect 112227 50085 112261 50113
rect 112289 50085 112323 50113
rect 112351 50085 112399 50113
rect 112089 50051 112399 50085
rect 112089 50023 112137 50051
rect 112165 50023 112199 50051
rect 112227 50023 112261 50051
rect 112289 50023 112323 50051
rect 112351 50023 112399 50051
rect 112089 49989 112399 50023
rect 112089 49961 112137 49989
rect 112165 49961 112199 49989
rect 112227 49961 112261 49989
rect 112289 49961 112323 49989
rect 112351 49961 112399 49989
rect 112089 41175 112399 49961
rect 123424 50175 123584 50192
rect 123424 50147 123459 50175
rect 123487 50147 123521 50175
rect 123549 50147 123584 50175
rect 123424 50113 123584 50147
rect 123424 50085 123459 50113
rect 123487 50085 123521 50113
rect 123549 50085 123584 50113
rect 123424 50051 123584 50085
rect 123424 50023 123459 50051
rect 123487 50023 123521 50051
rect 123549 50023 123584 50051
rect 123424 49989 123584 50023
rect 123424 49961 123459 49989
rect 123487 49961 123521 49989
rect 123549 49961 123584 49989
rect 123424 49944 123584 49961
rect 115744 47175 115904 47192
rect 115744 47147 115779 47175
rect 115807 47147 115841 47175
rect 115869 47147 115904 47175
rect 115744 47113 115904 47147
rect 115744 47085 115779 47113
rect 115807 47085 115841 47113
rect 115869 47085 115904 47113
rect 115744 47051 115904 47085
rect 115744 47023 115779 47051
rect 115807 47023 115841 47051
rect 115869 47023 115904 47051
rect 115744 46989 115904 47023
rect 115744 46961 115779 46989
rect 115807 46961 115841 46989
rect 115869 46961 115904 46989
rect 115744 46944 115904 46961
rect 125589 47175 125899 55961
rect 125589 47147 125637 47175
rect 125665 47147 125699 47175
rect 125727 47147 125761 47175
rect 125789 47147 125823 47175
rect 125851 47147 125899 47175
rect 125589 47113 125899 47147
rect 125589 47085 125637 47113
rect 125665 47085 125699 47113
rect 125727 47085 125761 47113
rect 125789 47085 125823 47113
rect 125851 47085 125899 47113
rect 125589 47051 125899 47085
rect 125589 47023 125637 47051
rect 125665 47023 125699 47051
rect 125727 47023 125761 47051
rect 125789 47023 125823 47051
rect 125851 47023 125899 47051
rect 125589 46989 125899 47023
rect 125589 46961 125637 46989
rect 125665 46961 125699 46989
rect 125727 46961 125761 46989
rect 125789 46961 125823 46989
rect 125851 46961 125899 46989
rect 112089 41147 112137 41175
rect 112165 41147 112199 41175
rect 112227 41147 112261 41175
rect 112289 41147 112323 41175
rect 112351 41147 112399 41175
rect 112089 41113 112399 41147
rect 112089 41085 112137 41113
rect 112165 41085 112199 41113
rect 112227 41085 112261 41113
rect 112289 41085 112323 41113
rect 112351 41085 112399 41113
rect 112089 41051 112399 41085
rect 112089 41023 112137 41051
rect 112165 41023 112199 41051
rect 112227 41023 112261 41051
rect 112289 41023 112323 41051
rect 112351 41023 112399 41051
rect 112089 40989 112399 41023
rect 112089 40961 112137 40989
rect 112165 40961 112199 40989
rect 112227 40961 112261 40989
rect 112289 40961 112323 40989
rect 112351 40961 112399 40989
rect 112089 32175 112399 40961
rect 123424 41175 123584 41192
rect 123424 41147 123459 41175
rect 123487 41147 123521 41175
rect 123549 41147 123584 41175
rect 123424 41113 123584 41147
rect 123424 41085 123459 41113
rect 123487 41085 123521 41113
rect 123549 41085 123584 41113
rect 123424 41051 123584 41085
rect 123424 41023 123459 41051
rect 123487 41023 123521 41051
rect 123549 41023 123584 41051
rect 123424 40989 123584 41023
rect 123424 40961 123459 40989
rect 123487 40961 123521 40989
rect 123549 40961 123584 40989
rect 123424 40944 123584 40961
rect 115744 38175 115904 38192
rect 115744 38147 115779 38175
rect 115807 38147 115841 38175
rect 115869 38147 115904 38175
rect 115744 38113 115904 38147
rect 115744 38085 115779 38113
rect 115807 38085 115841 38113
rect 115869 38085 115904 38113
rect 115744 38051 115904 38085
rect 115744 38023 115779 38051
rect 115807 38023 115841 38051
rect 115869 38023 115904 38051
rect 115744 37989 115904 38023
rect 115744 37961 115779 37989
rect 115807 37961 115841 37989
rect 115869 37961 115904 37989
rect 115744 37944 115904 37961
rect 125589 38175 125899 46961
rect 125589 38147 125637 38175
rect 125665 38147 125699 38175
rect 125727 38147 125761 38175
rect 125789 38147 125823 38175
rect 125851 38147 125899 38175
rect 125589 38113 125899 38147
rect 125589 38085 125637 38113
rect 125665 38085 125699 38113
rect 125727 38085 125761 38113
rect 125789 38085 125823 38113
rect 125851 38085 125899 38113
rect 125589 38051 125899 38085
rect 125589 38023 125637 38051
rect 125665 38023 125699 38051
rect 125727 38023 125761 38051
rect 125789 38023 125823 38051
rect 125851 38023 125899 38051
rect 125589 37989 125899 38023
rect 125589 37961 125637 37989
rect 125665 37961 125699 37989
rect 125727 37961 125761 37989
rect 125789 37961 125823 37989
rect 125851 37961 125899 37989
rect 112089 32147 112137 32175
rect 112165 32147 112199 32175
rect 112227 32147 112261 32175
rect 112289 32147 112323 32175
rect 112351 32147 112399 32175
rect 112089 32113 112399 32147
rect 112089 32085 112137 32113
rect 112165 32085 112199 32113
rect 112227 32085 112261 32113
rect 112289 32085 112323 32113
rect 112351 32085 112399 32113
rect 112089 32051 112399 32085
rect 112089 32023 112137 32051
rect 112165 32023 112199 32051
rect 112227 32023 112261 32051
rect 112289 32023 112323 32051
rect 112351 32023 112399 32051
rect 112089 31989 112399 32023
rect 112089 31961 112137 31989
rect 112165 31961 112199 31989
rect 112227 31961 112261 31989
rect 112289 31961 112323 31989
rect 112351 31961 112399 31989
rect 112089 23175 112399 31961
rect 123424 32175 123584 32192
rect 123424 32147 123459 32175
rect 123487 32147 123521 32175
rect 123549 32147 123584 32175
rect 123424 32113 123584 32147
rect 123424 32085 123459 32113
rect 123487 32085 123521 32113
rect 123549 32085 123584 32113
rect 123424 32051 123584 32085
rect 123424 32023 123459 32051
rect 123487 32023 123521 32051
rect 123549 32023 123584 32051
rect 123424 31989 123584 32023
rect 123424 31961 123459 31989
rect 123487 31961 123521 31989
rect 123549 31961 123584 31989
rect 123424 31944 123584 31961
rect 115744 29175 115904 29192
rect 115744 29147 115779 29175
rect 115807 29147 115841 29175
rect 115869 29147 115904 29175
rect 115744 29113 115904 29147
rect 115744 29085 115779 29113
rect 115807 29085 115841 29113
rect 115869 29085 115904 29113
rect 115744 29051 115904 29085
rect 115744 29023 115779 29051
rect 115807 29023 115841 29051
rect 115869 29023 115904 29051
rect 115744 28989 115904 29023
rect 115744 28961 115779 28989
rect 115807 28961 115841 28989
rect 115869 28961 115904 28989
rect 115744 28944 115904 28961
rect 125589 29175 125899 37961
rect 125589 29147 125637 29175
rect 125665 29147 125699 29175
rect 125727 29147 125761 29175
rect 125789 29147 125823 29175
rect 125851 29147 125899 29175
rect 125589 29113 125899 29147
rect 125589 29085 125637 29113
rect 125665 29085 125699 29113
rect 125727 29085 125761 29113
rect 125789 29085 125823 29113
rect 125851 29085 125899 29113
rect 125589 29051 125899 29085
rect 125589 29023 125637 29051
rect 125665 29023 125699 29051
rect 125727 29023 125761 29051
rect 125789 29023 125823 29051
rect 125851 29023 125899 29051
rect 125589 28989 125899 29023
rect 125589 28961 125637 28989
rect 125665 28961 125699 28989
rect 125727 28961 125761 28989
rect 125789 28961 125823 28989
rect 125851 28961 125899 28989
rect 112089 23147 112137 23175
rect 112165 23147 112199 23175
rect 112227 23147 112261 23175
rect 112289 23147 112323 23175
rect 112351 23147 112399 23175
rect 112089 23113 112399 23147
rect 112089 23085 112137 23113
rect 112165 23085 112199 23113
rect 112227 23085 112261 23113
rect 112289 23085 112323 23113
rect 112351 23085 112399 23113
rect 112089 23051 112399 23085
rect 112089 23023 112137 23051
rect 112165 23023 112199 23051
rect 112227 23023 112261 23051
rect 112289 23023 112323 23051
rect 112351 23023 112399 23051
rect 112089 22989 112399 23023
rect 112089 22961 112137 22989
rect 112165 22961 112199 22989
rect 112227 22961 112261 22989
rect 112289 22961 112323 22989
rect 112351 22961 112399 22989
rect 112089 14175 112399 22961
rect 123424 23175 123584 23192
rect 123424 23147 123459 23175
rect 123487 23147 123521 23175
rect 123549 23147 123584 23175
rect 123424 23113 123584 23147
rect 123424 23085 123459 23113
rect 123487 23085 123521 23113
rect 123549 23085 123584 23113
rect 123424 23051 123584 23085
rect 123424 23023 123459 23051
rect 123487 23023 123521 23051
rect 123549 23023 123584 23051
rect 123424 22989 123584 23023
rect 123424 22961 123459 22989
rect 123487 22961 123521 22989
rect 123549 22961 123584 22989
rect 123424 22944 123584 22961
rect 115744 20175 115904 20192
rect 115744 20147 115779 20175
rect 115807 20147 115841 20175
rect 115869 20147 115904 20175
rect 115744 20113 115904 20147
rect 115744 20085 115779 20113
rect 115807 20085 115841 20113
rect 115869 20085 115904 20113
rect 115744 20051 115904 20085
rect 115744 20023 115779 20051
rect 115807 20023 115841 20051
rect 115869 20023 115904 20051
rect 115744 19989 115904 20023
rect 115744 19961 115779 19989
rect 115807 19961 115841 19989
rect 115869 19961 115904 19989
rect 115744 19944 115904 19961
rect 125589 20175 125899 28961
rect 125589 20147 125637 20175
rect 125665 20147 125699 20175
rect 125727 20147 125761 20175
rect 125789 20147 125823 20175
rect 125851 20147 125899 20175
rect 125589 20113 125899 20147
rect 125589 20085 125637 20113
rect 125665 20085 125699 20113
rect 125727 20085 125761 20113
rect 125789 20085 125823 20113
rect 125851 20085 125899 20113
rect 125589 20051 125899 20085
rect 125589 20023 125637 20051
rect 125665 20023 125699 20051
rect 125727 20023 125761 20051
rect 125789 20023 125823 20051
rect 125851 20023 125899 20051
rect 125589 19989 125899 20023
rect 125589 19961 125637 19989
rect 125665 19961 125699 19989
rect 125727 19961 125761 19989
rect 125789 19961 125823 19989
rect 125851 19961 125899 19989
rect 112089 14147 112137 14175
rect 112165 14147 112199 14175
rect 112227 14147 112261 14175
rect 112289 14147 112323 14175
rect 112351 14147 112399 14175
rect 112089 14113 112399 14147
rect 112089 14085 112137 14113
rect 112165 14085 112199 14113
rect 112227 14085 112261 14113
rect 112289 14085 112323 14113
rect 112351 14085 112399 14113
rect 112089 14051 112399 14085
rect 112089 14023 112137 14051
rect 112165 14023 112199 14051
rect 112227 14023 112261 14051
rect 112289 14023 112323 14051
rect 112351 14023 112399 14051
rect 112089 13989 112399 14023
rect 112089 13961 112137 13989
rect 112165 13961 112199 13989
rect 112227 13961 112261 13989
rect 112289 13961 112323 13989
rect 112351 13961 112399 13989
rect 112089 5175 112399 13961
rect 123424 14175 123584 14192
rect 123424 14147 123459 14175
rect 123487 14147 123521 14175
rect 123549 14147 123584 14175
rect 123424 14113 123584 14147
rect 123424 14085 123459 14113
rect 123487 14085 123521 14113
rect 123549 14085 123584 14113
rect 123424 14051 123584 14085
rect 123424 14023 123459 14051
rect 123487 14023 123521 14051
rect 123549 14023 123584 14051
rect 123424 13989 123584 14023
rect 123424 13961 123459 13989
rect 123487 13961 123521 13989
rect 123549 13961 123584 13989
rect 123424 13944 123584 13961
rect 115744 11175 115904 11192
rect 115744 11147 115779 11175
rect 115807 11147 115841 11175
rect 115869 11147 115904 11175
rect 115744 11113 115904 11147
rect 115744 11085 115779 11113
rect 115807 11085 115841 11113
rect 115869 11085 115904 11113
rect 115744 11051 115904 11085
rect 115744 11023 115779 11051
rect 115807 11023 115841 11051
rect 115869 11023 115904 11051
rect 115744 10989 115904 11023
rect 115744 10961 115779 10989
rect 115807 10961 115841 10989
rect 115869 10961 115904 10989
rect 115744 10944 115904 10961
rect 125589 11175 125899 19961
rect 125589 11147 125637 11175
rect 125665 11147 125699 11175
rect 125727 11147 125761 11175
rect 125789 11147 125823 11175
rect 125851 11147 125899 11175
rect 125589 11113 125899 11147
rect 125589 11085 125637 11113
rect 125665 11085 125699 11113
rect 125727 11085 125761 11113
rect 125789 11085 125823 11113
rect 125851 11085 125899 11113
rect 125589 11051 125899 11085
rect 125589 11023 125637 11051
rect 125665 11023 125699 11051
rect 125727 11023 125761 11051
rect 125789 11023 125823 11051
rect 125851 11023 125899 11051
rect 125589 10989 125899 11023
rect 125589 10961 125637 10989
rect 125665 10961 125699 10989
rect 125727 10961 125761 10989
rect 125789 10961 125823 10989
rect 125851 10961 125899 10989
rect 112089 5147 112137 5175
rect 112165 5147 112199 5175
rect 112227 5147 112261 5175
rect 112289 5147 112323 5175
rect 112351 5147 112399 5175
rect 112089 5113 112399 5147
rect 112089 5085 112137 5113
rect 112165 5085 112199 5113
rect 112227 5085 112261 5113
rect 112289 5085 112323 5113
rect 112351 5085 112399 5113
rect 112089 5051 112399 5085
rect 112089 5023 112137 5051
rect 112165 5023 112199 5051
rect 112227 5023 112261 5051
rect 112289 5023 112323 5051
rect 112351 5023 112399 5051
rect 112089 4989 112399 5023
rect 112089 4961 112137 4989
rect 112165 4961 112199 4989
rect 112227 4961 112261 4989
rect 112289 4961 112323 4989
rect 112351 4961 112399 4989
rect 112089 -560 112399 4961
rect 123424 5175 123584 5192
rect 123424 5147 123459 5175
rect 123487 5147 123521 5175
rect 123549 5147 123584 5175
rect 123424 5113 123584 5147
rect 123424 5085 123459 5113
rect 123487 5085 123521 5113
rect 123549 5085 123584 5113
rect 123424 5051 123584 5085
rect 123424 5023 123459 5051
rect 123487 5023 123521 5051
rect 123549 5023 123584 5051
rect 123424 4989 123584 5023
rect 123424 4961 123459 4989
rect 123487 4961 123521 4989
rect 123549 4961 123584 4989
rect 123424 4944 123584 4961
rect 112089 -588 112137 -560
rect 112165 -588 112199 -560
rect 112227 -588 112261 -560
rect 112289 -588 112323 -560
rect 112351 -588 112399 -560
rect 112089 -622 112399 -588
rect 112089 -650 112137 -622
rect 112165 -650 112199 -622
rect 112227 -650 112261 -622
rect 112289 -650 112323 -622
rect 112351 -650 112399 -622
rect 112089 -684 112399 -650
rect 112089 -712 112137 -684
rect 112165 -712 112199 -684
rect 112227 -712 112261 -684
rect 112289 -712 112323 -684
rect 112351 -712 112399 -684
rect 112089 -746 112399 -712
rect 112089 -774 112137 -746
rect 112165 -774 112199 -746
rect 112227 -774 112261 -746
rect 112289 -774 112323 -746
rect 112351 -774 112399 -746
rect 112089 -822 112399 -774
rect 125589 2175 125899 10961
rect 125589 2147 125637 2175
rect 125665 2147 125699 2175
rect 125727 2147 125761 2175
rect 125789 2147 125823 2175
rect 125851 2147 125899 2175
rect 125589 2113 125899 2147
rect 125589 2085 125637 2113
rect 125665 2085 125699 2113
rect 125727 2085 125761 2113
rect 125789 2085 125823 2113
rect 125851 2085 125899 2113
rect 125589 2051 125899 2085
rect 125589 2023 125637 2051
rect 125665 2023 125699 2051
rect 125727 2023 125761 2051
rect 125789 2023 125823 2051
rect 125851 2023 125899 2051
rect 125589 1989 125899 2023
rect 125589 1961 125637 1989
rect 125665 1961 125699 1989
rect 125727 1961 125761 1989
rect 125789 1961 125823 1989
rect 125851 1961 125899 1989
rect 125589 -80 125899 1961
rect 125589 -108 125637 -80
rect 125665 -108 125699 -80
rect 125727 -108 125761 -80
rect 125789 -108 125823 -80
rect 125851 -108 125899 -80
rect 125589 -142 125899 -108
rect 125589 -170 125637 -142
rect 125665 -170 125699 -142
rect 125727 -170 125761 -142
rect 125789 -170 125823 -142
rect 125851 -170 125899 -142
rect 125589 -204 125899 -170
rect 125589 -232 125637 -204
rect 125665 -232 125699 -204
rect 125727 -232 125761 -204
rect 125789 -232 125823 -204
rect 125851 -232 125899 -204
rect 125589 -266 125899 -232
rect 125589 -294 125637 -266
rect 125665 -294 125699 -266
rect 125727 -294 125761 -266
rect 125789 -294 125823 -266
rect 125851 -294 125899 -266
rect 125589 -822 125899 -294
rect 127449 299086 127759 299134
rect 127449 299058 127497 299086
rect 127525 299058 127559 299086
rect 127587 299058 127621 299086
rect 127649 299058 127683 299086
rect 127711 299058 127759 299086
rect 127449 299024 127759 299058
rect 127449 298996 127497 299024
rect 127525 298996 127559 299024
rect 127587 298996 127621 299024
rect 127649 298996 127683 299024
rect 127711 298996 127759 299024
rect 127449 298962 127759 298996
rect 127449 298934 127497 298962
rect 127525 298934 127559 298962
rect 127587 298934 127621 298962
rect 127649 298934 127683 298962
rect 127711 298934 127759 298962
rect 127449 298900 127759 298934
rect 127449 298872 127497 298900
rect 127525 298872 127559 298900
rect 127587 298872 127621 298900
rect 127649 298872 127683 298900
rect 127711 298872 127759 298900
rect 127449 293175 127759 298872
rect 127449 293147 127497 293175
rect 127525 293147 127559 293175
rect 127587 293147 127621 293175
rect 127649 293147 127683 293175
rect 127711 293147 127759 293175
rect 127449 293113 127759 293147
rect 127449 293085 127497 293113
rect 127525 293085 127559 293113
rect 127587 293085 127621 293113
rect 127649 293085 127683 293113
rect 127711 293085 127759 293113
rect 127449 293051 127759 293085
rect 127449 293023 127497 293051
rect 127525 293023 127559 293051
rect 127587 293023 127621 293051
rect 127649 293023 127683 293051
rect 127711 293023 127759 293051
rect 127449 292989 127759 293023
rect 127449 292961 127497 292989
rect 127525 292961 127559 292989
rect 127587 292961 127621 292989
rect 127649 292961 127683 292989
rect 127711 292961 127759 292989
rect 127449 284175 127759 292961
rect 127449 284147 127497 284175
rect 127525 284147 127559 284175
rect 127587 284147 127621 284175
rect 127649 284147 127683 284175
rect 127711 284147 127759 284175
rect 127449 284113 127759 284147
rect 127449 284085 127497 284113
rect 127525 284085 127559 284113
rect 127587 284085 127621 284113
rect 127649 284085 127683 284113
rect 127711 284085 127759 284113
rect 127449 284051 127759 284085
rect 127449 284023 127497 284051
rect 127525 284023 127559 284051
rect 127587 284023 127621 284051
rect 127649 284023 127683 284051
rect 127711 284023 127759 284051
rect 127449 283989 127759 284023
rect 127449 283961 127497 283989
rect 127525 283961 127559 283989
rect 127587 283961 127621 283989
rect 127649 283961 127683 283989
rect 127711 283961 127759 283989
rect 127449 275175 127759 283961
rect 127449 275147 127497 275175
rect 127525 275147 127559 275175
rect 127587 275147 127621 275175
rect 127649 275147 127683 275175
rect 127711 275147 127759 275175
rect 127449 275113 127759 275147
rect 127449 275085 127497 275113
rect 127525 275085 127559 275113
rect 127587 275085 127621 275113
rect 127649 275085 127683 275113
rect 127711 275085 127759 275113
rect 127449 275051 127759 275085
rect 127449 275023 127497 275051
rect 127525 275023 127559 275051
rect 127587 275023 127621 275051
rect 127649 275023 127683 275051
rect 127711 275023 127759 275051
rect 127449 274989 127759 275023
rect 127449 274961 127497 274989
rect 127525 274961 127559 274989
rect 127587 274961 127621 274989
rect 127649 274961 127683 274989
rect 127711 274961 127759 274989
rect 127449 266175 127759 274961
rect 127449 266147 127497 266175
rect 127525 266147 127559 266175
rect 127587 266147 127621 266175
rect 127649 266147 127683 266175
rect 127711 266147 127759 266175
rect 127449 266113 127759 266147
rect 127449 266085 127497 266113
rect 127525 266085 127559 266113
rect 127587 266085 127621 266113
rect 127649 266085 127683 266113
rect 127711 266085 127759 266113
rect 127449 266051 127759 266085
rect 127449 266023 127497 266051
rect 127525 266023 127559 266051
rect 127587 266023 127621 266051
rect 127649 266023 127683 266051
rect 127711 266023 127759 266051
rect 127449 265989 127759 266023
rect 127449 265961 127497 265989
rect 127525 265961 127559 265989
rect 127587 265961 127621 265989
rect 127649 265961 127683 265989
rect 127711 265961 127759 265989
rect 127449 257175 127759 265961
rect 127449 257147 127497 257175
rect 127525 257147 127559 257175
rect 127587 257147 127621 257175
rect 127649 257147 127683 257175
rect 127711 257147 127759 257175
rect 127449 257113 127759 257147
rect 127449 257085 127497 257113
rect 127525 257085 127559 257113
rect 127587 257085 127621 257113
rect 127649 257085 127683 257113
rect 127711 257085 127759 257113
rect 127449 257051 127759 257085
rect 127449 257023 127497 257051
rect 127525 257023 127559 257051
rect 127587 257023 127621 257051
rect 127649 257023 127683 257051
rect 127711 257023 127759 257051
rect 127449 256989 127759 257023
rect 127449 256961 127497 256989
rect 127525 256961 127559 256989
rect 127587 256961 127621 256989
rect 127649 256961 127683 256989
rect 127711 256961 127759 256989
rect 127449 248175 127759 256961
rect 127449 248147 127497 248175
rect 127525 248147 127559 248175
rect 127587 248147 127621 248175
rect 127649 248147 127683 248175
rect 127711 248147 127759 248175
rect 127449 248113 127759 248147
rect 127449 248085 127497 248113
rect 127525 248085 127559 248113
rect 127587 248085 127621 248113
rect 127649 248085 127683 248113
rect 127711 248085 127759 248113
rect 127449 248051 127759 248085
rect 127449 248023 127497 248051
rect 127525 248023 127559 248051
rect 127587 248023 127621 248051
rect 127649 248023 127683 248051
rect 127711 248023 127759 248051
rect 127449 247989 127759 248023
rect 127449 247961 127497 247989
rect 127525 247961 127559 247989
rect 127587 247961 127621 247989
rect 127649 247961 127683 247989
rect 127711 247961 127759 247989
rect 127449 239175 127759 247961
rect 127449 239147 127497 239175
rect 127525 239147 127559 239175
rect 127587 239147 127621 239175
rect 127649 239147 127683 239175
rect 127711 239147 127759 239175
rect 127449 239113 127759 239147
rect 127449 239085 127497 239113
rect 127525 239085 127559 239113
rect 127587 239085 127621 239113
rect 127649 239085 127683 239113
rect 127711 239085 127759 239113
rect 127449 239051 127759 239085
rect 127449 239023 127497 239051
rect 127525 239023 127559 239051
rect 127587 239023 127621 239051
rect 127649 239023 127683 239051
rect 127711 239023 127759 239051
rect 127449 238989 127759 239023
rect 127449 238961 127497 238989
rect 127525 238961 127559 238989
rect 127587 238961 127621 238989
rect 127649 238961 127683 238989
rect 127711 238961 127759 238989
rect 127449 230175 127759 238961
rect 127449 230147 127497 230175
rect 127525 230147 127559 230175
rect 127587 230147 127621 230175
rect 127649 230147 127683 230175
rect 127711 230147 127759 230175
rect 127449 230113 127759 230147
rect 127449 230085 127497 230113
rect 127525 230085 127559 230113
rect 127587 230085 127621 230113
rect 127649 230085 127683 230113
rect 127711 230085 127759 230113
rect 127449 230051 127759 230085
rect 127449 230023 127497 230051
rect 127525 230023 127559 230051
rect 127587 230023 127621 230051
rect 127649 230023 127683 230051
rect 127711 230023 127759 230051
rect 127449 229989 127759 230023
rect 127449 229961 127497 229989
rect 127525 229961 127559 229989
rect 127587 229961 127621 229989
rect 127649 229961 127683 229989
rect 127711 229961 127759 229989
rect 127449 221175 127759 229961
rect 127449 221147 127497 221175
rect 127525 221147 127559 221175
rect 127587 221147 127621 221175
rect 127649 221147 127683 221175
rect 127711 221147 127759 221175
rect 127449 221113 127759 221147
rect 127449 221085 127497 221113
rect 127525 221085 127559 221113
rect 127587 221085 127621 221113
rect 127649 221085 127683 221113
rect 127711 221085 127759 221113
rect 127449 221051 127759 221085
rect 127449 221023 127497 221051
rect 127525 221023 127559 221051
rect 127587 221023 127621 221051
rect 127649 221023 127683 221051
rect 127711 221023 127759 221051
rect 127449 220989 127759 221023
rect 127449 220961 127497 220989
rect 127525 220961 127559 220989
rect 127587 220961 127621 220989
rect 127649 220961 127683 220989
rect 127711 220961 127759 220989
rect 127449 212175 127759 220961
rect 127449 212147 127497 212175
rect 127525 212147 127559 212175
rect 127587 212147 127621 212175
rect 127649 212147 127683 212175
rect 127711 212147 127759 212175
rect 127449 212113 127759 212147
rect 127449 212085 127497 212113
rect 127525 212085 127559 212113
rect 127587 212085 127621 212113
rect 127649 212085 127683 212113
rect 127711 212085 127759 212113
rect 127449 212051 127759 212085
rect 127449 212023 127497 212051
rect 127525 212023 127559 212051
rect 127587 212023 127621 212051
rect 127649 212023 127683 212051
rect 127711 212023 127759 212051
rect 127449 211989 127759 212023
rect 127449 211961 127497 211989
rect 127525 211961 127559 211989
rect 127587 211961 127621 211989
rect 127649 211961 127683 211989
rect 127711 211961 127759 211989
rect 127449 203175 127759 211961
rect 127449 203147 127497 203175
rect 127525 203147 127559 203175
rect 127587 203147 127621 203175
rect 127649 203147 127683 203175
rect 127711 203147 127759 203175
rect 127449 203113 127759 203147
rect 127449 203085 127497 203113
rect 127525 203085 127559 203113
rect 127587 203085 127621 203113
rect 127649 203085 127683 203113
rect 127711 203085 127759 203113
rect 127449 203051 127759 203085
rect 127449 203023 127497 203051
rect 127525 203023 127559 203051
rect 127587 203023 127621 203051
rect 127649 203023 127683 203051
rect 127711 203023 127759 203051
rect 127449 202989 127759 203023
rect 127449 202961 127497 202989
rect 127525 202961 127559 202989
rect 127587 202961 127621 202989
rect 127649 202961 127683 202989
rect 127711 202961 127759 202989
rect 127449 194175 127759 202961
rect 127449 194147 127497 194175
rect 127525 194147 127559 194175
rect 127587 194147 127621 194175
rect 127649 194147 127683 194175
rect 127711 194147 127759 194175
rect 127449 194113 127759 194147
rect 127449 194085 127497 194113
rect 127525 194085 127559 194113
rect 127587 194085 127621 194113
rect 127649 194085 127683 194113
rect 127711 194085 127759 194113
rect 127449 194051 127759 194085
rect 127449 194023 127497 194051
rect 127525 194023 127559 194051
rect 127587 194023 127621 194051
rect 127649 194023 127683 194051
rect 127711 194023 127759 194051
rect 127449 193989 127759 194023
rect 127449 193961 127497 193989
rect 127525 193961 127559 193989
rect 127587 193961 127621 193989
rect 127649 193961 127683 193989
rect 127711 193961 127759 193989
rect 127449 185175 127759 193961
rect 127449 185147 127497 185175
rect 127525 185147 127559 185175
rect 127587 185147 127621 185175
rect 127649 185147 127683 185175
rect 127711 185147 127759 185175
rect 127449 185113 127759 185147
rect 127449 185085 127497 185113
rect 127525 185085 127559 185113
rect 127587 185085 127621 185113
rect 127649 185085 127683 185113
rect 127711 185085 127759 185113
rect 127449 185051 127759 185085
rect 127449 185023 127497 185051
rect 127525 185023 127559 185051
rect 127587 185023 127621 185051
rect 127649 185023 127683 185051
rect 127711 185023 127759 185051
rect 127449 184989 127759 185023
rect 127449 184961 127497 184989
rect 127525 184961 127559 184989
rect 127587 184961 127621 184989
rect 127649 184961 127683 184989
rect 127711 184961 127759 184989
rect 127449 176175 127759 184961
rect 127449 176147 127497 176175
rect 127525 176147 127559 176175
rect 127587 176147 127621 176175
rect 127649 176147 127683 176175
rect 127711 176147 127759 176175
rect 127449 176113 127759 176147
rect 127449 176085 127497 176113
rect 127525 176085 127559 176113
rect 127587 176085 127621 176113
rect 127649 176085 127683 176113
rect 127711 176085 127759 176113
rect 127449 176051 127759 176085
rect 127449 176023 127497 176051
rect 127525 176023 127559 176051
rect 127587 176023 127621 176051
rect 127649 176023 127683 176051
rect 127711 176023 127759 176051
rect 127449 175989 127759 176023
rect 127449 175961 127497 175989
rect 127525 175961 127559 175989
rect 127587 175961 127621 175989
rect 127649 175961 127683 175989
rect 127711 175961 127759 175989
rect 127449 167175 127759 175961
rect 140949 298606 141259 299134
rect 140949 298578 140997 298606
rect 141025 298578 141059 298606
rect 141087 298578 141121 298606
rect 141149 298578 141183 298606
rect 141211 298578 141259 298606
rect 140949 298544 141259 298578
rect 140949 298516 140997 298544
rect 141025 298516 141059 298544
rect 141087 298516 141121 298544
rect 141149 298516 141183 298544
rect 141211 298516 141259 298544
rect 140949 298482 141259 298516
rect 140949 298454 140997 298482
rect 141025 298454 141059 298482
rect 141087 298454 141121 298482
rect 141149 298454 141183 298482
rect 141211 298454 141259 298482
rect 140949 298420 141259 298454
rect 140949 298392 140997 298420
rect 141025 298392 141059 298420
rect 141087 298392 141121 298420
rect 141149 298392 141183 298420
rect 141211 298392 141259 298420
rect 140949 290175 141259 298392
rect 140949 290147 140997 290175
rect 141025 290147 141059 290175
rect 141087 290147 141121 290175
rect 141149 290147 141183 290175
rect 141211 290147 141259 290175
rect 140949 290113 141259 290147
rect 140949 290085 140997 290113
rect 141025 290085 141059 290113
rect 141087 290085 141121 290113
rect 141149 290085 141183 290113
rect 141211 290085 141259 290113
rect 140949 290051 141259 290085
rect 140949 290023 140997 290051
rect 141025 290023 141059 290051
rect 141087 290023 141121 290051
rect 141149 290023 141183 290051
rect 141211 290023 141259 290051
rect 140949 289989 141259 290023
rect 140949 289961 140997 289989
rect 141025 289961 141059 289989
rect 141087 289961 141121 289989
rect 141149 289961 141183 289989
rect 141211 289961 141259 289989
rect 140949 281175 141259 289961
rect 140949 281147 140997 281175
rect 141025 281147 141059 281175
rect 141087 281147 141121 281175
rect 141149 281147 141183 281175
rect 141211 281147 141259 281175
rect 140949 281113 141259 281147
rect 140949 281085 140997 281113
rect 141025 281085 141059 281113
rect 141087 281085 141121 281113
rect 141149 281085 141183 281113
rect 141211 281085 141259 281113
rect 140949 281051 141259 281085
rect 140949 281023 140997 281051
rect 141025 281023 141059 281051
rect 141087 281023 141121 281051
rect 141149 281023 141183 281051
rect 141211 281023 141259 281051
rect 140949 280989 141259 281023
rect 140949 280961 140997 280989
rect 141025 280961 141059 280989
rect 141087 280961 141121 280989
rect 141149 280961 141183 280989
rect 141211 280961 141259 280989
rect 140949 272175 141259 280961
rect 140949 272147 140997 272175
rect 141025 272147 141059 272175
rect 141087 272147 141121 272175
rect 141149 272147 141183 272175
rect 141211 272147 141259 272175
rect 140949 272113 141259 272147
rect 140949 272085 140997 272113
rect 141025 272085 141059 272113
rect 141087 272085 141121 272113
rect 141149 272085 141183 272113
rect 141211 272085 141259 272113
rect 140949 272051 141259 272085
rect 140949 272023 140997 272051
rect 141025 272023 141059 272051
rect 141087 272023 141121 272051
rect 141149 272023 141183 272051
rect 141211 272023 141259 272051
rect 140949 271989 141259 272023
rect 140949 271961 140997 271989
rect 141025 271961 141059 271989
rect 141087 271961 141121 271989
rect 141149 271961 141183 271989
rect 141211 271961 141259 271989
rect 140949 263175 141259 271961
rect 140949 263147 140997 263175
rect 141025 263147 141059 263175
rect 141087 263147 141121 263175
rect 141149 263147 141183 263175
rect 141211 263147 141259 263175
rect 140949 263113 141259 263147
rect 140949 263085 140997 263113
rect 141025 263085 141059 263113
rect 141087 263085 141121 263113
rect 141149 263085 141183 263113
rect 141211 263085 141259 263113
rect 140949 263051 141259 263085
rect 140949 263023 140997 263051
rect 141025 263023 141059 263051
rect 141087 263023 141121 263051
rect 141149 263023 141183 263051
rect 141211 263023 141259 263051
rect 140949 262989 141259 263023
rect 140949 262961 140997 262989
rect 141025 262961 141059 262989
rect 141087 262961 141121 262989
rect 141149 262961 141183 262989
rect 141211 262961 141259 262989
rect 140949 254175 141259 262961
rect 140949 254147 140997 254175
rect 141025 254147 141059 254175
rect 141087 254147 141121 254175
rect 141149 254147 141183 254175
rect 141211 254147 141259 254175
rect 140949 254113 141259 254147
rect 140949 254085 140997 254113
rect 141025 254085 141059 254113
rect 141087 254085 141121 254113
rect 141149 254085 141183 254113
rect 141211 254085 141259 254113
rect 140949 254051 141259 254085
rect 140949 254023 140997 254051
rect 141025 254023 141059 254051
rect 141087 254023 141121 254051
rect 141149 254023 141183 254051
rect 141211 254023 141259 254051
rect 140949 253989 141259 254023
rect 140949 253961 140997 253989
rect 141025 253961 141059 253989
rect 141087 253961 141121 253989
rect 141149 253961 141183 253989
rect 141211 253961 141259 253989
rect 140949 245175 141259 253961
rect 140949 245147 140997 245175
rect 141025 245147 141059 245175
rect 141087 245147 141121 245175
rect 141149 245147 141183 245175
rect 141211 245147 141259 245175
rect 140949 245113 141259 245147
rect 140949 245085 140997 245113
rect 141025 245085 141059 245113
rect 141087 245085 141121 245113
rect 141149 245085 141183 245113
rect 141211 245085 141259 245113
rect 140949 245051 141259 245085
rect 140949 245023 140997 245051
rect 141025 245023 141059 245051
rect 141087 245023 141121 245051
rect 141149 245023 141183 245051
rect 141211 245023 141259 245051
rect 140949 244989 141259 245023
rect 140949 244961 140997 244989
rect 141025 244961 141059 244989
rect 141087 244961 141121 244989
rect 141149 244961 141183 244989
rect 141211 244961 141259 244989
rect 140949 236175 141259 244961
rect 140949 236147 140997 236175
rect 141025 236147 141059 236175
rect 141087 236147 141121 236175
rect 141149 236147 141183 236175
rect 141211 236147 141259 236175
rect 140949 236113 141259 236147
rect 140949 236085 140997 236113
rect 141025 236085 141059 236113
rect 141087 236085 141121 236113
rect 141149 236085 141183 236113
rect 141211 236085 141259 236113
rect 140949 236051 141259 236085
rect 140949 236023 140997 236051
rect 141025 236023 141059 236051
rect 141087 236023 141121 236051
rect 141149 236023 141183 236051
rect 141211 236023 141259 236051
rect 140949 235989 141259 236023
rect 140949 235961 140997 235989
rect 141025 235961 141059 235989
rect 141087 235961 141121 235989
rect 141149 235961 141183 235989
rect 141211 235961 141259 235989
rect 140949 227175 141259 235961
rect 140949 227147 140997 227175
rect 141025 227147 141059 227175
rect 141087 227147 141121 227175
rect 141149 227147 141183 227175
rect 141211 227147 141259 227175
rect 140949 227113 141259 227147
rect 140949 227085 140997 227113
rect 141025 227085 141059 227113
rect 141087 227085 141121 227113
rect 141149 227085 141183 227113
rect 141211 227085 141259 227113
rect 140949 227051 141259 227085
rect 140949 227023 140997 227051
rect 141025 227023 141059 227051
rect 141087 227023 141121 227051
rect 141149 227023 141183 227051
rect 141211 227023 141259 227051
rect 140949 226989 141259 227023
rect 140949 226961 140997 226989
rect 141025 226961 141059 226989
rect 141087 226961 141121 226989
rect 141149 226961 141183 226989
rect 141211 226961 141259 226989
rect 140949 218175 141259 226961
rect 140949 218147 140997 218175
rect 141025 218147 141059 218175
rect 141087 218147 141121 218175
rect 141149 218147 141183 218175
rect 141211 218147 141259 218175
rect 140949 218113 141259 218147
rect 140949 218085 140997 218113
rect 141025 218085 141059 218113
rect 141087 218085 141121 218113
rect 141149 218085 141183 218113
rect 141211 218085 141259 218113
rect 140949 218051 141259 218085
rect 140949 218023 140997 218051
rect 141025 218023 141059 218051
rect 141087 218023 141121 218051
rect 141149 218023 141183 218051
rect 141211 218023 141259 218051
rect 140949 217989 141259 218023
rect 140949 217961 140997 217989
rect 141025 217961 141059 217989
rect 141087 217961 141121 217989
rect 141149 217961 141183 217989
rect 141211 217961 141259 217989
rect 140949 209175 141259 217961
rect 140949 209147 140997 209175
rect 141025 209147 141059 209175
rect 141087 209147 141121 209175
rect 141149 209147 141183 209175
rect 141211 209147 141259 209175
rect 140949 209113 141259 209147
rect 140949 209085 140997 209113
rect 141025 209085 141059 209113
rect 141087 209085 141121 209113
rect 141149 209085 141183 209113
rect 141211 209085 141259 209113
rect 140949 209051 141259 209085
rect 140949 209023 140997 209051
rect 141025 209023 141059 209051
rect 141087 209023 141121 209051
rect 141149 209023 141183 209051
rect 141211 209023 141259 209051
rect 140949 208989 141259 209023
rect 140949 208961 140997 208989
rect 141025 208961 141059 208989
rect 141087 208961 141121 208989
rect 141149 208961 141183 208989
rect 141211 208961 141259 208989
rect 140949 200175 141259 208961
rect 140949 200147 140997 200175
rect 141025 200147 141059 200175
rect 141087 200147 141121 200175
rect 141149 200147 141183 200175
rect 141211 200147 141259 200175
rect 140949 200113 141259 200147
rect 140949 200085 140997 200113
rect 141025 200085 141059 200113
rect 141087 200085 141121 200113
rect 141149 200085 141183 200113
rect 141211 200085 141259 200113
rect 140949 200051 141259 200085
rect 140949 200023 140997 200051
rect 141025 200023 141059 200051
rect 141087 200023 141121 200051
rect 141149 200023 141183 200051
rect 141211 200023 141259 200051
rect 140949 199989 141259 200023
rect 140949 199961 140997 199989
rect 141025 199961 141059 199989
rect 141087 199961 141121 199989
rect 141149 199961 141183 199989
rect 141211 199961 141259 199989
rect 140949 191175 141259 199961
rect 140949 191147 140997 191175
rect 141025 191147 141059 191175
rect 141087 191147 141121 191175
rect 141149 191147 141183 191175
rect 141211 191147 141259 191175
rect 140949 191113 141259 191147
rect 140949 191085 140997 191113
rect 141025 191085 141059 191113
rect 141087 191085 141121 191113
rect 141149 191085 141183 191113
rect 141211 191085 141259 191113
rect 140949 191051 141259 191085
rect 140949 191023 140997 191051
rect 141025 191023 141059 191051
rect 141087 191023 141121 191051
rect 141149 191023 141183 191051
rect 141211 191023 141259 191051
rect 140949 190989 141259 191023
rect 140949 190961 140997 190989
rect 141025 190961 141059 190989
rect 141087 190961 141121 190989
rect 141149 190961 141183 190989
rect 141211 190961 141259 190989
rect 140949 182175 141259 190961
rect 140949 182147 140997 182175
rect 141025 182147 141059 182175
rect 141087 182147 141121 182175
rect 141149 182147 141183 182175
rect 141211 182147 141259 182175
rect 140949 182113 141259 182147
rect 140949 182085 140997 182113
rect 141025 182085 141059 182113
rect 141087 182085 141121 182113
rect 141149 182085 141183 182113
rect 141211 182085 141259 182113
rect 140949 182051 141259 182085
rect 140949 182023 140997 182051
rect 141025 182023 141059 182051
rect 141087 182023 141121 182051
rect 141149 182023 141183 182051
rect 141211 182023 141259 182051
rect 140949 181989 141259 182023
rect 140949 181961 140997 181989
rect 141025 181961 141059 181989
rect 141087 181961 141121 181989
rect 141149 181961 141183 181989
rect 141211 181961 141259 181989
rect 131104 173175 131264 173192
rect 131104 173147 131139 173175
rect 131167 173147 131201 173175
rect 131229 173147 131264 173175
rect 131104 173113 131264 173147
rect 131104 173085 131139 173113
rect 131167 173085 131201 173113
rect 131229 173085 131264 173113
rect 131104 173051 131264 173085
rect 131104 173023 131139 173051
rect 131167 173023 131201 173051
rect 131229 173023 131264 173051
rect 131104 172989 131264 173023
rect 131104 172961 131139 172989
rect 131167 172961 131201 172989
rect 131229 172961 131264 172989
rect 131104 172944 131264 172961
rect 140949 173175 141259 181961
rect 140949 173147 140997 173175
rect 141025 173147 141059 173175
rect 141087 173147 141121 173175
rect 141149 173147 141183 173175
rect 141211 173147 141259 173175
rect 140949 173113 141259 173147
rect 140949 173085 140997 173113
rect 141025 173085 141059 173113
rect 141087 173085 141121 173113
rect 141149 173085 141183 173113
rect 141211 173085 141259 173113
rect 140949 173051 141259 173085
rect 140949 173023 140997 173051
rect 141025 173023 141059 173051
rect 141087 173023 141121 173051
rect 141149 173023 141183 173051
rect 141211 173023 141259 173051
rect 140949 172989 141259 173023
rect 140949 172961 140997 172989
rect 141025 172961 141059 172989
rect 141087 172961 141121 172989
rect 141149 172961 141183 172989
rect 141211 172961 141259 172989
rect 127449 167147 127497 167175
rect 127525 167147 127559 167175
rect 127587 167147 127621 167175
rect 127649 167147 127683 167175
rect 127711 167147 127759 167175
rect 127449 167113 127759 167147
rect 127449 167085 127497 167113
rect 127525 167085 127559 167113
rect 127587 167085 127621 167113
rect 127649 167085 127683 167113
rect 127711 167085 127759 167113
rect 127449 167051 127759 167085
rect 127449 167023 127497 167051
rect 127525 167023 127559 167051
rect 127587 167023 127621 167051
rect 127649 167023 127683 167051
rect 127711 167023 127759 167051
rect 127449 166989 127759 167023
rect 127449 166961 127497 166989
rect 127525 166961 127559 166989
rect 127587 166961 127621 166989
rect 127649 166961 127683 166989
rect 127711 166961 127759 166989
rect 127449 158175 127759 166961
rect 138784 167175 138944 167192
rect 138784 167147 138819 167175
rect 138847 167147 138881 167175
rect 138909 167147 138944 167175
rect 138784 167113 138944 167147
rect 138784 167085 138819 167113
rect 138847 167085 138881 167113
rect 138909 167085 138944 167113
rect 138784 167051 138944 167085
rect 138784 167023 138819 167051
rect 138847 167023 138881 167051
rect 138909 167023 138944 167051
rect 138784 166989 138944 167023
rect 138784 166961 138819 166989
rect 138847 166961 138881 166989
rect 138909 166961 138944 166989
rect 138784 166944 138944 166961
rect 131104 164175 131264 164192
rect 131104 164147 131139 164175
rect 131167 164147 131201 164175
rect 131229 164147 131264 164175
rect 131104 164113 131264 164147
rect 131104 164085 131139 164113
rect 131167 164085 131201 164113
rect 131229 164085 131264 164113
rect 131104 164051 131264 164085
rect 131104 164023 131139 164051
rect 131167 164023 131201 164051
rect 131229 164023 131264 164051
rect 131104 163989 131264 164023
rect 131104 163961 131139 163989
rect 131167 163961 131201 163989
rect 131229 163961 131264 163989
rect 131104 163944 131264 163961
rect 140949 164175 141259 172961
rect 140949 164147 140997 164175
rect 141025 164147 141059 164175
rect 141087 164147 141121 164175
rect 141149 164147 141183 164175
rect 141211 164147 141259 164175
rect 140949 164113 141259 164147
rect 140949 164085 140997 164113
rect 141025 164085 141059 164113
rect 141087 164085 141121 164113
rect 141149 164085 141183 164113
rect 141211 164085 141259 164113
rect 140949 164051 141259 164085
rect 140949 164023 140997 164051
rect 141025 164023 141059 164051
rect 141087 164023 141121 164051
rect 141149 164023 141183 164051
rect 141211 164023 141259 164051
rect 140949 163989 141259 164023
rect 140949 163961 140997 163989
rect 141025 163961 141059 163989
rect 141087 163961 141121 163989
rect 141149 163961 141183 163989
rect 141211 163961 141259 163989
rect 127449 158147 127497 158175
rect 127525 158147 127559 158175
rect 127587 158147 127621 158175
rect 127649 158147 127683 158175
rect 127711 158147 127759 158175
rect 127449 158113 127759 158147
rect 127449 158085 127497 158113
rect 127525 158085 127559 158113
rect 127587 158085 127621 158113
rect 127649 158085 127683 158113
rect 127711 158085 127759 158113
rect 127449 158051 127759 158085
rect 127449 158023 127497 158051
rect 127525 158023 127559 158051
rect 127587 158023 127621 158051
rect 127649 158023 127683 158051
rect 127711 158023 127759 158051
rect 127449 157989 127759 158023
rect 127449 157961 127497 157989
rect 127525 157961 127559 157989
rect 127587 157961 127621 157989
rect 127649 157961 127683 157989
rect 127711 157961 127759 157989
rect 127449 149175 127759 157961
rect 138784 158175 138944 158192
rect 138784 158147 138819 158175
rect 138847 158147 138881 158175
rect 138909 158147 138944 158175
rect 138784 158113 138944 158147
rect 138784 158085 138819 158113
rect 138847 158085 138881 158113
rect 138909 158085 138944 158113
rect 138784 158051 138944 158085
rect 138784 158023 138819 158051
rect 138847 158023 138881 158051
rect 138909 158023 138944 158051
rect 138784 157989 138944 158023
rect 138784 157961 138819 157989
rect 138847 157961 138881 157989
rect 138909 157961 138944 157989
rect 138784 157944 138944 157961
rect 131104 155175 131264 155192
rect 131104 155147 131139 155175
rect 131167 155147 131201 155175
rect 131229 155147 131264 155175
rect 131104 155113 131264 155147
rect 131104 155085 131139 155113
rect 131167 155085 131201 155113
rect 131229 155085 131264 155113
rect 131104 155051 131264 155085
rect 131104 155023 131139 155051
rect 131167 155023 131201 155051
rect 131229 155023 131264 155051
rect 131104 154989 131264 155023
rect 131104 154961 131139 154989
rect 131167 154961 131201 154989
rect 131229 154961 131264 154989
rect 131104 154944 131264 154961
rect 140949 155175 141259 163961
rect 140949 155147 140997 155175
rect 141025 155147 141059 155175
rect 141087 155147 141121 155175
rect 141149 155147 141183 155175
rect 141211 155147 141259 155175
rect 140949 155113 141259 155147
rect 140949 155085 140997 155113
rect 141025 155085 141059 155113
rect 141087 155085 141121 155113
rect 141149 155085 141183 155113
rect 141211 155085 141259 155113
rect 140949 155051 141259 155085
rect 140949 155023 140997 155051
rect 141025 155023 141059 155051
rect 141087 155023 141121 155051
rect 141149 155023 141183 155051
rect 141211 155023 141259 155051
rect 140949 154989 141259 155023
rect 140949 154961 140997 154989
rect 141025 154961 141059 154989
rect 141087 154961 141121 154989
rect 141149 154961 141183 154989
rect 141211 154961 141259 154989
rect 127449 149147 127497 149175
rect 127525 149147 127559 149175
rect 127587 149147 127621 149175
rect 127649 149147 127683 149175
rect 127711 149147 127759 149175
rect 127449 149113 127759 149147
rect 127449 149085 127497 149113
rect 127525 149085 127559 149113
rect 127587 149085 127621 149113
rect 127649 149085 127683 149113
rect 127711 149085 127759 149113
rect 127449 149051 127759 149085
rect 127449 149023 127497 149051
rect 127525 149023 127559 149051
rect 127587 149023 127621 149051
rect 127649 149023 127683 149051
rect 127711 149023 127759 149051
rect 127449 148989 127759 149023
rect 127449 148961 127497 148989
rect 127525 148961 127559 148989
rect 127587 148961 127621 148989
rect 127649 148961 127683 148989
rect 127711 148961 127759 148989
rect 127449 140175 127759 148961
rect 138784 149175 138944 149192
rect 138784 149147 138819 149175
rect 138847 149147 138881 149175
rect 138909 149147 138944 149175
rect 138784 149113 138944 149147
rect 138784 149085 138819 149113
rect 138847 149085 138881 149113
rect 138909 149085 138944 149113
rect 138784 149051 138944 149085
rect 138784 149023 138819 149051
rect 138847 149023 138881 149051
rect 138909 149023 138944 149051
rect 138784 148989 138944 149023
rect 138784 148961 138819 148989
rect 138847 148961 138881 148989
rect 138909 148961 138944 148989
rect 138784 148944 138944 148961
rect 131104 146175 131264 146192
rect 131104 146147 131139 146175
rect 131167 146147 131201 146175
rect 131229 146147 131264 146175
rect 131104 146113 131264 146147
rect 131104 146085 131139 146113
rect 131167 146085 131201 146113
rect 131229 146085 131264 146113
rect 131104 146051 131264 146085
rect 131104 146023 131139 146051
rect 131167 146023 131201 146051
rect 131229 146023 131264 146051
rect 131104 145989 131264 146023
rect 131104 145961 131139 145989
rect 131167 145961 131201 145989
rect 131229 145961 131264 145989
rect 131104 145944 131264 145961
rect 140949 146175 141259 154961
rect 140949 146147 140997 146175
rect 141025 146147 141059 146175
rect 141087 146147 141121 146175
rect 141149 146147 141183 146175
rect 141211 146147 141259 146175
rect 140949 146113 141259 146147
rect 140949 146085 140997 146113
rect 141025 146085 141059 146113
rect 141087 146085 141121 146113
rect 141149 146085 141183 146113
rect 141211 146085 141259 146113
rect 140949 146051 141259 146085
rect 140949 146023 140997 146051
rect 141025 146023 141059 146051
rect 141087 146023 141121 146051
rect 141149 146023 141183 146051
rect 141211 146023 141259 146051
rect 140949 145989 141259 146023
rect 140949 145961 140997 145989
rect 141025 145961 141059 145989
rect 141087 145961 141121 145989
rect 141149 145961 141183 145989
rect 141211 145961 141259 145989
rect 127449 140147 127497 140175
rect 127525 140147 127559 140175
rect 127587 140147 127621 140175
rect 127649 140147 127683 140175
rect 127711 140147 127759 140175
rect 127449 140113 127759 140147
rect 127449 140085 127497 140113
rect 127525 140085 127559 140113
rect 127587 140085 127621 140113
rect 127649 140085 127683 140113
rect 127711 140085 127759 140113
rect 127449 140051 127759 140085
rect 127449 140023 127497 140051
rect 127525 140023 127559 140051
rect 127587 140023 127621 140051
rect 127649 140023 127683 140051
rect 127711 140023 127759 140051
rect 127449 139989 127759 140023
rect 127449 139961 127497 139989
rect 127525 139961 127559 139989
rect 127587 139961 127621 139989
rect 127649 139961 127683 139989
rect 127711 139961 127759 139989
rect 127449 131175 127759 139961
rect 138784 140175 138944 140192
rect 138784 140147 138819 140175
rect 138847 140147 138881 140175
rect 138909 140147 138944 140175
rect 138784 140113 138944 140147
rect 138784 140085 138819 140113
rect 138847 140085 138881 140113
rect 138909 140085 138944 140113
rect 138784 140051 138944 140085
rect 138784 140023 138819 140051
rect 138847 140023 138881 140051
rect 138909 140023 138944 140051
rect 138784 139989 138944 140023
rect 138784 139961 138819 139989
rect 138847 139961 138881 139989
rect 138909 139961 138944 139989
rect 138784 139944 138944 139961
rect 131104 137175 131264 137192
rect 131104 137147 131139 137175
rect 131167 137147 131201 137175
rect 131229 137147 131264 137175
rect 131104 137113 131264 137147
rect 131104 137085 131139 137113
rect 131167 137085 131201 137113
rect 131229 137085 131264 137113
rect 131104 137051 131264 137085
rect 131104 137023 131139 137051
rect 131167 137023 131201 137051
rect 131229 137023 131264 137051
rect 131104 136989 131264 137023
rect 131104 136961 131139 136989
rect 131167 136961 131201 136989
rect 131229 136961 131264 136989
rect 131104 136944 131264 136961
rect 140949 137175 141259 145961
rect 140949 137147 140997 137175
rect 141025 137147 141059 137175
rect 141087 137147 141121 137175
rect 141149 137147 141183 137175
rect 141211 137147 141259 137175
rect 140949 137113 141259 137147
rect 140949 137085 140997 137113
rect 141025 137085 141059 137113
rect 141087 137085 141121 137113
rect 141149 137085 141183 137113
rect 141211 137085 141259 137113
rect 140949 137051 141259 137085
rect 140949 137023 140997 137051
rect 141025 137023 141059 137051
rect 141087 137023 141121 137051
rect 141149 137023 141183 137051
rect 141211 137023 141259 137051
rect 140949 136989 141259 137023
rect 140949 136961 140997 136989
rect 141025 136961 141059 136989
rect 141087 136961 141121 136989
rect 141149 136961 141183 136989
rect 141211 136961 141259 136989
rect 127449 131147 127497 131175
rect 127525 131147 127559 131175
rect 127587 131147 127621 131175
rect 127649 131147 127683 131175
rect 127711 131147 127759 131175
rect 127449 131113 127759 131147
rect 127449 131085 127497 131113
rect 127525 131085 127559 131113
rect 127587 131085 127621 131113
rect 127649 131085 127683 131113
rect 127711 131085 127759 131113
rect 127449 131051 127759 131085
rect 127449 131023 127497 131051
rect 127525 131023 127559 131051
rect 127587 131023 127621 131051
rect 127649 131023 127683 131051
rect 127711 131023 127759 131051
rect 127449 130989 127759 131023
rect 127449 130961 127497 130989
rect 127525 130961 127559 130989
rect 127587 130961 127621 130989
rect 127649 130961 127683 130989
rect 127711 130961 127759 130989
rect 127449 122175 127759 130961
rect 138784 131175 138944 131192
rect 138784 131147 138819 131175
rect 138847 131147 138881 131175
rect 138909 131147 138944 131175
rect 138784 131113 138944 131147
rect 138784 131085 138819 131113
rect 138847 131085 138881 131113
rect 138909 131085 138944 131113
rect 138784 131051 138944 131085
rect 138784 131023 138819 131051
rect 138847 131023 138881 131051
rect 138909 131023 138944 131051
rect 138784 130989 138944 131023
rect 138784 130961 138819 130989
rect 138847 130961 138881 130989
rect 138909 130961 138944 130989
rect 138784 130944 138944 130961
rect 131104 128175 131264 128192
rect 131104 128147 131139 128175
rect 131167 128147 131201 128175
rect 131229 128147 131264 128175
rect 131104 128113 131264 128147
rect 131104 128085 131139 128113
rect 131167 128085 131201 128113
rect 131229 128085 131264 128113
rect 131104 128051 131264 128085
rect 131104 128023 131139 128051
rect 131167 128023 131201 128051
rect 131229 128023 131264 128051
rect 131104 127989 131264 128023
rect 131104 127961 131139 127989
rect 131167 127961 131201 127989
rect 131229 127961 131264 127989
rect 131104 127944 131264 127961
rect 140949 128175 141259 136961
rect 140949 128147 140997 128175
rect 141025 128147 141059 128175
rect 141087 128147 141121 128175
rect 141149 128147 141183 128175
rect 141211 128147 141259 128175
rect 140949 128113 141259 128147
rect 140949 128085 140997 128113
rect 141025 128085 141059 128113
rect 141087 128085 141121 128113
rect 141149 128085 141183 128113
rect 141211 128085 141259 128113
rect 140949 128051 141259 128085
rect 140949 128023 140997 128051
rect 141025 128023 141059 128051
rect 141087 128023 141121 128051
rect 141149 128023 141183 128051
rect 141211 128023 141259 128051
rect 140949 127989 141259 128023
rect 140949 127961 140997 127989
rect 141025 127961 141059 127989
rect 141087 127961 141121 127989
rect 141149 127961 141183 127989
rect 141211 127961 141259 127989
rect 127449 122147 127497 122175
rect 127525 122147 127559 122175
rect 127587 122147 127621 122175
rect 127649 122147 127683 122175
rect 127711 122147 127759 122175
rect 127449 122113 127759 122147
rect 127449 122085 127497 122113
rect 127525 122085 127559 122113
rect 127587 122085 127621 122113
rect 127649 122085 127683 122113
rect 127711 122085 127759 122113
rect 127449 122051 127759 122085
rect 127449 122023 127497 122051
rect 127525 122023 127559 122051
rect 127587 122023 127621 122051
rect 127649 122023 127683 122051
rect 127711 122023 127759 122051
rect 127449 121989 127759 122023
rect 127449 121961 127497 121989
rect 127525 121961 127559 121989
rect 127587 121961 127621 121989
rect 127649 121961 127683 121989
rect 127711 121961 127759 121989
rect 127449 113175 127759 121961
rect 138784 122175 138944 122192
rect 138784 122147 138819 122175
rect 138847 122147 138881 122175
rect 138909 122147 138944 122175
rect 138784 122113 138944 122147
rect 138784 122085 138819 122113
rect 138847 122085 138881 122113
rect 138909 122085 138944 122113
rect 138784 122051 138944 122085
rect 138784 122023 138819 122051
rect 138847 122023 138881 122051
rect 138909 122023 138944 122051
rect 138784 121989 138944 122023
rect 138784 121961 138819 121989
rect 138847 121961 138881 121989
rect 138909 121961 138944 121989
rect 138784 121944 138944 121961
rect 131104 119175 131264 119192
rect 131104 119147 131139 119175
rect 131167 119147 131201 119175
rect 131229 119147 131264 119175
rect 131104 119113 131264 119147
rect 131104 119085 131139 119113
rect 131167 119085 131201 119113
rect 131229 119085 131264 119113
rect 131104 119051 131264 119085
rect 131104 119023 131139 119051
rect 131167 119023 131201 119051
rect 131229 119023 131264 119051
rect 131104 118989 131264 119023
rect 131104 118961 131139 118989
rect 131167 118961 131201 118989
rect 131229 118961 131264 118989
rect 131104 118944 131264 118961
rect 140949 119175 141259 127961
rect 140949 119147 140997 119175
rect 141025 119147 141059 119175
rect 141087 119147 141121 119175
rect 141149 119147 141183 119175
rect 141211 119147 141259 119175
rect 140949 119113 141259 119147
rect 140949 119085 140997 119113
rect 141025 119085 141059 119113
rect 141087 119085 141121 119113
rect 141149 119085 141183 119113
rect 141211 119085 141259 119113
rect 140949 119051 141259 119085
rect 140949 119023 140997 119051
rect 141025 119023 141059 119051
rect 141087 119023 141121 119051
rect 141149 119023 141183 119051
rect 141211 119023 141259 119051
rect 140949 118989 141259 119023
rect 140949 118961 140997 118989
rect 141025 118961 141059 118989
rect 141087 118961 141121 118989
rect 141149 118961 141183 118989
rect 141211 118961 141259 118989
rect 127449 113147 127497 113175
rect 127525 113147 127559 113175
rect 127587 113147 127621 113175
rect 127649 113147 127683 113175
rect 127711 113147 127759 113175
rect 127449 113113 127759 113147
rect 127449 113085 127497 113113
rect 127525 113085 127559 113113
rect 127587 113085 127621 113113
rect 127649 113085 127683 113113
rect 127711 113085 127759 113113
rect 127449 113051 127759 113085
rect 127449 113023 127497 113051
rect 127525 113023 127559 113051
rect 127587 113023 127621 113051
rect 127649 113023 127683 113051
rect 127711 113023 127759 113051
rect 127449 112989 127759 113023
rect 127449 112961 127497 112989
rect 127525 112961 127559 112989
rect 127587 112961 127621 112989
rect 127649 112961 127683 112989
rect 127711 112961 127759 112989
rect 127449 104175 127759 112961
rect 138784 113175 138944 113192
rect 138784 113147 138819 113175
rect 138847 113147 138881 113175
rect 138909 113147 138944 113175
rect 138784 113113 138944 113147
rect 138784 113085 138819 113113
rect 138847 113085 138881 113113
rect 138909 113085 138944 113113
rect 138784 113051 138944 113085
rect 138784 113023 138819 113051
rect 138847 113023 138881 113051
rect 138909 113023 138944 113051
rect 138784 112989 138944 113023
rect 138784 112961 138819 112989
rect 138847 112961 138881 112989
rect 138909 112961 138944 112989
rect 138784 112944 138944 112961
rect 131104 110175 131264 110192
rect 131104 110147 131139 110175
rect 131167 110147 131201 110175
rect 131229 110147 131264 110175
rect 131104 110113 131264 110147
rect 131104 110085 131139 110113
rect 131167 110085 131201 110113
rect 131229 110085 131264 110113
rect 131104 110051 131264 110085
rect 131104 110023 131139 110051
rect 131167 110023 131201 110051
rect 131229 110023 131264 110051
rect 131104 109989 131264 110023
rect 131104 109961 131139 109989
rect 131167 109961 131201 109989
rect 131229 109961 131264 109989
rect 131104 109944 131264 109961
rect 140949 110175 141259 118961
rect 140949 110147 140997 110175
rect 141025 110147 141059 110175
rect 141087 110147 141121 110175
rect 141149 110147 141183 110175
rect 141211 110147 141259 110175
rect 140949 110113 141259 110147
rect 140949 110085 140997 110113
rect 141025 110085 141059 110113
rect 141087 110085 141121 110113
rect 141149 110085 141183 110113
rect 141211 110085 141259 110113
rect 140949 110051 141259 110085
rect 140949 110023 140997 110051
rect 141025 110023 141059 110051
rect 141087 110023 141121 110051
rect 141149 110023 141183 110051
rect 141211 110023 141259 110051
rect 140949 109989 141259 110023
rect 140949 109961 140997 109989
rect 141025 109961 141059 109989
rect 141087 109961 141121 109989
rect 141149 109961 141183 109989
rect 141211 109961 141259 109989
rect 127449 104147 127497 104175
rect 127525 104147 127559 104175
rect 127587 104147 127621 104175
rect 127649 104147 127683 104175
rect 127711 104147 127759 104175
rect 127449 104113 127759 104147
rect 127449 104085 127497 104113
rect 127525 104085 127559 104113
rect 127587 104085 127621 104113
rect 127649 104085 127683 104113
rect 127711 104085 127759 104113
rect 127449 104051 127759 104085
rect 127449 104023 127497 104051
rect 127525 104023 127559 104051
rect 127587 104023 127621 104051
rect 127649 104023 127683 104051
rect 127711 104023 127759 104051
rect 127449 103989 127759 104023
rect 127449 103961 127497 103989
rect 127525 103961 127559 103989
rect 127587 103961 127621 103989
rect 127649 103961 127683 103989
rect 127711 103961 127759 103989
rect 127449 95175 127759 103961
rect 138784 104175 138944 104192
rect 138784 104147 138819 104175
rect 138847 104147 138881 104175
rect 138909 104147 138944 104175
rect 138784 104113 138944 104147
rect 138784 104085 138819 104113
rect 138847 104085 138881 104113
rect 138909 104085 138944 104113
rect 138784 104051 138944 104085
rect 138784 104023 138819 104051
rect 138847 104023 138881 104051
rect 138909 104023 138944 104051
rect 138784 103989 138944 104023
rect 138784 103961 138819 103989
rect 138847 103961 138881 103989
rect 138909 103961 138944 103989
rect 138784 103944 138944 103961
rect 131104 101175 131264 101192
rect 131104 101147 131139 101175
rect 131167 101147 131201 101175
rect 131229 101147 131264 101175
rect 131104 101113 131264 101147
rect 131104 101085 131139 101113
rect 131167 101085 131201 101113
rect 131229 101085 131264 101113
rect 131104 101051 131264 101085
rect 131104 101023 131139 101051
rect 131167 101023 131201 101051
rect 131229 101023 131264 101051
rect 131104 100989 131264 101023
rect 131104 100961 131139 100989
rect 131167 100961 131201 100989
rect 131229 100961 131264 100989
rect 131104 100944 131264 100961
rect 140949 101175 141259 109961
rect 140949 101147 140997 101175
rect 141025 101147 141059 101175
rect 141087 101147 141121 101175
rect 141149 101147 141183 101175
rect 141211 101147 141259 101175
rect 140949 101113 141259 101147
rect 140949 101085 140997 101113
rect 141025 101085 141059 101113
rect 141087 101085 141121 101113
rect 141149 101085 141183 101113
rect 141211 101085 141259 101113
rect 140949 101051 141259 101085
rect 140949 101023 140997 101051
rect 141025 101023 141059 101051
rect 141087 101023 141121 101051
rect 141149 101023 141183 101051
rect 141211 101023 141259 101051
rect 140949 100989 141259 101023
rect 140949 100961 140997 100989
rect 141025 100961 141059 100989
rect 141087 100961 141121 100989
rect 141149 100961 141183 100989
rect 141211 100961 141259 100989
rect 127449 95147 127497 95175
rect 127525 95147 127559 95175
rect 127587 95147 127621 95175
rect 127649 95147 127683 95175
rect 127711 95147 127759 95175
rect 127449 95113 127759 95147
rect 127449 95085 127497 95113
rect 127525 95085 127559 95113
rect 127587 95085 127621 95113
rect 127649 95085 127683 95113
rect 127711 95085 127759 95113
rect 127449 95051 127759 95085
rect 127449 95023 127497 95051
rect 127525 95023 127559 95051
rect 127587 95023 127621 95051
rect 127649 95023 127683 95051
rect 127711 95023 127759 95051
rect 127449 94989 127759 95023
rect 127449 94961 127497 94989
rect 127525 94961 127559 94989
rect 127587 94961 127621 94989
rect 127649 94961 127683 94989
rect 127711 94961 127759 94989
rect 127449 86175 127759 94961
rect 138784 95175 138944 95192
rect 138784 95147 138819 95175
rect 138847 95147 138881 95175
rect 138909 95147 138944 95175
rect 138784 95113 138944 95147
rect 138784 95085 138819 95113
rect 138847 95085 138881 95113
rect 138909 95085 138944 95113
rect 138784 95051 138944 95085
rect 138784 95023 138819 95051
rect 138847 95023 138881 95051
rect 138909 95023 138944 95051
rect 138784 94989 138944 95023
rect 138784 94961 138819 94989
rect 138847 94961 138881 94989
rect 138909 94961 138944 94989
rect 138784 94944 138944 94961
rect 131104 92175 131264 92192
rect 131104 92147 131139 92175
rect 131167 92147 131201 92175
rect 131229 92147 131264 92175
rect 131104 92113 131264 92147
rect 131104 92085 131139 92113
rect 131167 92085 131201 92113
rect 131229 92085 131264 92113
rect 131104 92051 131264 92085
rect 131104 92023 131139 92051
rect 131167 92023 131201 92051
rect 131229 92023 131264 92051
rect 131104 91989 131264 92023
rect 131104 91961 131139 91989
rect 131167 91961 131201 91989
rect 131229 91961 131264 91989
rect 131104 91944 131264 91961
rect 140949 92175 141259 100961
rect 140949 92147 140997 92175
rect 141025 92147 141059 92175
rect 141087 92147 141121 92175
rect 141149 92147 141183 92175
rect 141211 92147 141259 92175
rect 140949 92113 141259 92147
rect 140949 92085 140997 92113
rect 141025 92085 141059 92113
rect 141087 92085 141121 92113
rect 141149 92085 141183 92113
rect 141211 92085 141259 92113
rect 140949 92051 141259 92085
rect 140949 92023 140997 92051
rect 141025 92023 141059 92051
rect 141087 92023 141121 92051
rect 141149 92023 141183 92051
rect 141211 92023 141259 92051
rect 140949 91989 141259 92023
rect 140949 91961 140997 91989
rect 141025 91961 141059 91989
rect 141087 91961 141121 91989
rect 141149 91961 141183 91989
rect 141211 91961 141259 91989
rect 127449 86147 127497 86175
rect 127525 86147 127559 86175
rect 127587 86147 127621 86175
rect 127649 86147 127683 86175
rect 127711 86147 127759 86175
rect 127449 86113 127759 86147
rect 127449 86085 127497 86113
rect 127525 86085 127559 86113
rect 127587 86085 127621 86113
rect 127649 86085 127683 86113
rect 127711 86085 127759 86113
rect 127449 86051 127759 86085
rect 127449 86023 127497 86051
rect 127525 86023 127559 86051
rect 127587 86023 127621 86051
rect 127649 86023 127683 86051
rect 127711 86023 127759 86051
rect 127449 85989 127759 86023
rect 127449 85961 127497 85989
rect 127525 85961 127559 85989
rect 127587 85961 127621 85989
rect 127649 85961 127683 85989
rect 127711 85961 127759 85989
rect 127449 77175 127759 85961
rect 138784 86175 138944 86192
rect 138784 86147 138819 86175
rect 138847 86147 138881 86175
rect 138909 86147 138944 86175
rect 138784 86113 138944 86147
rect 138784 86085 138819 86113
rect 138847 86085 138881 86113
rect 138909 86085 138944 86113
rect 138784 86051 138944 86085
rect 138784 86023 138819 86051
rect 138847 86023 138881 86051
rect 138909 86023 138944 86051
rect 138784 85989 138944 86023
rect 138784 85961 138819 85989
rect 138847 85961 138881 85989
rect 138909 85961 138944 85989
rect 138784 85944 138944 85961
rect 131104 83175 131264 83192
rect 131104 83147 131139 83175
rect 131167 83147 131201 83175
rect 131229 83147 131264 83175
rect 131104 83113 131264 83147
rect 131104 83085 131139 83113
rect 131167 83085 131201 83113
rect 131229 83085 131264 83113
rect 131104 83051 131264 83085
rect 131104 83023 131139 83051
rect 131167 83023 131201 83051
rect 131229 83023 131264 83051
rect 131104 82989 131264 83023
rect 131104 82961 131139 82989
rect 131167 82961 131201 82989
rect 131229 82961 131264 82989
rect 131104 82944 131264 82961
rect 140949 83175 141259 91961
rect 140949 83147 140997 83175
rect 141025 83147 141059 83175
rect 141087 83147 141121 83175
rect 141149 83147 141183 83175
rect 141211 83147 141259 83175
rect 140949 83113 141259 83147
rect 140949 83085 140997 83113
rect 141025 83085 141059 83113
rect 141087 83085 141121 83113
rect 141149 83085 141183 83113
rect 141211 83085 141259 83113
rect 140949 83051 141259 83085
rect 140949 83023 140997 83051
rect 141025 83023 141059 83051
rect 141087 83023 141121 83051
rect 141149 83023 141183 83051
rect 141211 83023 141259 83051
rect 140949 82989 141259 83023
rect 140949 82961 140997 82989
rect 141025 82961 141059 82989
rect 141087 82961 141121 82989
rect 141149 82961 141183 82989
rect 141211 82961 141259 82989
rect 127449 77147 127497 77175
rect 127525 77147 127559 77175
rect 127587 77147 127621 77175
rect 127649 77147 127683 77175
rect 127711 77147 127759 77175
rect 127449 77113 127759 77147
rect 127449 77085 127497 77113
rect 127525 77085 127559 77113
rect 127587 77085 127621 77113
rect 127649 77085 127683 77113
rect 127711 77085 127759 77113
rect 127449 77051 127759 77085
rect 127449 77023 127497 77051
rect 127525 77023 127559 77051
rect 127587 77023 127621 77051
rect 127649 77023 127683 77051
rect 127711 77023 127759 77051
rect 127449 76989 127759 77023
rect 127449 76961 127497 76989
rect 127525 76961 127559 76989
rect 127587 76961 127621 76989
rect 127649 76961 127683 76989
rect 127711 76961 127759 76989
rect 127449 68175 127759 76961
rect 138784 77175 138944 77192
rect 138784 77147 138819 77175
rect 138847 77147 138881 77175
rect 138909 77147 138944 77175
rect 138784 77113 138944 77147
rect 138784 77085 138819 77113
rect 138847 77085 138881 77113
rect 138909 77085 138944 77113
rect 138784 77051 138944 77085
rect 138784 77023 138819 77051
rect 138847 77023 138881 77051
rect 138909 77023 138944 77051
rect 138784 76989 138944 77023
rect 138784 76961 138819 76989
rect 138847 76961 138881 76989
rect 138909 76961 138944 76989
rect 138784 76944 138944 76961
rect 131104 74175 131264 74192
rect 131104 74147 131139 74175
rect 131167 74147 131201 74175
rect 131229 74147 131264 74175
rect 131104 74113 131264 74147
rect 131104 74085 131139 74113
rect 131167 74085 131201 74113
rect 131229 74085 131264 74113
rect 131104 74051 131264 74085
rect 131104 74023 131139 74051
rect 131167 74023 131201 74051
rect 131229 74023 131264 74051
rect 131104 73989 131264 74023
rect 131104 73961 131139 73989
rect 131167 73961 131201 73989
rect 131229 73961 131264 73989
rect 131104 73944 131264 73961
rect 140949 74175 141259 82961
rect 140949 74147 140997 74175
rect 141025 74147 141059 74175
rect 141087 74147 141121 74175
rect 141149 74147 141183 74175
rect 141211 74147 141259 74175
rect 140949 74113 141259 74147
rect 140949 74085 140997 74113
rect 141025 74085 141059 74113
rect 141087 74085 141121 74113
rect 141149 74085 141183 74113
rect 141211 74085 141259 74113
rect 140949 74051 141259 74085
rect 140949 74023 140997 74051
rect 141025 74023 141059 74051
rect 141087 74023 141121 74051
rect 141149 74023 141183 74051
rect 141211 74023 141259 74051
rect 140949 73989 141259 74023
rect 140949 73961 140997 73989
rect 141025 73961 141059 73989
rect 141087 73961 141121 73989
rect 141149 73961 141183 73989
rect 141211 73961 141259 73989
rect 127449 68147 127497 68175
rect 127525 68147 127559 68175
rect 127587 68147 127621 68175
rect 127649 68147 127683 68175
rect 127711 68147 127759 68175
rect 127449 68113 127759 68147
rect 127449 68085 127497 68113
rect 127525 68085 127559 68113
rect 127587 68085 127621 68113
rect 127649 68085 127683 68113
rect 127711 68085 127759 68113
rect 127449 68051 127759 68085
rect 127449 68023 127497 68051
rect 127525 68023 127559 68051
rect 127587 68023 127621 68051
rect 127649 68023 127683 68051
rect 127711 68023 127759 68051
rect 127449 67989 127759 68023
rect 127449 67961 127497 67989
rect 127525 67961 127559 67989
rect 127587 67961 127621 67989
rect 127649 67961 127683 67989
rect 127711 67961 127759 67989
rect 127449 59175 127759 67961
rect 138784 68175 138944 68192
rect 138784 68147 138819 68175
rect 138847 68147 138881 68175
rect 138909 68147 138944 68175
rect 138784 68113 138944 68147
rect 138784 68085 138819 68113
rect 138847 68085 138881 68113
rect 138909 68085 138944 68113
rect 138784 68051 138944 68085
rect 138784 68023 138819 68051
rect 138847 68023 138881 68051
rect 138909 68023 138944 68051
rect 138784 67989 138944 68023
rect 138784 67961 138819 67989
rect 138847 67961 138881 67989
rect 138909 67961 138944 67989
rect 138784 67944 138944 67961
rect 131104 65175 131264 65192
rect 131104 65147 131139 65175
rect 131167 65147 131201 65175
rect 131229 65147 131264 65175
rect 131104 65113 131264 65147
rect 131104 65085 131139 65113
rect 131167 65085 131201 65113
rect 131229 65085 131264 65113
rect 131104 65051 131264 65085
rect 131104 65023 131139 65051
rect 131167 65023 131201 65051
rect 131229 65023 131264 65051
rect 131104 64989 131264 65023
rect 131104 64961 131139 64989
rect 131167 64961 131201 64989
rect 131229 64961 131264 64989
rect 131104 64944 131264 64961
rect 140949 65175 141259 73961
rect 140949 65147 140997 65175
rect 141025 65147 141059 65175
rect 141087 65147 141121 65175
rect 141149 65147 141183 65175
rect 141211 65147 141259 65175
rect 140949 65113 141259 65147
rect 140949 65085 140997 65113
rect 141025 65085 141059 65113
rect 141087 65085 141121 65113
rect 141149 65085 141183 65113
rect 141211 65085 141259 65113
rect 140949 65051 141259 65085
rect 140949 65023 140997 65051
rect 141025 65023 141059 65051
rect 141087 65023 141121 65051
rect 141149 65023 141183 65051
rect 141211 65023 141259 65051
rect 140949 64989 141259 65023
rect 140949 64961 140997 64989
rect 141025 64961 141059 64989
rect 141087 64961 141121 64989
rect 141149 64961 141183 64989
rect 141211 64961 141259 64989
rect 127449 59147 127497 59175
rect 127525 59147 127559 59175
rect 127587 59147 127621 59175
rect 127649 59147 127683 59175
rect 127711 59147 127759 59175
rect 127449 59113 127759 59147
rect 127449 59085 127497 59113
rect 127525 59085 127559 59113
rect 127587 59085 127621 59113
rect 127649 59085 127683 59113
rect 127711 59085 127759 59113
rect 127449 59051 127759 59085
rect 127449 59023 127497 59051
rect 127525 59023 127559 59051
rect 127587 59023 127621 59051
rect 127649 59023 127683 59051
rect 127711 59023 127759 59051
rect 127449 58989 127759 59023
rect 127449 58961 127497 58989
rect 127525 58961 127559 58989
rect 127587 58961 127621 58989
rect 127649 58961 127683 58989
rect 127711 58961 127759 58989
rect 127449 50175 127759 58961
rect 138784 59175 138944 59192
rect 138784 59147 138819 59175
rect 138847 59147 138881 59175
rect 138909 59147 138944 59175
rect 138784 59113 138944 59147
rect 138784 59085 138819 59113
rect 138847 59085 138881 59113
rect 138909 59085 138944 59113
rect 138784 59051 138944 59085
rect 138784 59023 138819 59051
rect 138847 59023 138881 59051
rect 138909 59023 138944 59051
rect 138784 58989 138944 59023
rect 138784 58961 138819 58989
rect 138847 58961 138881 58989
rect 138909 58961 138944 58989
rect 138784 58944 138944 58961
rect 131104 56175 131264 56192
rect 131104 56147 131139 56175
rect 131167 56147 131201 56175
rect 131229 56147 131264 56175
rect 131104 56113 131264 56147
rect 131104 56085 131139 56113
rect 131167 56085 131201 56113
rect 131229 56085 131264 56113
rect 131104 56051 131264 56085
rect 131104 56023 131139 56051
rect 131167 56023 131201 56051
rect 131229 56023 131264 56051
rect 131104 55989 131264 56023
rect 131104 55961 131139 55989
rect 131167 55961 131201 55989
rect 131229 55961 131264 55989
rect 131104 55944 131264 55961
rect 140949 56175 141259 64961
rect 140949 56147 140997 56175
rect 141025 56147 141059 56175
rect 141087 56147 141121 56175
rect 141149 56147 141183 56175
rect 141211 56147 141259 56175
rect 140949 56113 141259 56147
rect 140949 56085 140997 56113
rect 141025 56085 141059 56113
rect 141087 56085 141121 56113
rect 141149 56085 141183 56113
rect 141211 56085 141259 56113
rect 140949 56051 141259 56085
rect 140949 56023 140997 56051
rect 141025 56023 141059 56051
rect 141087 56023 141121 56051
rect 141149 56023 141183 56051
rect 141211 56023 141259 56051
rect 140949 55989 141259 56023
rect 140949 55961 140997 55989
rect 141025 55961 141059 55989
rect 141087 55961 141121 55989
rect 141149 55961 141183 55989
rect 141211 55961 141259 55989
rect 127449 50147 127497 50175
rect 127525 50147 127559 50175
rect 127587 50147 127621 50175
rect 127649 50147 127683 50175
rect 127711 50147 127759 50175
rect 127449 50113 127759 50147
rect 127449 50085 127497 50113
rect 127525 50085 127559 50113
rect 127587 50085 127621 50113
rect 127649 50085 127683 50113
rect 127711 50085 127759 50113
rect 127449 50051 127759 50085
rect 127449 50023 127497 50051
rect 127525 50023 127559 50051
rect 127587 50023 127621 50051
rect 127649 50023 127683 50051
rect 127711 50023 127759 50051
rect 127449 49989 127759 50023
rect 127449 49961 127497 49989
rect 127525 49961 127559 49989
rect 127587 49961 127621 49989
rect 127649 49961 127683 49989
rect 127711 49961 127759 49989
rect 127449 41175 127759 49961
rect 138784 50175 138944 50192
rect 138784 50147 138819 50175
rect 138847 50147 138881 50175
rect 138909 50147 138944 50175
rect 138784 50113 138944 50147
rect 138784 50085 138819 50113
rect 138847 50085 138881 50113
rect 138909 50085 138944 50113
rect 138784 50051 138944 50085
rect 138784 50023 138819 50051
rect 138847 50023 138881 50051
rect 138909 50023 138944 50051
rect 138784 49989 138944 50023
rect 138784 49961 138819 49989
rect 138847 49961 138881 49989
rect 138909 49961 138944 49989
rect 138784 49944 138944 49961
rect 131104 47175 131264 47192
rect 131104 47147 131139 47175
rect 131167 47147 131201 47175
rect 131229 47147 131264 47175
rect 131104 47113 131264 47147
rect 131104 47085 131139 47113
rect 131167 47085 131201 47113
rect 131229 47085 131264 47113
rect 131104 47051 131264 47085
rect 131104 47023 131139 47051
rect 131167 47023 131201 47051
rect 131229 47023 131264 47051
rect 131104 46989 131264 47023
rect 131104 46961 131139 46989
rect 131167 46961 131201 46989
rect 131229 46961 131264 46989
rect 131104 46944 131264 46961
rect 140949 47175 141259 55961
rect 140949 47147 140997 47175
rect 141025 47147 141059 47175
rect 141087 47147 141121 47175
rect 141149 47147 141183 47175
rect 141211 47147 141259 47175
rect 140949 47113 141259 47147
rect 140949 47085 140997 47113
rect 141025 47085 141059 47113
rect 141087 47085 141121 47113
rect 141149 47085 141183 47113
rect 141211 47085 141259 47113
rect 140949 47051 141259 47085
rect 140949 47023 140997 47051
rect 141025 47023 141059 47051
rect 141087 47023 141121 47051
rect 141149 47023 141183 47051
rect 141211 47023 141259 47051
rect 140949 46989 141259 47023
rect 140949 46961 140997 46989
rect 141025 46961 141059 46989
rect 141087 46961 141121 46989
rect 141149 46961 141183 46989
rect 141211 46961 141259 46989
rect 127449 41147 127497 41175
rect 127525 41147 127559 41175
rect 127587 41147 127621 41175
rect 127649 41147 127683 41175
rect 127711 41147 127759 41175
rect 127449 41113 127759 41147
rect 127449 41085 127497 41113
rect 127525 41085 127559 41113
rect 127587 41085 127621 41113
rect 127649 41085 127683 41113
rect 127711 41085 127759 41113
rect 127449 41051 127759 41085
rect 127449 41023 127497 41051
rect 127525 41023 127559 41051
rect 127587 41023 127621 41051
rect 127649 41023 127683 41051
rect 127711 41023 127759 41051
rect 127449 40989 127759 41023
rect 127449 40961 127497 40989
rect 127525 40961 127559 40989
rect 127587 40961 127621 40989
rect 127649 40961 127683 40989
rect 127711 40961 127759 40989
rect 127449 32175 127759 40961
rect 138784 41175 138944 41192
rect 138784 41147 138819 41175
rect 138847 41147 138881 41175
rect 138909 41147 138944 41175
rect 138784 41113 138944 41147
rect 138784 41085 138819 41113
rect 138847 41085 138881 41113
rect 138909 41085 138944 41113
rect 138784 41051 138944 41085
rect 138784 41023 138819 41051
rect 138847 41023 138881 41051
rect 138909 41023 138944 41051
rect 138784 40989 138944 41023
rect 138784 40961 138819 40989
rect 138847 40961 138881 40989
rect 138909 40961 138944 40989
rect 138784 40944 138944 40961
rect 131104 38175 131264 38192
rect 131104 38147 131139 38175
rect 131167 38147 131201 38175
rect 131229 38147 131264 38175
rect 131104 38113 131264 38147
rect 131104 38085 131139 38113
rect 131167 38085 131201 38113
rect 131229 38085 131264 38113
rect 131104 38051 131264 38085
rect 131104 38023 131139 38051
rect 131167 38023 131201 38051
rect 131229 38023 131264 38051
rect 131104 37989 131264 38023
rect 131104 37961 131139 37989
rect 131167 37961 131201 37989
rect 131229 37961 131264 37989
rect 131104 37944 131264 37961
rect 140949 38175 141259 46961
rect 140949 38147 140997 38175
rect 141025 38147 141059 38175
rect 141087 38147 141121 38175
rect 141149 38147 141183 38175
rect 141211 38147 141259 38175
rect 140949 38113 141259 38147
rect 140949 38085 140997 38113
rect 141025 38085 141059 38113
rect 141087 38085 141121 38113
rect 141149 38085 141183 38113
rect 141211 38085 141259 38113
rect 140949 38051 141259 38085
rect 140949 38023 140997 38051
rect 141025 38023 141059 38051
rect 141087 38023 141121 38051
rect 141149 38023 141183 38051
rect 141211 38023 141259 38051
rect 140949 37989 141259 38023
rect 140949 37961 140997 37989
rect 141025 37961 141059 37989
rect 141087 37961 141121 37989
rect 141149 37961 141183 37989
rect 141211 37961 141259 37989
rect 127449 32147 127497 32175
rect 127525 32147 127559 32175
rect 127587 32147 127621 32175
rect 127649 32147 127683 32175
rect 127711 32147 127759 32175
rect 127449 32113 127759 32147
rect 127449 32085 127497 32113
rect 127525 32085 127559 32113
rect 127587 32085 127621 32113
rect 127649 32085 127683 32113
rect 127711 32085 127759 32113
rect 127449 32051 127759 32085
rect 127449 32023 127497 32051
rect 127525 32023 127559 32051
rect 127587 32023 127621 32051
rect 127649 32023 127683 32051
rect 127711 32023 127759 32051
rect 127449 31989 127759 32023
rect 127449 31961 127497 31989
rect 127525 31961 127559 31989
rect 127587 31961 127621 31989
rect 127649 31961 127683 31989
rect 127711 31961 127759 31989
rect 127449 23175 127759 31961
rect 138784 32175 138944 32192
rect 138784 32147 138819 32175
rect 138847 32147 138881 32175
rect 138909 32147 138944 32175
rect 138784 32113 138944 32147
rect 138784 32085 138819 32113
rect 138847 32085 138881 32113
rect 138909 32085 138944 32113
rect 138784 32051 138944 32085
rect 138784 32023 138819 32051
rect 138847 32023 138881 32051
rect 138909 32023 138944 32051
rect 138784 31989 138944 32023
rect 138784 31961 138819 31989
rect 138847 31961 138881 31989
rect 138909 31961 138944 31989
rect 138784 31944 138944 31961
rect 131104 29175 131264 29192
rect 131104 29147 131139 29175
rect 131167 29147 131201 29175
rect 131229 29147 131264 29175
rect 131104 29113 131264 29147
rect 131104 29085 131139 29113
rect 131167 29085 131201 29113
rect 131229 29085 131264 29113
rect 131104 29051 131264 29085
rect 131104 29023 131139 29051
rect 131167 29023 131201 29051
rect 131229 29023 131264 29051
rect 131104 28989 131264 29023
rect 131104 28961 131139 28989
rect 131167 28961 131201 28989
rect 131229 28961 131264 28989
rect 131104 28944 131264 28961
rect 140949 29175 141259 37961
rect 140949 29147 140997 29175
rect 141025 29147 141059 29175
rect 141087 29147 141121 29175
rect 141149 29147 141183 29175
rect 141211 29147 141259 29175
rect 140949 29113 141259 29147
rect 140949 29085 140997 29113
rect 141025 29085 141059 29113
rect 141087 29085 141121 29113
rect 141149 29085 141183 29113
rect 141211 29085 141259 29113
rect 140949 29051 141259 29085
rect 140949 29023 140997 29051
rect 141025 29023 141059 29051
rect 141087 29023 141121 29051
rect 141149 29023 141183 29051
rect 141211 29023 141259 29051
rect 140949 28989 141259 29023
rect 140949 28961 140997 28989
rect 141025 28961 141059 28989
rect 141087 28961 141121 28989
rect 141149 28961 141183 28989
rect 141211 28961 141259 28989
rect 127449 23147 127497 23175
rect 127525 23147 127559 23175
rect 127587 23147 127621 23175
rect 127649 23147 127683 23175
rect 127711 23147 127759 23175
rect 127449 23113 127759 23147
rect 127449 23085 127497 23113
rect 127525 23085 127559 23113
rect 127587 23085 127621 23113
rect 127649 23085 127683 23113
rect 127711 23085 127759 23113
rect 127449 23051 127759 23085
rect 127449 23023 127497 23051
rect 127525 23023 127559 23051
rect 127587 23023 127621 23051
rect 127649 23023 127683 23051
rect 127711 23023 127759 23051
rect 127449 22989 127759 23023
rect 127449 22961 127497 22989
rect 127525 22961 127559 22989
rect 127587 22961 127621 22989
rect 127649 22961 127683 22989
rect 127711 22961 127759 22989
rect 127449 14175 127759 22961
rect 138784 23175 138944 23192
rect 138784 23147 138819 23175
rect 138847 23147 138881 23175
rect 138909 23147 138944 23175
rect 138784 23113 138944 23147
rect 138784 23085 138819 23113
rect 138847 23085 138881 23113
rect 138909 23085 138944 23113
rect 138784 23051 138944 23085
rect 138784 23023 138819 23051
rect 138847 23023 138881 23051
rect 138909 23023 138944 23051
rect 138784 22989 138944 23023
rect 138784 22961 138819 22989
rect 138847 22961 138881 22989
rect 138909 22961 138944 22989
rect 138784 22944 138944 22961
rect 131104 20175 131264 20192
rect 131104 20147 131139 20175
rect 131167 20147 131201 20175
rect 131229 20147 131264 20175
rect 131104 20113 131264 20147
rect 131104 20085 131139 20113
rect 131167 20085 131201 20113
rect 131229 20085 131264 20113
rect 131104 20051 131264 20085
rect 131104 20023 131139 20051
rect 131167 20023 131201 20051
rect 131229 20023 131264 20051
rect 131104 19989 131264 20023
rect 131104 19961 131139 19989
rect 131167 19961 131201 19989
rect 131229 19961 131264 19989
rect 131104 19944 131264 19961
rect 140949 20175 141259 28961
rect 140949 20147 140997 20175
rect 141025 20147 141059 20175
rect 141087 20147 141121 20175
rect 141149 20147 141183 20175
rect 141211 20147 141259 20175
rect 140949 20113 141259 20147
rect 140949 20085 140997 20113
rect 141025 20085 141059 20113
rect 141087 20085 141121 20113
rect 141149 20085 141183 20113
rect 141211 20085 141259 20113
rect 140949 20051 141259 20085
rect 140949 20023 140997 20051
rect 141025 20023 141059 20051
rect 141087 20023 141121 20051
rect 141149 20023 141183 20051
rect 141211 20023 141259 20051
rect 140949 19989 141259 20023
rect 140949 19961 140997 19989
rect 141025 19961 141059 19989
rect 141087 19961 141121 19989
rect 141149 19961 141183 19989
rect 141211 19961 141259 19989
rect 127449 14147 127497 14175
rect 127525 14147 127559 14175
rect 127587 14147 127621 14175
rect 127649 14147 127683 14175
rect 127711 14147 127759 14175
rect 127449 14113 127759 14147
rect 127449 14085 127497 14113
rect 127525 14085 127559 14113
rect 127587 14085 127621 14113
rect 127649 14085 127683 14113
rect 127711 14085 127759 14113
rect 127449 14051 127759 14085
rect 127449 14023 127497 14051
rect 127525 14023 127559 14051
rect 127587 14023 127621 14051
rect 127649 14023 127683 14051
rect 127711 14023 127759 14051
rect 127449 13989 127759 14023
rect 127449 13961 127497 13989
rect 127525 13961 127559 13989
rect 127587 13961 127621 13989
rect 127649 13961 127683 13989
rect 127711 13961 127759 13989
rect 127449 5175 127759 13961
rect 138784 14175 138944 14192
rect 138784 14147 138819 14175
rect 138847 14147 138881 14175
rect 138909 14147 138944 14175
rect 138784 14113 138944 14147
rect 138784 14085 138819 14113
rect 138847 14085 138881 14113
rect 138909 14085 138944 14113
rect 138784 14051 138944 14085
rect 138784 14023 138819 14051
rect 138847 14023 138881 14051
rect 138909 14023 138944 14051
rect 138784 13989 138944 14023
rect 138784 13961 138819 13989
rect 138847 13961 138881 13989
rect 138909 13961 138944 13989
rect 138784 13944 138944 13961
rect 131104 11175 131264 11192
rect 131104 11147 131139 11175
rect 131167 11147 131201 11175
rect 131229 11147 131264 11175
rect 131104 11113 131264 11147
rect 131104 11085 131139 11113
rect 131167 11085 131201 11113
rect 131229 11085 131264 11113
rect 131104 11051 131264 11085
rect 131104 11023 131139 11051
rect 131167 11023 131201 11051
rect 131229 11023 131264 11051
rect 131104 10989 131264 11023
rect 131104 10961 131139 10989
rect 131167 10961 131201 10989
rect 131229 10961 131264 10989
rect 131104 10944 131264 10961
rect 140949 11175 141259 19961
rect 140949 11147 140997 11175
rect 141025 11147 141059 11175
rect 141087 11147 141121 11175
rect 141149 11147 141183 11175
rect 141211 11147 141259 11175
rect 140949 11113 141259 11147
rect 140949 11085 140997 11113
rect 141025 11085 141059 11113
rect 141087 11085 141121 11113
rect 141149 11085 141183 11113
rect 141211 11085 141259 11113
rect 140949 11051 141259 11085
rect 140949 11023 140997 11051
rect 141025 11023 141059 11051
rect 141087 11023 141121 11051
rect 141149 11023 141183 11051
rect 141211 11023 141259 11051
rect 140949 10989 141259 11023
rect 140949 10961 140997 10989
rect 141025 10961 141059 10989
rect 141087 10961 141121 10989
rect 141149 10961 141183 10989
rect 141211 10961 141259 10989
rect 127449 5147 127497 5175
rect 127525 5147 127559 5175
rect 127587 5147 127621 5175
rect 127649 5147 127683 5175
rect 127711 5147 127759 5175
rect 127449 5113 127759 5147
rect 127449 5085 127497 5113
rect 127525 5085 127559 5113
rect 127587 5085 127621 5113
rect 127649 5085 127683 5113
rect 127711 5085 127759 5113
rect 127449 5051 127759 5085
rect 127449 5023 127497 5051
rect 127525 5023 127559 5051
rect 127587 5023 127621 5051
rect 127649 5023 127683 5051
rect 127711 5023 127759 5051
rect 127449 4989 127759 5023
rect 127449 4961 127497 4989
rect 127525 4961 127559 4989
rect 127587 4961 127621 4989
rect 127649 4961 127683 4989
rect 127711 4961 127759 4989
rect 127449 -560 127759 4961
rect 138784 5175 138944 5192
rect 138784 5147 138819 5175
rect 138847 5147 138881 5175
rect 138909 5147 138944 5175
rect 138784 5113 138944 5147
rect 138784 5085 138819 5113
rect 138847 5085 138881 5113
rect 138909 5085 138944 5113
rect 138784 5051 138944 5085
rect 138784 5023 138819 5051
rect 138847 5023 138881 5051
rect 138909 5023 138944 5051
rect 138784 4989 138944 5023
rect 138784 4961 138819 4989
rect 138847 4961 138881 4989
rect 138909 4961 138944 4989
rect 138784 4944 138944 4961
rect 127449 -588 127497 -560
rect 127525 -588 127559 -560
rect 127587 -588 127621 -560
rect 127649 -588 127683 -560
rect 127711 -588 127759 -560
rect 127449 -622 127759 -588
rect 127449 -650 127497 -622
rect 127525 -650 127559 -622
rect 127587 -650 127621 -622
rect 127649 -650 127683 -622
rect 127711 -650 127759 -622
rect 127449 -684 127759 -650
rect 127449 -712 127497 -684
rect 127525 -712 127559 -684
rect 127587 -712 127621 -684
rect 127649 -712 127683 -684
rect 127711 -712 127759 -684
rect 127449 -746 127759 -712
rect 127449 -774 127497 -746
rect 127525 -774 127559 -746
rect 127587 -774 127621 -746
rect 127649 -774 127683 -746
rect 127711 -774 127759 -746
rect 127449 -822 127759 -774
rect 140949 2175 141259 10961
rect 140949 2147 140997 2175
rect 141025 2147 141059 2175
rect 141087 2147 141121 2175
rect 141149 2147 141183 2175
rect 141211 2147 141259 2175
rect 140949 2113 141259 2147
rect 140949 2085 140997 2113
rect 141025 2085 141059 2113
rect 141087 2085 141121 2113
rect 141149 2085 141183 2113
rect 141211 2085 141259 2113
rect 140949 2051 141259 2085
rect 140949 2023 140997 2051
rect 141025 2023 141059 2051
rect 141087 2023 141121 2051
rect 141149 2023 141183 2051
rect 141211 2023 141259 2051
rect 140949 1989 141259 2023
rect 140949 1961 140997 1989
rect 141025 1961 141059 1989
rect 141087 1961 141121 1989
rect 141149 1961 141183 1989
rect 141211 1961 141259 1989
rect 140949 -80 141259 1961
rect 140949 -108 140997 -80
rect 141025 -108 141059 -80
rect 141087 -108 141121 -80
rect 141149 -108 141183 -80
rect 141211 -108 141259 -80
rect 140949 -142 141259 -108
rect 140949 -170 140997 -142
rect 141025 -170 141059 -142
rect 141087 -170 141121 -142
rect 141149 -170 141183 -142
rect 141211 -170 141259 -142
rect 140949 -204 141259 -170
rect 140949 -232 140997 -204
rect 141025 -232 141059 -204
rect 141087 -232 141121 -204
rect 141149 -232 141183 -204
rect 141211 -232 141259 -204
rect 140949 -266 141259 -232
rect 140949 -294 140997 -266
rect 141025 -294 141059 -266
rect 141087 -294 141121 -266
rect 141149 -294 141183 -266
rect 141211 -294 141259 -266
rect 140949 -822 141259 -294
rect 142809 299086 143119 299134
rect 142809 299058 142857 299086
rect 142885 299058 142919 299086
rect 142947 299058 142981 299086
rect 143009 299058 143043 299086
rect 143071 299058 143119 299086
rect 142809 299024 143119 299058
rect 142809 298996 142857 299024
rect 142885 298996 142919 299024
rect 142947 298996 142981 299024
rect 143009 298996 143043 299024
rect 143071 298996 143119 299024
rect 142809 298962 143119 298996
rect 142809 298934 142857 298962
rect 142885 298934 142919 298962
rect 142947 298934 142981 298962
rect 143009 298934 143043 298962
rect 143071 298934 143119 298962
rect 142809 298900 143119 298934
rect 142809 298872 142857 298900
rect 142885 298872 142919 298900
rect 142947 298872 142981 298900
rect 143009 298872 143043 298900
rect 143071 298872 143119 298900
rect 142809 293175 143119 298872
rect 142809 293147 142857 293175
rect 142885 293147 142919 293175
rect 142947 293147 142981 293175
rect 143009 293147 143043 293175
rect 143071 293147 143119 293175
rect 142809 293113 143119 293147
rect 142809 293085 142857 293113
rect 142885 293085 142919 293113
rect 142947 293085 142981 293113
rect 143009 293085 143043 293113
rect 143071 293085 143119 293113
rect 142809 293051 143119 293085
rect 142809 293023 142857 293051
rect 142885 293023 142919 293051
rect 142947 293023 142981 293051
rect 143009 293023 143043 293051
rect 143071 293023 143119 293051
rect 142809 292989 143119 293023
rect 142809 292961 142857 292989
rect 142885 292961 142919 292989
rect 142947 292961 142981 292989
rect 143009 292961 143043 292989
rect 143071 292961 143119 292989
rect 142809 284175 143119 292961
rect 142809 284147 142857 284175
rect 142885 284147 142919 284175
rect 142947 284147 142981 284175
rect 143009 284147 143043 284175
rect 143071 284147 143119 284175
rect 142809 284113 143119 284147
rect 142809 284085 142857 284113
rect 142885 284085 142919 284113
rect 142947 284085 142981 284113
rect 143009 284085 143043 284113
rect 143071 284085 143119 284113
rect 142809 284051 143119 284085
rect 142809 284023 142857 284051
rect 142885 284023 142919 284051
rect 142947 284023 142981 284051
rect 143009 284023 143043 284051
rect 143071 284023 143119 284051
rect 142809 283989 143119 284023
rect 142809 283961 142857 283989
rect 142885 283961 142919 283989
rect 142947 283961 142981 283989
rect 143009 283961 143043 283989
rect 143071 283961 143119 283989
rect 142809 275175 143119 283961
rect 142809 275147 142857 275175
rect 142885 275147 142919 275175
rect 142947 275147 142981 275175
rect 143009 275147 143043 275175
rect 143071 275147 143119 275175
rect 142809 275113 143119 275147
rect 142809 275085 142857 275113
rect 142885 275085 142919 275113
rect 142947 275085 142981 275113
rect 143009 275085 143043 275113
rect 143071 275085 143119 275113
rect 142809 275051 143119 275085
rect 142809 275023 142857 275051
rect 142885 275023 142919 275051
rect 142947 275023 142981 275051
rect 143009 275023 143043 275051
rect 143071 275023 143119 275051
rect 142809 274989 143119 275023
rect 142809 274961 142857 274989
rect 142885 274961 142919 274989
rect 142947 274961 142981 274989
rect 143009 274961 143043 274989
rect 143071 274961 143119 274989
rect 142809 266175 143119 274961
rect 142809 266147 142857 266175
rect 142885 266147 142919 266175
rect 142947 266147 142981 266175
rect 143009 266147 143043 266175
rect 143071 266147 143119 266175
rect 142809 266113 143119 266147
rect 142809 266085 142857 266113
rect 142885 266085 142919 266113
rect 142947 266085 142981 266113
rect 143009 266085 143043 266113
rect 143071 266085 143119 266113
rect 142809 266051 143119 266085
rect 142809 266023 142857 266051
rect 142885 266023 142919 266051
rect 142947 266023 142981 266051
rect 143009 266023 143043 266051
rect 143071 266023 143119 266051
rect 142809 265989 143119 266023
rect 142809 265961 142857 265989
rect 142885 265961 142919 265989
rect 142947 265961 142981 265989
rect 143009 265961 143043 265989
rect 143071 265961 143119 265989
rect 142809 257175 143119 265961
rect 142809 257147 142857 257175
rect 142885 257147 142919 257175
rect 142947 257147 142981 257175
rect 143009 257147 143043 257175
rect 143071 257147 143119 257175
rect 142809 257113 143119 257147
rect 142809 257085 142857 257113
rect 142885 257085 142919 257113
rect 142947 257085 142981 257113
rect 143009 257085 143043 257113
rect 143071 257085 143119 257113
rect 142809 257051 143119 257085
rect 142809 257023 142857 257051
rect 142885 257023 142919 257051
rect 142947 257023 142981 257051
rect 143009 257023 143043 257051
rect 143071 257023 143119 257051
rect 142809 256989 143119 257023
rect 142809 256961 142857 256989
rect 142885 256961 142919 256989
rect 142947 256961 142981 256989
rect 143009 256961 143043 256989
rect 143071 256961 143119 256989
rect 142809 248175 143119 256961
rect 142809 248147 142857 248175
rect 142885 248147 142919 248175
rect 142947 248147 142981 248175
rect 143009 248147 143043 248175
rect 143071 248147 143119 248175
rect 142809 248113 143119 248147
rect 142809 248085 142857 248113
rect 142885 248085 142919 248113
rect 142947 248085 142981 248113
rect 143009 248085 143043 248113
rect 143071 248085 143119 248113
rect 142809 248051 143119 248085
rect 142809 248023 142857 248051
rect 142885 248023 142919 248051
rect 142947 248023 142981 248051
rect 143009 248023 143043 248051
rect 143071 248023 143119 248051
rect 142809 247989 143119 248023
rect 142809 247961 142857 247989
rect 142885 247961 142919 247989
rect 142947 247961 142981 247989
rect 143009 247961 143043 247989
rect 143071 247961 143119 247989
rect 142809 239175 143119 247961
rect 142809 239147 142857 239175
rect 142885 239147 142919 239175
rect 142947 239147 142981 239175
rect 143009 239147 143043 239175
rect 143071 239147 143119 239175
rect 142809 239113 143119 239147
rect 142809 239085 142857 239113
rect 142885 239085 142919 239113
rect 142947 239085 142981 239113
rect 143009 239085 143043 239113
rect 143071 239085 143119 239113
rect 142809 239051 143119 239085
rect 142809 239023 142857 239051
rect 142885 239023 142919 239051
rect 142947 239023 142981 239051
rect 143009 239023 143043 239051
rect 143071 239023 143119 239051
rect 142809 238989 143119 239023
rect 142809 238961 142857 238989
rect 142885 238961 142919 238989
rect 142947 238961 142981 238989
rect 143009 238961 143043 238989
rect 143071 238961 143119 238989
rect 142809 230175 143119 238961
rect 142809 230147 142857 230175
rect 142885 230147 142919 230175
rect 142947 230147 142981 230175
rect 143009 230147 143043 230175
rect 143071 230147 143119 230175
rect 142809 230113 143119 230147
rect 142809 230085 142857 230113
rect 142885 230085 142919 230113
rect 142947 230085 142981 230113
rect 143009 230085 143043 230113
rect 143071 230085 143119 230113
rect 142809 230051 143119 230085
rect 142809 230023 142857 230051
rect 142885 230023 142919 230051
rect 142947 230023 142981 230051
rect 143009 230023 143043 230051
rect 143071 230023 143119 230051
rect 142809 229989 143119 230023
rect 142809 229961 142857 229989
rect 142885 229961 142919 229989
rect 142947 229961 142981 229989
rect 143009 229961 143043 229989
rect 143071 229961 143119 229989
rect 142809 221175 143119 229961
rect 142809 221147 142857 221175
rect 142885 221147 142919 221175
rect 142947 221147 142981 221175
rect 143009 221147 143043 221175
rect 143071 221147 143119 221175
rect 142809 221113 143119 221147
rect 142809 221085 142857 221113
rect 142885 221085 142919 221113
rect 142947 221085 142981 221113
rect 143009 221085 143043 221113
rect 143071 221085 143119 221113
rect 142809 221051 143119 221085
rect 142809 221023 142857 221051
rect 142885 221023 142919 221051
rect 142947 221023 142981 221051
rect 143009 221023 143043 221051
rect 143071 221023 143119 221051
rect 142809 220989 143119 221023
rect 142809 220961 142857 220989
rect 142885 220961 142919 220989
rect 142947 220961 142981 220989
rect 143009 220961 143043 220989
rect 143071 220961 143119 220989
rect 142809 212175 143119 220961
rect 142809 212147 142857 212175
rect 142885 212147 142919 212175
rect 142947 212147 142981 212175
rect 143009 212147 143043 212175
rect 143071 212147 143119 212175
rect 142809 212113 143119 212147
rect 142809 212085 142857 212113
rect 142885 212085 142919 212113
rect 142947 212085 142981 212113
rect 143009 212085 143043 212113
rect 143071 212085 143119 212113
rect 142809 212051 143119 212085
rect 142809 212023 142857 212051
rect 142885 212023 142919 212051
rect 142947 212023 142981 212051
rect 143009 212023 143043 212051
rect 143071 212023 143119 212051
rect 142809 211989 143119 212023
rect 142809 211961 142857 211989
rect 142885 211961 142919 211989
rect 142947 211961 142981 211989
rect 143009 211961 143043 211989
rect 143071 211961 143119 211989
rect 142809 203175 143119 211961
rect 142809 203147 142857 203175
rect 142885 203147 142919 203175
rect 142947 203147 142981 203175
rect 143009 203147 143043 203175
rect 143071 203147 143119 203175
rect 142809 203113 143119 203147
rect 142809 203085 142857 203113
rect 142885 203085 142919 203113
rect 142947 203085 142981 203113
rect 143009 203085 143043 203113
rect 143071 203085 143119 203113
rect 142809 203051 143119 203085
rect 142809 203023 142857 203051
rect 142885 203023 142919 203051
rect 142947 203023 142981 203051
rect 143009 203023 143043 203051
rect 143071 203023 143119 203051
rect 142809 202989 143119 203023
rect 142809 202961 142857 202989
rect 142885 202961 142919 202989
rect 142947 202961 142981 202989
rect 143009 202961 143043 202989
rect 143071 202961 143119 202989
rect 142809 194175 143119 202961
rect 142809 194147 142857 194175
rect 142885 194147 142919 194175
rect 142947 194147 142981 194175
rect 143009 194147 143043 194175
rect 143071 194147 143119 194175
rect 142809 194113 143119 194147
rect 142809 194085 142857 194113
rect 142885 194085 142919 194113
rect 142947 194085 142981 194113
rect 143009 194085 143043 194113
rect 143071 194085 143119 194113
rect 142809 194051 143119 194085
rect 142809 194023 142857 194051
rect 142885 194023 142919 194051
rect 142947 194023 142981 194051
rect 143009 194023 143043 194051
rect 143071 194023 143119 194051
rect 142809 193989 143119 194023
rect 142809 193961 142857 193989
rect 142885 193961 142919 193989
rect 142947 193961 142981 193989
rect 143009 193961 143043 193989
rect 143071 193961 143119 193989
rect 142809 185175 143119 193961
rect 142809 185147 142857 185175
rect 142885 185147 142919 185175
rect 142947 185147 142981 185175
rect 143009 185147 143043 185175
rect 143071 185147 143119 185175
rect 142809 185113 143119 185147
rect 142809 185085 142857 185113
rect 142885 185085 142919 185113
rect 142947 185085 142981 185113
rect 143009 185085 143043 185113
rect 143071 185085 143119 185113
rect 142809 185051 143119 185085
rect 142809 185023 142857 185051
rect 142885 185023 142919 185051
rect 142947 185023 142981 185051
rect 143009 185023 143043 185051
rect 143071 185023 143119 185051
rect 142809 184989 143119 185023
rect 142809 184961 142857 184989
rect 142885 184961 142919 184989
rect 142947 184961 142981 184989
rect 143009 184961 143043 184989
rect 143071 184961 143119 184989
rect 142809 176175 143119 184961
rect 142809 176147 142857 176175
rect 142885 176147 142919 176175
rect 142947 176147 142981 176175
rect 143009 176147 143043 176175
rect 143071 176147 143119 176175
rect 142809 176113 143119 176147
rect 142809 176085 142857 176113
rect 142885 176085 142919 176113
rect 142947 176085 142981 176113
rect 143009 176085 143043 176113
rect 143071 176085 143119 176113
rect 142809 176051 143119 176085
rect 142809 176023 142857 176051
rect 142885 176023 142919 176051
rect 142947 176023 142981 176051
rect 143009 176023 143043 176051
rect 143071 176023 143119 176051
rect 142809 175989 143119 176023
rect 142809 175961 142857 175989
rect 142885 175961 142919 175989
rect 142947 175961 142981 175989
rect 143009 175961 143043 175989
rect 143071 175961 143119 175989
rect 142809 167175 143119 175961
rect 156309 298606 156619 299134
rect 156309 298578 156357 298606
rect 156385 298578 156419 298606
rect 156447 298578 156481 298606
rect 156509 298578 156543 298606
rect 156571 298578 156619 298606
rect 156309 298544 156619 298578
rect 156309 298516 156357 298544
rect 156385 298516 156419 298544
rect 156447 298516 156481 298544
rect 156509 298516 156543 298544
rect 156571 298516 156619 298544
rect 156309 298482 156619 298516
rect 156309 298454 156357 298482
rect 156385 298454 156419 298482
rect 156447 298454 156481 298482
rect 156509 298454 156543 298482
rect 156571 298454 156619 298482
rect 156309 298420 156619 298454
rect 156309 298392 156357 298420
rect 156385 298392 156419 298420
rect 156447 298392 156481 298420
rect 156509 298392 156543 298420
rect 156571 298392 156619 298420
rect 156309 290175 156619 298392
rect 156309 290147 156357 290175
rect 156385 290147 156419 290175
rect 156447 290147 156481 290175
rect 156509 290147 156543 290175
rect 156571 290147 156619 290175
rect 156309 290113 156619 290147
rect 156309 290085 156357 290113
rect 156385 290085 156419 290113
rect 156447 290085 156481 290113
rect 156509 290085 156543 290113
rect 156571 290085 156619 290113
rect 156309 290051 156619 290085
rect 156309 290023 156357 290051
rect 156385 290023 156419 290051
rect 156447 290023 156481 290051
rect 156509 290023 156543 290051
rect 156571 290023 156619 290051
rect 156309 289989 156619 290023
rect 156309 289961 156357 289989
rect 156385 289961 156419 289989
rect 156447 289961 156481 289989
rect 156509 289961 156543 289989
rect 156571 289961 156619 289989
rect 156309 281175 156619 289961
rect 156309 281147 156357 281175
rect 156385 281147 156419 281175
rect 156447 281147 156481 281175
rect 156509 281147 156543 281175
rect 156571 281147 156619 281175
rect 156309 281113 156619 281147
rect 156309 281085 156357 281113
rect 156385 281085 156419 281113
rect 156447 281085 156481 281113
rect 156509 281085 156543 281113
rect 156571 281085 156619 281113
rect 156309 281051 156619 281085
rect 156309 281023 156357 281051
rect 156385 281023 156419 281051
rect 156447 281023 156481 281051
rect 156509 281023 156543 281051
rect 156571 281023 156619 281051
rect 156309 280989 156619 281023
rect 156309 280961 156357 280989
rect 156385 280961 156419 280989
rect 156447 280961 156481 280989
rect 156509 280961 156543 280989
rect 156571 280961 156619 280989
rect 156309 272175 156619 280961
rect 156309 272147 156357 272175
rect 156385 272147 156419 272175
rect 156447 272147 156481 272175
rect 156509 272147 156543 272175
rect 156571 272147 156619 272175
rect 156309 272113 156619 272147
rect 156309 272085 156357 272113
rect 156385 272085 156419 272113
rect 156447 272085 156481 272113
rect 156509 272085 156543 272113
rect 156571 272085 156619 272113
rect 156309 272051 156619 272085
rect 156309 272023 156357 272051
rect 156385 272023 156419 272051
rect 156447 272023 156481 272051
rect 156509 272023 156543 272051
rect 156571 272023 156619 272051
rect 156309 271989 156619 272023
rect 156309 271961 156357 271989
rect 156385 271961 156419 271989
rect 156447 271961 156481 271989
rect 156509 271961 156543 271989
rect 156571 271961 156619 271989
rect 156309 263175 156619 271961
rect 156309 263147 156357 263175
rect 156385 263147 156419 263175
rect 156447 263147 156481 263175
rect 156509 263147 156543 263175
rect 156571 263147 156619 263175
rect 156309 263113 156619 263147
rect 156309 263085 156357 263113
rect 156385 263085 156419 263113
rect 156447 263085 156481 263113
rect 156509 263085 156543 263113
rect 156571 263085 156619 263113
rect 156309 263051 156619 263085
rect 156309 263023 156357 263051
rect 156385 263023 156419 263051
rect 156447 263023 156481 263051
rect 156509 263023 156543 263051
rect 156571 263023 156619 263051
rect 156309 262989 156619 263023
rect 156309 262961 156357 262989
rect 156385 262961 156419 262989
rect 156447 262961 156481 262989
rect 156509 262961 156543 262989
rect 156571 262961 156619 262989
rect 156309 254175 156619 262961
rect 156309 254147 156357 254175
rect 156385 254147 156419 254175
rect 156447 254147 156481 254175
rect 156509 254147 156543 254175
rect 156571 254147 156619 254175
rect 156309 254113 156619 254147
rect 156309 254085 156357 254113
rect 156385 254085 156419 254113
rect 156447 254085 156481 254113
rect 156509 254085 156543 254113
rect 156571 254085 156619 254113
rect 156309 254051 156619 254085
rect 156309 254023 156357 254051
rect 156385 254023 156419 254051
rect 156447 254023 156481 254051
rect 156509 254023 156543 254051
rect 156571 254023 156619 254051
rect 156309 253989 156619 254023
rect 156309 253961 156357 253989
rect 156385 253961 156419 253989
rect 156447 253961 156481 253989
rect 156509 253961 156543 253989
rect 156571 253961 156619 253989
rect 156309 245175 156619 253961
rect 156309 245147 156357 245175
rect 156385 245147 156419 245175
rect 156447 245147 156481 245175
rect 156509 245147 156543 245175
rect 156571 245147 156619 245175
rect 156309 245113 156619 245147
rect 156309 245085 156357 245113
rect 156385 245085 156419 245113
rect 156447 245085 156481 245113
rect 156509 245085 156543 245113
rect 156571 245085 156619 245113
rect 156309 245051 156619 245085
rect 156309 245023 156357 245051
rect 156385 245023 156419 245051
rect 156447 245023 156481 245051
rect 156509 245023 156543 245051
rect 156571 245023 156619 245051
rect 156309 244989 156619 245023
rect 156309 244961 156357 244989
rect 156385 244961 156419 244989
rect 156447 244961 156481 244989
rect 156509 244961 156543 244989
rect 156571 244961 156619 244989
rect 156309 236175 156619 244961
rect 156309 236147 156357 236175
rect 156385 236147 156419 236175
rect 156447 236147 156481 236175
rect 156509 236147 156543 236175
rect 156571 236147 156619 236175
rect 156309 236113 156619 236147
rect 156309 236085 156357 236113
rect 156385 236085 156419 236113
rect 156447 236085 156481 236113
rect 156509 236085 156543 236113
rect 156571 236085 156619 236113
rect 156309 236051 156619 236085
rect 156309 236023 156357 236051
rect 156385 236023 156419 236051
rect 156447 236023 156481 236051
rect 156509 236023 156543 236051
rect 156571 236023 156619 236051
rect 156309 235989 156619 236023
rect 156309 235961 156357 235989
rect 156385 235961 156419 235989
rect 156447 235961 156481 235989
rect 156509 235961 156543 235989
rect 156571 235961 156619 235989
rect 156309 227175 156619 235961
rect 156309 227147 156357 227175
rect 156385 227147 156419 227175
rect 156447 227147 156481 227175
rect 156509 227147 156543 227175
rect 156571 227147 156619 227175
rect 156309 227113 156619 227147
rect 156309 227085 156357 227113
rect 156385 227085 156419 227113
rect 156447 227085 156481 227113
rect 156509 227085 156543 227113
rect 156571 227085 156619 227113
rect 156309 227051 156619 227085
rect 156309 227023 156357 227051
rect 156385 227023 156419 227051
rect 156447 227023 156481 227051
rect 156509 227023 156543 227051
rect 156571 227023 156619 227051
rect 156309 226989 156619 227023
rect 156309 226961 156357 226989
rect 156385 226961 156419 226989
rect 156447 226961 156481 226989
rect 156509 226961 156543 226989
rect 156571 226961 156619 226989
rect 156309 218175 156619 226961
rect 156309 218147 156357 218175
rect 156385 218147 156419 218175
rect 156447 218147 156481 218175
rect 156509 218147 156543 218175
rect 156571 218147 156619 218175
rect 156309 218113 156619 218147
rect 156309 218085 156357 218113
rect 156385 218085 156419 218113
rect 156447 218085 156481 218113
rect 156509 218085 156543 218113
rect 156571 218085 156619 218113
rect 156309 218051 156619 218085
rect 156309 218023 156357 218051
rect 156385 218023 156419 218051
rect 156447 218023 156481 218051
rect 156509 218023 156543 218051
rect 156571 218023 156619 218051
rect 156309 217989 156619 218023
rect 156309 217961 156357 217989
rect 156385 217961 156419 217989
rect 156447 217961 156481 217989
rect 156509 217961 156543 217989
rect 156571 217961 156619 217989
rect 156309 209175 156619 217961
rect 156309 209147 156357 209175
rect 156385 209147 156419 209175
rect 156447 209147 156481 209175
rect 156509 209147 156543 209175
rect 156571 209147 156619 209175
rect 156309 209113 156619 209147
rect 156309 209085 156357 209113
rect 156385 209085 156419 209113
rect 156447 209085 156481 209113
rect 156509 209085 156543 209113
rect 156571 209085 156619 209113
rect 156309 209051 156619 209085
rect 156309 209023 156357 209051
rect 156385 209023 156419 209051
rect 156447 209023 156481 209051
rect 156509 209023 156543 209051
rect 156571 209023 156619 209051
rect 156309 208989 156619 209023
rect 156309 208961 156357 208989
rect 156385 208961 156419 208989
rect 156447 208961 156481 208989
rect 156509 208961 156543 208989
rect 156571 208961 156619 208989
rect 156309 200175 156619 208961
rect 156309 200147 156357 200175
rect 156385 200147 156419 200175
rect 156447 200147 156481 200175
rect 156509 200147 156543 200175
rect 156571 200147 156619 200175
rect 156309 200113 156619 200147
rect 156309 200085 156357 200113
rect 156385 200085 156419 200113
rect 156447 200085 156481 200113
rect 156509 200085 156543 200113
rect 156571 200085 156619 200113
rect 156309 200051 156619 200085
rect 156309 200023 156357 200051
rect 156385 200023 156419 200051
rect 156447 200023 156481 200051
rect 156509 200023 156543 200051
rect 156571 200023 156619 200051
rect 156309 199989 156619 200023
rect 156309 199961 156357 199989
rect 156385 199961 156419 199989
rect 156447 199961 156481 199989
rect 156509 199961 156543 199989
rect 156571 199961 156619 199989
rect 156309 191175 156619 199961
rect 156309 191147 156357 191175
rect 156385 191147 156419 191175
rect 156447 191147 156481 191175
rect 156509 191147 156543 191175
rect 156571 191147 156619 191175
rect 156309 191113 156619 191147
rect 156309 191085 156357 191113
rect 156385 191085 156419 191113
rect 156447 191085 156481 191113
rect 156509 191085 156543 191113
rect 156571 191085 156619 191113
rect 156309 191051 156619 191085
rect 156309 191023 156357 191051
rect 156385 191023 156419 191051
rect 156447 191023 156481 191051
rect 156509 191023 156543 191051
rect 156571 191023 156619 191051
rect 156309 190989 156619 191023
rect 156309 190961 156357 190989
rect 156385 190961 156419 190989
rect 156447 190961 156481 190989
rect 156509 190961 156543 190989
rect 156571 190961 156619 190989
rect 156309 182175 156619 190961
rect 156309 182147 156357 182175
rect 156385 182147 156419 182175
rect 156447 182147 156481 182175
rect 156509 182147 156543 182175
rect 156571 182147 156619 182175
rect 156309 182113 156619 182147
rect 156309 182085 156357 182113
rect 156385 182085 156419 182113
rect 156447 182085 156481 182113
rect 156509 182085 156543 182113
rect 156571 182085 156619 182113
rect 156309 182051 156619 182085
rect 156309 182023 156357 182051
rect 156385 182023 156419 182051
rect 156447 182023 156481 182051
rect 156509 182023 156543 182051
rect 156571 182023 156619 182051
rect 156309 181989 156619 182023
rect 156309 181961 156357 181989
rect 156385 181961 156419 181989
rect 156447 181961 156481 181989
rect 156509 181961 156543 181989
rect 156571 181961 156619 181989
rect 146464 173175 146624 173192
rect 146464 173147 146499 173175
rect 146527 173147 146561 173175
rect 146589 173147 146624 173175
rect 146464 173113 146624 173147
rect 146464 173085 146499 173113
rect 146527 173085 146561 173113
rect 146589 173085 146624 173113
rect 146464 173051 146624 173085
rect 146464 173023 146499 173051
rect 146527 173023 146561 173051
rect 146589 173023 146624 173051
rect 146464 172989 146624 173023
rect 146464 172961 146499 172989
rect 146527 172961 146561 172989
rect 146589 172961 146624 172989
rect 146464 172944 146624 172961
rect 156309 173175 156619 181961
rect 156309 173147 156357 173175
rect 156385 173147 156419 173175
rect 156447 173147 156481 173175
rect 156509 173147 156543 173175
rect 156571 173147 156619 173175
rect 156309 173113 156619 173147
rect 156309 173085 156357 173113
rect 156385 173085 156419 173113
rect 156447 173085 156481 173113
rect 156509 173085 156543 173113
rect 156571 173085 156619 173113
rect 156309 173051 156619 173085
rect 156309 173023 156357 173051
rect 156385 173023 156419 173051
rect 156447 173023 156481 173051
rect 156509 173023 156543 173051
rect 156571 173023 156619 173051
rect 156309 172989 156619 173023
rect 156309 172961 156357 172989
rect 156385 172961 156419 172989
rect 156447 172961 156481 172989
rect 156509 172961 156543 172989
rect 156571 172961 156619 172989
rect 142809 167147 142857 167175
rect 142885 167147 142919 167175
rect 142947 167147 142981 167175
rect 143009 167147 143043 167175
rect 143071 167147 143119 167175
rect 142809 167113 143119 167147
rect 142809 167085 142857 167113
rect 142885 167085 142919 167113
rect 142947 167085 142981 167113
rect 143009 167085 143043 167113
rect 143071 167085 143119 167113
rect 142809 167051 143119 167085
rect 142809 167023 142857 167051
rect 142885 167023 142919 167051
rect 142947 167023 142981 167051
rect 143009 167023 143043 167051
rect 143071 167023 143119 167051
rect 142809 166989 143119 167023
rect 142809 166961 142857 166989
rect 142885 166961 142919 166989
rect 142947 166961 142981 166989
rect 143009 166961 143043 166989
rect 143071 166961 143119 166989
rect 142809 158175 143119 166961
rect 154144 167175 154304 167192
rect 154144 167147 154179 167175
rect 154207 167147 154241 167175
rect 154269 167147 154304 167175
rect 154144 167113 154304 167147
rect 154144 167085 154179 167113
rect 154207 167085 154241 167113
rect 154269 167085 154304 167113
rect 154144 167051 154304 167085
rect 154144 167023 154179 167051
rect 154207 167023 154241 167051
rect 154269 167023 154304 167051
rect 154144 166989 154304 167023
rect 154144 166961 154179 166989
rect 154207 166961 154241 166989
rect 154269 166961 154304 166989
rect 154144 166944 154304 166961
rect 146464 164175 146624 164192
rect 146464 164147 146499 164175
rect 146527 164147 146561 164175
rect 146589 164147 146624 164175
rect 146464 164113 146624 164147
rect 146464 164085 146499 164113
rect 146527 164085 146561 164113
rect 146589 164085 146624 164113
rect 146464 164051 146624 164085
rect 146464 164023 146499 164051
rect 146527 164023 146561 164051
rect 146589 164023 146624 164051
rect 146464 163989 146624 164023
rect 146464 163961 146499 163989
rect 146527 163961 146561 163989
rect 146589 163961 146624 163989
rect 146464 163944 146624 163961
rect 156309 164175 156619 172961
rect 156309 164147 156357 164175
rect 156385 164147 156419 164175
rect 156447 164147 156481 164175
rect 156509 164147 156543 164175
rect 156571 164147 156619 164175
rect 156309 164113 156619 164147
rect 156309 164085 156357 164113
rect 156385 164085 156419 164113
rect 156447 164085 156481 164113
rect 156509 164085 156543 164113
rect 156571 164085 156619 164113
rect 156309 164051 156619 164085
rect 156309 164023 156357 164051
rect 156385 164023 156419 164051
rect 156447 164023 156481 164051
rect 156509 164023 156543 164051
rect 156571 164023 156619 164051
rect 156309 163989 156619 164023
rect 156309 163961 156357 163989
rect 156385 163961 156419 163989
rect 156447 163961 156481 163989
rect 156509 163961 156543 163989
rect 156571 163961 156619 163989
rect 142809 158147 142857 158175
rect 142885 158147 142919 158175
rect 142947 158147 142981 158175
rect 143009 158147 143043 158175
rect 143071 158147 143119 158175
rect 142809 158113 143119 158147
rect 142809 158085 142857 158113
rect 142885 158085 142919 158113
rect 142947 158085 142981 158113
rect 143009 158085 143043 158113
rect 143071 158085 143119 158113
rect 142809 158051 143119 158085
rect 142809 158023 142857 158051
rect 142885 158023 142919 158051
rect 142947 158023 142981 158051
rect 143009 158023 143043 158051
rect 143071 158023 143119 158051
rect 142809 157989 143119 158023
rect 142809 157961 142857 157989
rect 142885 157961 142919 157989
rect 142947 157961 142981 157989
rect 143009 157961 143043 157989
rect 143071 157961 143119 157989
rect 142809 149175 143119 157961
rect 154144 158175 154304 158192
rect 154144 158147 154179 158175
rect 154207 158147 154241 158175
rect 154269 158147 154304 158175
rect 154144 158113 154304 158147
rect 154144 158085 154179 158113
rect 154207 158085 154241 158113
rect 154269 158085 154304 158113
rect 154144 158051 154304 158085
rect 154144 158023 154179 158051
rect 154207 158023 154241 158051
rect 154269 158023 154304 158051
rect 154144 157989 154304 158023
rect 154144 157961 154179 157989
rect 154207 157961 154241 157989
rect 154269 157961 154304 157989
rect 154144 157944 154304 157961
rect 146464 155175 146624 155192
rect 146464 155147 146499 155175
rect 146527 155147 146561 155175
rect 146589 155147 146624 155175
rect 146464 155113 146624 155147
rect 146464 155085 146499 155113
rect 146527 155085 146561 155113
rect 146589 155085 146624 155113
rect 146464 155051 146624 155085
rect 146464 155023 146499 155051
rect 146527 155023 146561 155051
rect 146589 155023 146624 155051
rect 146464 154989 146624 155023
rect 146464 154961 146499 154989
rect 146527 154961 146561 154989
rect 146589 154961 146624 154989
rect 146464 154944 146624 154961
rect 156309 155175 156619 163961
rect 156309 155147 156357 155175
rect 156385 155147 156419 155175
rect 156447 155147 156481 155175
rect 156509 155147 156543 155175
rect 156571 155147 156619 155175
rect 156309 155113 156619 155147
rect 156309 155085 156357 155113
rect 156385 155085 156419 155113
rect 156447 155085 156481 155113
rect 156509 155085 156543 155113
rect 156571 155085 156619 155113
rect 156309 155051 156619 155085
rect 156309 155023 156357 155051
rect 156385 155023 156419 155051
rect 156447 155023 156481 155051
rect 156509 155023 156543 155051
rect 156571 155023 156619 155051
rect 156309 154989 156619 155023
rect 156309 154961 156357 154989
rect 156385 154961 156419 154989
rect 156447 154961 156481 154989
rect 156509 154961 156543 154989
rect 156571 154961 156619 154989
rect 142809 149147 142857 149175
rect 142885 149147 142919 149175
rect 142947 149147 142981 149175
rect 143009 149147 143043 149175
rect 143071 149147 143119 149175
rect 142809 149113 143119 149147
rect 142809 149085 142857 149113
rect 142885 149085 142919 149113
rect 142947 149085 142981 149113
rect 143009 149085 143043 149113
rect 143071 149085 143119 149113
rect 142809 149051 143119 149085
rect 142809 149023 142857 149051
rect 142885 149023 142919 149051
rect 142947 149023 142981 149051
rect 143009 149023 143043 149051
rect 143071 149023 143119 149051
rect 142809 148989 143119 149023
rect 142809 148961 142857 148989
rect 142885 148961 142919 148989
rect 142947 148961 142981 148989
rect 143009 148961 143043 148989
rect 143071 148961 143119 148989
rect 142809 140175 143119 148961
rect 154144 149175 154304 149192
rect 154144 149147 154179 149175
rect 154207 149147 154241 149175
rect 154269 149147 154304 149175
rect 154144 149113 154304 149147
rect 154144 149085 154179 149113
rect 154207 149085 154241 149113
rect 154269 149085 154304 149113
rect 154144 149051 154304 149085
rect 154144 149023 154179 149051
rect 154207 149023 154241 149051
rect 154269 149023 154304 149051
rect 154144 148989 154304 149023
rect 154144 148961 154179 148989
rect 154207 148961 154241 148989
rect 154269 148961 154304 148989
rect 154144 148944 154304 148961
rect 146464 146175 146624 146192
rect 146464 146147 146499 146175
rect 146527 146147 146561 146175
rect 146589 146147 146624 146175
rect 146464 146113 146624 146147
rect 146464 146085 146499 146113
rect 146527 146085 146561 146113
rect 146589 146085 146624 146113
rect 146464 146051 146624 146085
rect 146464 146023 146499 146051
rect 146527 146023 146561 146051
rect 146589 146023 146624 146051
rect 146464 145989 146624 146023
rect 146464 145961 146499 145989
rect 146527 145961 146561 145989
rect 146589 145961 146624 145989
rect 146464 145944 146624 145961
rect 156309 146175 156619 154961
rect 156309 146147 156357 146175
rect 156385 146147 156419 146175
rect 156447 146147 156481 146175
rect 156509 146147 156543 146175
rect 156571 146147 156619 146175
rect 156309 146113 156619 146147
rect 156309 146085 156357 146113
rect 156385 146085 156419 146113
rect 156447 146085 156481 146113
rect 156509 146085 156543 146113
rect 156571 146085 156619 146113
rect 156309 146051 156619 146085
rect 156309 146023 156357 146051
rect 156385 146023 156419 146051
rect 156447 146023 156481 146051
rect 156509 146023 156543 146051
rect 156571 146023 156619 146051
rect 156309 145989 156619 146023
rect 156309 145961 156357 145989
rect 156385 145961 156419 145989
rect 156447 145961 156481 145989
rect 156509 145961 156543 145989
rect 156571 145961 156619 145989
rect 142809 140147 142857 140175
rect 142885 140147 142919 140175
rect 142947 140147 142981 140175
rect 143009 140147 143043 140175
rect 143071 140147 143119 140175
rect 142809 140113 143119 140147
rect 142809 140085 142857 140113
rect 142885 140085 142919 140113
rect 142947 140085 142981 140113
rect 143009 140085 143043 140113
rect 143071 140085 143119 140113
rect 142809 140051 143119 140085
rect 142809 140023 142857 140051
rect 142885 140023 142919 140051
rect 142947 140023 142981 140051
rect 143009 140023 143043 140051
rect 143071 140023 143119 140051
rect 142809 139989 143119 140023
rect 142809 139961 142857 139989
rect 142885 139961 142919 139989
rect 142947 139961 142981 139989
rect 143009 139961 143043 139989
rect 143071 139961 143119 139989
rect 142809 131175 143119 139961
rect 154144 140175 154304 140192
rect 154144 140147 154179 140175
rect 154207 140147 154241 140175
rect 154269 140147 154304 140175
rect 154144 140113 154304 140147
rect 154144 140085 154179 140113
rect 154207 140085 154241 140113
rect 154269 140085 154304 140113
rect 154144 140051 154304 140085
rect 154144 140023 154179 140051
rect 154207 140023 154241 140051
rect 154269 140023 154304 140051
rect 154144 139989 154304 140023
rect 154144 139961 154179 139989
rect 154207 139961 154241 139989
rect 154269 139961 154304 139989
rect 154144 139944 154304 139961
rect 146464 137175 146624 137192
rect 146464 137147 146499 137175
rect 146527 137147 146561 137175
rect 146589 137147 146624 137175
rect 146464 137113 146624 137147
rect 146464 137085 146499 137113
rect 146527 137085 146561 137113
rect 146589 137085 146624 137113
rect 146464 137051 146624 137085
rect 146464 137023 146499 137051
rect 146527 137023 146561 137051
rect 146589 137023 146624 137051
rect 146464 136989 146624 137023
rect 146464 136961 146499 136989
rect 146527 136961 146561 136989
rect 146589 136961 146624 136989
rect 146464 136944 146624 136961
rect 156309 137175 156619 145961
rect 156309 137147 156357 137175
rect 156385 137147 156419 137175
rect 156447 137147 156481 137175
rect 156509 137147 156543 137175
rect 156571 137147 156619 137175
rect 156309 137113 156619 137147
rect 156309 137085 156357 137113
rect 156385 137085 156419 137113
rect 156447 137085 156481 137113
rect 156509 137085 156543 137113
rect 156571 137085 156619 137113
rect 156309 137051 156619 137085
rect 156309 137023 156357 137051
rect 156385 137023 156419 137051
rect 156447 137023 156481 137051
rect 156509 137023 156543 137051
rect 156571 137023 156619 137051
rect 156309 136989 156619 137023
rect 156309 136961 156357 136989
rect 156385 136961 156419 136989
rect 156447 136961 156481 136989
rect 156509 136961 156543 136989
rect 156571 136961 156619 136989
rect 142809 131147 142857 131175
rect 142885 131147 142919 131175
rect 142947 131147 142981 131175
rect 143009 131147 143043 131175
rect 143071 131147 143119 131175
rect 142809 131113 143119 131147
rect 142809 131085 142857 131113
rect 142885 131085 142919 131113
rect 142947 131085 142981 131113
rect 143009 131085 143043 131113
rect 143071 131085 143119 131113
rect 142809 131051 143119 131085
rect 142809 131023 142857 131051
rect 142885 131023 142919 131051
rect 142947 131023 142981 131051
rect 143009 131023 143043 131051
rect 143071 131023 143119 131051
rect 142809 130989 143119 131023
rect 142809 130961 142857 130989
rect 142885 130961 142919 130989
rect 142947 130961 142981 130989
rect 143009 130961 143043 130989
rect 143071 130961 143119 130989
rect 142809 122175 143119 130961
rect 154144 131175 154304 131192
rect 154144 131147 154179 131175
rect 154207 131147 154241 131175
rect 154269 131147 154304 131175
rect 154144 131113 154304 131147
rect 154144 131085 154179 131113
rect 154207 131085 154241 131113
rect 154269 131085 154304 131113
rect 154144 131051 154304 131085
rect 154144 131023 154179 131051
rect 154207 131023 154241 131051
rect 154269 131023 154304 131051
rect 154144 130989 154304 131023
rect 154144 130961 154179 130989
rect 154207 130961 154241 130989
rect 154269 130961 154304 130989
rect 154144 130944 154304 130961
rect 146464 128175 146624 128192
rect 146464 128147 146499 128175
rect 146527 128147 146561 128175
rect 146589 128147 146624 128175
rect 146464 128113 146624 128147
rect 146464 128085 146499 128113
rect 146527 128085 146561 128113
rect 146589 128085 146624 128113
rect 146464 128051 146624 128085
rect 146464 128023 146499 128051
rect 146527 128023 146561 128051
rect 146589 128023 146624 128051
rect 146464 127989 146624 128023
rect 146464 127961 146499 127989
rect 146527 127961 146561 127989
rect 146589 127961 146624 127989
rect 146464 127944 146624 127961
rect 156309 128175 156619 136961
rect 156309 128147 156357 128175
rect 156385 128147 156419 128175
rect 156447 128147 156481 128175
rect 156509 128147 156543 128175
rect 156571 128147 156619 128175
rect 156309 128113 156619 128147
rect 156309 128085 156357 128113
rect 156385 128085 156419 128113
rect 156447 128085 156481 128113
rect 156509 128085 156543 128113
rect 156571 128085 156619 128113
rect 156309 128051 156619 128085
rect 156309 128023 156357 128051
rect 156385 128023 156419 128051
rect 156447 128023 156481 128051
rect 156509 128023 156543 128051
rect 156571 128023 156619 128051
rect 156309 127989 156619 128023
rect 156309 127961 156357 127989
rect 156385 127961 156419 127989
rect 156447 127961 156481 127989
rect 156509 127961 156543 127989
rect 156571 127961 156619 127989
rect 142809 122147 142857 122175
rect 142885 122147 142919 122175
rect 142947 122147 142981 122175
rect 143009 122147 143043 122175
rect 143071 122147 143119 122175
rect 142809 122113 143119 122147
rect 142809 122085 142857 122113
rect 142885 122085 142919 122113
rect 142947 122085 142981 122113
rect 143009 122085 143043 122113
rect 143071 122085 143119 122113
rect 142809 122051 143119 122085
rect 142809 122023 142857 122051
rect 142885 122023 142919 122051
rect 142947 122023 142981 122051
rect 143009 122023 143043 122051
rect 143071 122023 143119 122051
rect 142809 121989 143119 122023
rect 142809 121961 142857 121989
rect 142885 121961 142919 121989
rect 142947 121961 142981 121989
rect 143009 121961 143043 121989
rect 143071 121961 143119 121989
rect 142809 113175 143119 121961
rect 154144 122175 154304 122192
rect 154144 122147 154179 122175
rect 154207 122147 154241 122175
rect 154269 122147 154304 122175
rect 154144 122113 154304 122147
rect 154144 122085 154179 122113
rect 154207 122085 154241 122113
rect 154269 122085 154304 122113
rect 154144 122051 154304 122085
rect 154144 122023 154179 122051
rect 154207 122023 154241 122051
rect 154269 122023 154304 122051
rect 154144 121989 154304 122023
rect 154144 121961 154179 121989
rect 154207 121961 154241 121989
rect 154269 121961 154304 121989
rect 154144 121944 154304 121961
rect 146464 119175 146624 119192
rect 146464 119147 146499 119175
rect 146527 119147 146561 119175
rect 146589 119147 146624 119175
rect 146464 119113 146624 119147
rect 146464 119085 146499 119113
rect 146527 119085 146561 119113
rect 146589 119085 146624 119113
rect 146464 119051 146624 119085
rect 146464 119023 146499 119051
rect 146527 119023 146561 119051
rect 146589 119023 146624 119051
rect 146464 118989 146624 119023
rect 146464 118961 146499 118989
rect 146527 118961 146561 118989
rect 146589 118961 146624 118989
rect 146464 118944 146624 118961
rect 156309 119175 156619 127961
rect 156309 119147 156357 119175
rect 156385 119147 156419 119175
rect 156447 119147 156481 119175
rect 156509 119147 156543 119175
rect 156571 119147 156619 119175
rect 156309 119113 156619 119147
rect 156309 119085 156357 119113
rect 156385 119085 156419 119113
rect 156447 119085 156481 119113
rect 156509 119085 156543 119113
rect 156571 119085 156619 119113
rect 156309 119051 156619 119085
rect 156309 119023 156357 119051
rect 156385 119023 156419 119051
rect 156447 119023 156481 119051
rect 156509 119023 156543 119051
rect 156571 119023 156619 119051
rect 156309 118989 156619 119023
rect 156309 118961 156357 118989
rect 156385 118961 156419 118989
rect 156447 118961 156481 118989
rect 156509 118961 156543 118989
rect 156571 118961 156619 118989
rect 142809 113147 142857 113175
rect 142885 113147 142919 113175
rect 142947 113147 142981 113175
rect 143009 113147 143043 113175
rect 143071 113147 143119 113175
rect 142809 113113 143119 113147
rect 142809 113085 142857 113113
rect 142885 113085 142919 113113
rect 142947 113085 142981 113113
rect 143009 113085 143043 113113
rect 143071 113085 143119 113113
rect 142809 113051 143119 113085
rect 142809 113023 142857 113051
rect 142885 113023 142919 113051
rect 142947 113023 142981 113051
rect 143009 113023 143043 113051
rect 143071 113023 143119 113051
rect 142809 112989 143119 113023
rect 142809 112961 142857 112989
rect 142885 112961 142919 112989
rect 142947 112961 142981 112989
rect 143009 112961 143043 112989
rect 143071 112961 143119 112989
rect 142809 104175 143119 112961
rect 154144 113175 154304 113192
rect 154144 113147 154179 113175
rect 154207 113147 154241 113175
rect 154269 113147 154304 113175
rect 154144 113113 154304 113147
rect 154144 113085 154179 113113
rect 154207 113085 154241 113113
rect 154269 113085 154304 113113
rect 154144 113051 154304 113085
rect 154144 113023 154179 113051
rect 154207 113023 154241 113051
rect 154269 113023 154304 113051
rect 154144 112989 154304 113023
rect 154144 112961 154179 112989
rect 154207 112961 154241 112989
rect 154269 112961 154304 112989
rect 154144 112944 154304 112961
rect 146464 110175 146624 110192
rect 146464 110147 146499 110175
rect 146527 110147 146561 110175
rect 146589 110147 146624 110175
rect 146464 110113 146624 110147
rect 146464 110085 146499 110113
rect 146527 110085 146561 110113
rect 146589 110085 146624 110113
rect 146464 110051 146624 110085
rect 146464 110023 146499 110051
rect 146527 110023 146561 110051
rect 146589 110023 146624 110051
rect 146464 109989 146624 110023
rect 146464 109961 146499 109989
rect 146527 109961 146561 109989
rect 146589 109961 146624 109989
rect 146464 109944 146624 109961
rect 156309 110175 156619 118961
rect 156309 110147 156357 110175
rect 156385 110147 156419 110175
rect 156447 110147 156481 110175
rect 156509 110147 156543 110175
rect 156571 110147 156619 110175
rect 156309 110113 156619 110147
rect 156309 110085 156357 110113
rect 156385 110085 156419 110113
rect 156447 110085 156481 110113
rect 156509 110085 156543 110113
rect 156571 110085 156619 110113
rect 156309 110051 156619 110085
rect 156309 110023 156357 110051
rect 156385 110023 156419 110051
rect 156447 110023 156481 110051
rect 156509 110023 156543 110051
rect 156571 110023 156619 110051
rect 156309 109989 156619 110023
rect 156309 109961 156357 109989
rect 156385 109961 156419 109989
rect 156447 109961 156481 109989
rect 156509 109961 156543 109989
rect 156571 109961 156619 109989
rect 142809 104147 142857 104175
rect 142885 104147 142919 104175
rect 142947 104147 142981 104175
rect 143009 104147 143043 104175
rect 143071 104147 143119 104175
rect 142809 104113 143119 104147
rect 142809 104085 142857 104113
rect 142885 104085 142919 104113
rect 142947 104085 142981 104113
rect 143009 104085 143043 104113
rect 143071 104085 143119 104113
rect 142809 104051 143119 104085
rect 142809 104023 142857 104051
rect 142885 104023 142919 104051
rect 142947 104023 142981 104051
rect 143009 104023 143043 104051
rect 143071 104023 143119 104051
rect 142809 103989 143119 104023
rect 142809 103961 142857 103989
rect 142885 103961 142919 103989
rect 142947 103961 142981 103989
rect 143009 103961 143043 103989
rect 143071 103961 143119 103989
rect 142809 95175 143119 103961
rect 154144 104175 154304 104192
rect 154144 104147 154179 104175
rect 154207 104147 154241 104175
rect 154269 104147 154304 104175
rect 154144 104113 154304 104147
rect 154144 104085 154179 104113
rect 154207 104085 154241 104113
rect 154269 104085 154304 104113
rect 154144 104051 154304 104085
rect 154144 104023 154179 104051
rect 154207 104023 154241 104051
rect 154269 104023 154304 104051
rect 154144 103989 154304 104023
rect 154144 103961 154179 103989
rect 154207 103961 154241 103989
rect 154269 103961 154304 103989
rect 154144 103944 154304 103961
rect 146464 101175 146624 101192
rect 146464 101147 146499 101175
rect 146527 101147 146561 101175
rect 146589 101147 146624 101175
rect 146464 101113 146624 101147
rect 146464 101085 146499 101113
rect 146527 101085 146561 101113
rect 146589 101085 146624 101113
rect 146464 101051 146624 101085
rect 146464 101023 146499 101051
rect 146527 101023 146561 101051
rect 146589 101023 146624 101051
rect 146464 100989 146624 101023
rect 146464 100961 146499 100989
rect 146527 100961 146561 100989
rect 146589 100961 146624 100989
rect 146464 100944 146624 100961
rect 156309 101175 156619 109961
rect 156309 101147 156357 101175
rect 156385 101147 156419 101175
rect 156447 101147 156481 101175
rect 156509 101147 156543 101175
rect 156571 101147 156619 101175
rect 156309 101113 156619 101147
rect 156309 101085 156357 101113
rect 156385 101085 156419 101113
rect 156447 101085 156481 101113
rect 156509 101085 156543 101113
rect 156571 101085 156619 101113
rect 156309 101051 156619 101085
rect 156309 101023 156357 101051
rect 156385 101023 156419 101051
rect 156447 101023 156481 101051
rect 156509 101023 156543 101051
rect 156571 101023 156619 101051
rect 156309 100989 156619 101023
rect 156309 100961 156357 100989
rect 156385 100961 156419 100989
rect 156447 100961 156481 100989
rect 156509 100961 156543 100989
rect 156571 100961 156619 100989
rect 142809 95147 142857 95175
rect 142885 95147 142919 95175
rect 142947 95147 142981 95175
rect 143009 95147 143043 95175
rect 143071 95147 143119 95175
rect 142809 95113 143119 95147
rect 142809 95085 142857 95113
rect 142885 95085 142919 95113
rect 142947 95085 142981 95113
rect 143009 95085 143043 95113
rect 143071 95085 143119 95113
rect 142809 95051 143119 95085
rect 142809 95023 142857 95051
rect 142885 95023 142919 95051
rect 142947 95023 142981 95051
rect 143009 95023 143043 95051
rect 143071 95023 143119 95051
rect 142809 94989 143119 95023
rect 142809 94961 142857 94989
rect 142885 94961 142919 94989
rect 142947 94961 142981 94989
rect 143009 94961 143043 94989
rect 143071 94961 143119 94989
rect 142809 86175 143119 94961
rect 154144 95175 154304 95192
rect 154144 95147 154179 95175
rect 154207 95147 154241 95175
rect 154269 95147 154304 95175
rect 154144 95113 154304 95147
rect 154144 95085 154179 95113
rect 154207 95085 154241 95113
rect 154269 95085 154304 95113
rect 154144 95051 154304 95085
rect 154144 95023 154179 95051
rect 154207 95023 154241 95051
rect 154269 95023 154304 95051
rect 154144 94989 154304 95023
rect 154144 94961 154179 94989
rect 154207 94961 154241 94989
rect 154269 94961 154304 94989
rect 154144 94944 154304 94961
rect 146464 92175 146624 92192
rect 146464 92147 146499 92175
rect 146527 92147 146561 92175
rect 146589 92147 146624 92175
rect 146464 92113 146624 92147
rect 146464 92085 146499 92113
rect 146527 92085 146561 92113
rect 146589 92085 146624 92113
rect 146464 92051 146624 92085
rect 146464 92023 146499 92051
rect 146527 92023 146561 92051
rect 146589 92023 146624 92051
rect 146464 91989 146624 92023
rect 146464 91961 146499 91989
rect 146527 91961 146561 91989
rect 146589 91961 146624 91989
rect 146464 91944 146624 91961
rect 156309 92175 156619 100961
rect 156309 92147 156357 92175
rect 156385 92147 156419 92175
rect 156447 92147 156481 92175
rect 156509 92147 156543 92175
rect 156571 92147 156619 92175
rect 156309 92113 156619 92147
rect 156309 92085 156357 92113
rect 156385 92085 156419 92113
rect 156447 92085 156481 92113
rect 156509 92085 156543 92113
rect 156571 92085 156619 92113
rect 156309 92051 156619 92085
rect 156309 92023 156357 92051
rect 156385 92023 156419 92051
rect 156447 92023 156481 92051
rect 156509 92023 156543 92051
rect 156571 92023 156619 92051
rect 156309 91989 156619 92023
rect 156309 91961 156357 91989
rect 156385 91961 156419 91989
rect 156447 91961 156481 91989
rect 156509 91961 156543 91989
rect 156571 91961 156619 91989
rect 142809 86147 142857 86175
rect 142885 86147 142919 86175
rect 142947 86147 142981 86175
rect 143009 86147 143043 86175
rect 143071 86147 143119 86175
rect 142809 86113 143119 86147
rect 142809 86085 142857 86113
rect 142885 86085 142919 86113
rect 142947 86085 142981 86113
rect 143009 86085 143043 86113
rect 143071 86085 143119 86113
rect 142809 86051 143119 86085
rect 142809 86023 142857 86051
rect 142885 86023 142919 86051
rect 142947 86023 142981 86051
rect 143009 86023 143043 86051
rect 143071 86023 143119 86051
rect 142809 85989 143119 86023
rect 142809 85961 142857 85989
rect 142885 85961 142919 85989
rect 142947 85961 142981 85989
rect 143009 85961 143043 85989
rect 143071 85961 143119 85989
rect 142809 77175 143119 85961
rect 154144 86175 154304 86192
rect 154144 86147 154179 86175
rect 154207 86147 154241 86175
rect 154269 86147 154304 86175
rect 154144 86113 154304 86147
rect 154144 86085 154179 86113
rect 154207 86085 154241 86113
rect 154269 86085 154304 86113
rect 154144 86051 154304 86085
rect 154144 86023 154179 86051
rect 154207 86023 154241 86051
rect 154269 86023 154304 86051
rect 154144 85989 154304 86023
rect 154144 85961 154179 85989
rect 154207 85961 154241 85989
rect 154269 85961 154304 85989
rect 154144 85944 154304 85961
rect 146464 83175 146624 83192
rect 146464 83147 146499 83175
rect 146527 83147 146561 83175
rect 146589 83147 146624 83175
rect 146464 83113 146624 83147
rect 146464 83085 146499 83113
rect 146527 83085 146561 83113
rect 146589 83085 146624 83113
rect 146464 83051 146624 83085
rect 146464 83023 146499 83051
rect 146527 83023 146561 83051
rect 146589 83023 146624 83051
rect 146464 82989 146624 83023
rect 146464 82961 146499 82989
rect 146527 82961 146561 82989
rect 146589 82961 146624 82989
rect 146464 82944 146624 82961
rect 156309 83175 156619 91961
rect 156309 83147 156357 83175
rect 156385 83147 156419 83175
rect 156447 83147 156481 83175
rect 156509 83147 156543 83175
rect 156571 83147 156619 83175
rect 156309 83113 156619 83147
rect 156309 83085 156357 83113
rect 156385 83085 156419 83113
rect 156447 83085 156481 83113
rect 156509 83085 156543 83113
rect 156571 83085 156619 83113
rect 156309 83051 156619 83085
rect 156309 83023 156357 83051
rect 156385 83023 156419 83051
rect 156447 83023 156481 83051
rect 156509 83023 156543 83051
rect 156571 83023 156619 83051
rect 156309 82989 156619 83023
rect 156309 82961 156357 82989
rect 156385 82961 156419 82989
rect 156447 82961 156481 82989
rect 156509 82961 156543 82989
rect 156571 82961 156619 82989
rect 142809 77147 142857 77175
rect 142885 77147 142919 77175
rect 142947 77147 142981 77175
rect 143009 77147 143043 77175
rect 143071 77147 143119 77175
rect 142809 77113 143119 77147
rect 142809 77085 142857 77113
rect 142885 77085 142919 77113
rect 142947 77085 142981 77113
rect 143009 77085 143043 77113
rect 143071 77085 143119 77113
rect 142809 77051 143119 77085
rect 142809 77023 142857 77051
rect 142885 77023 142919 77051
rect 142947 77023 142981 77051
rect 143009 77023 143043 77051
rect 143071 77023 143119 77051
rect 142809 76989 143119 77023
rect 142809 76961 142857 76989
rect 142885 76961 142919 76989
rect 142947 76961 142981 76989
rect 143009 76961 143043 76989
rect 143071 76961 143119 76989
rect 142809 68175 143119 76961
rect 154144 77175 154304 77192
rect 154144 77147 154179 77175
rect 154207 77147 154241 77175
rect 154269 77147 154304 77175
rect 154144 77113 154304 77147
rect 154144 77085 154179 77113
rect 154207 77085 154241 77113
rect 154269 77085 154304 77113
rect 154144 77051 154304 77085
rect 154144 77023 154179 77051
rect 154207 77023 154241 77051
rect 154269 77023 154304 77051
rect 154144 76989 154304 77023
rect 154144 76961 154179 76989
rect 154207 76961 154241 76989
rect 154269 76961 154304 76989
rect 154144 76944 154304 76961
rect 146464 74175 146624 74192
rect 146464 74147 146499 74175
rect 146527 74147 146561 74175
rect 146589 74147 146624 74175
rect 146464 74113 146624 74147
rect 146464 74085 146499 74113
rect 146527 74085 146561 74113
rect 146589 74085 146624 74113
rect 146464 74051 146624 74085
rect 146464 74023 146499 74051
rect 146527 74023 146561 74051
rect 146589 74023 146624 74051
rect 146464 73989 146624 74023
rect 146464 73961 146499 73989
rect 146527 73961 146561 73989
rect 146589 73961 146624 73989
rect 146464 73944 146624 73961
rect 156309 74175 156619 82961
rect 156309 74147 156357 74175
rect 156385 74147 156419 74175
rect 156447 74147 156481 74175
rect 156509 74147 156543 74175
rect 156571 74147 156619 74175
rect 156309 74113 156619 74147
rect 156309 74085 156357 74113
rect 156385 74085 156419 74113
rect 156447 74085 156481 74113
rect 156509 74085 156543 74113
rect 156571 74085 156619 74113
rect 156309 74051 156619 74085
rect 156309 74023 156357 74051
rect 156385 74023 156419 74051
rect 156447 74023 156481 74051
rect 156509 74023 156543 74051
rect 156571 74023 156619 74051
rect 156309 73989 156619 74023
rect 156309 73961 156357 73989
rect 156385 73961 156419 73989
rect 156447 73961 156481 73989
rect 156509 73961 156543 73989
rect 156571 73961 156619 73989
rect 142809 68147 142857 68175
rect 142885 68147 142919 68175
rect 142947 68147 142981 68175
rect 143009 68147 143043 68175
rect 143071 68147 143119 68175
rect 142809 68113 143119 68147
rect 142809 68085 142857 68113
rect 142885 68085 142919 68113
rect 142947 68085 142981 68113
rect 143009 68085 143043 68113
rect 143071 68085 143119 68113
rect 142809 68051 143119 68085
rect 142809 68023 142857 68051
rect 142885 68023 142919 68051
rect 142947 68023 142981 68051
rect 143009 68023 143043 68051
rect 143071 68023 143119 68051
rect 142809 67989 143119 68023
rect 142809 67961 142857 67989
rect 142885 67961 142919 67989
rect 142947 67961 142981 67989
rect 143009 67961 143043 67989
rect 143071 67961 143119 67989
rect 142809 59175 143119 67961
rect 154144 68175 154304 68192
rect 154144 68147 154179 68175
rect 154207 68147 154241 68175
rect 154269 68147 154304 68175
rect 154144 68113 154304 68147
rect 154144 68085 154179 68113
rect 154207 68085 154241 68113
rect 154269 68085 154304 68113
rect 154144 68051 154304 68085
rect 154144 68023 154179 68051
rect 154207 68023 154241 68051
rect 154269 68023 154304 68051
rect 154144 67989 154304 68023
rect 154144 67961 154179 67989
rect 154207 67961 154241 67989
rect 154269 67961 154304 67989
rect 154144 67944 154304 67961
rect 146464 65175 146624 65192
rect 146464 65147 146499 65175
rect 146527 65147 146561 65175
rect 146589 65147 146624 65175
rect 146464 65113 146624 65147
rect 146464 65085 146499 65113
rect 146527 65085 146561 65113
rect 146589 65085 146624 65113
rect 146464 65051 146624 65085
rect 146464 65023 146499 65051
rect 146527 65023 146561 65051
rect 146589 65023 146624 65051
rect 146464 64989 146624 65023
rect 146464 64961 146499 64989
rect 146527 64961 146561 64989
rect 146589 64961 146624 64989
rect 146464 64944 146624 64961
rect 156309 65175 156619 73961
rect 156309 65147 156357 65175
rect 156385 65147 156419 65175
rect 156447 65147 156481 65175
rect 156509 65147 156543 65175
rect 156571 65147 156619 65175
rect 156309 65113 156619 65147
rect 156309 65085 156357 65113
rect 156385 65085 156419 65113
rect 156447 65085 156481 65113
rect 156509 65085 156543 65113
rect 156571 65085 156619 65113
rect 156309 65051 156619 65085
rect 156309 65023 156357 65051
rect 156385 65023 156419 65051
rect 156447 65023 156481 65051
rect 156509 65023 156543 65051
rect 156571 65023 156619 65051
rect 156309 64989 156619 65023
rect 156309 64961 156357 64989
rect 156385 64961 156419 64989
rect 156447 64961 156481 64989
rect 156509 64961 156543 64989
rect 156571 64961 156619 64989
rect 142809 59147 142857 59175
rect 142885 59147 142919 59175
rect 142947 59147 142981 59175
rect 143009 59147 143043 59175
rect 143071 59147 143119 59175
rect 142809 59113 143119 59147
rect 142809 59085 142857 59113
rect 142885 59085 142919 59113
rect 142947 59085 142981 59113
rect 143009 59085 143043 59113
rect 143071 59085 143119 59113
rect 142809 59051 143119 59085
rect 142809 59023 142857 59051
rect 142885 59023 142919 59051
rect 142947 59023 142981 59051
rect 143009 59023 143043 59051
rect 143071 59023 143119 59051
rect 142809 58989 143119 59023
rect 142809 58961 142857 58989
rect 142885 58961 142919 58989
rect 142947 58961 142981 58989
rect 143009 58961 143043 58989
rect 143071 58961 143119 58989
rect 142809 50175 143119 58961
rect 154144 59175 154304 59192
rect 154144 59147 154179 59175
rect 154207 59147 154241 59175
rect 154269 59147 154304 59175
rect 154144 59113 154304 59147
rect 154144 59085 154179 59113
rect 154207 59085 154241 59113
rect 154269 59085 154304 59113
rect 154144 59051 154304 59085
rect 154144 59023 154179 59051
rect 154207 59023 154241 59051
rect 154269 59023 154304 59051
rect 154144 58989 154304 59023
rect 154144 58961 154179 58989
rect 154207 58961 154241 58989
rect 154269 58961 154304 58989
rect 154144 58944 154304 58961
rect 146464 56175 146624 56192
rect 146464 56147 146499 56175
rect 146527 56147 146561 56175
rect 146589 56147 146624 56175
rect 146464 56113 146624 56147
rect 146464 56085 146499 56113
rect 146527 56085 146561 56113
rect 146589 56085 146624 56113
rect 146464 56051 146624 56085
rect 146464 56023 146499 56051
rect 146527 56023 146561 56051
rect 146589 56023 146624 56051
rect 146464 55989 146624 56023
rect 146464 55961 146499 55989
rect 146527 55961 146561 55989
rect 146589 55961 146624 55989
rect 146464 55944 146624 55961
rect 156309 56175 156619 64961
rect 156309 56147 156357 56175
rect 156385 56147 156419 56175
rect 156447 56147 156481 56175
rect 156509 56147 156543 56175
rect 156571 56147 156619 56175
rect 156309 56113 156619 56147
rect 156309 56085 156357 56113
rect 156385 56085 156419 56113
rect 156447 56085 156481 56113
rect 156509 56085 156543 56113
rect 156571 56085 156619 56113
rect 156309 56051 156619 56085
rect 156309 56023 156357 56051
rect 156385 56023 156419 56051
rect 156447 56023 156481 56051
rect 156509 56023 156543 56051
rect 156571 56023 156619 56051
rect 156309 55989 156619 56023
rect 156309 55961 156357 55989
rect 156385 55961 156419 55989
rect 156447 55961 156481 55989
rect 156509 55961 156543 55989
rect 156571 55961 156619 55989
rect 142809 50147 142857 50175
rect 142885 50147 142919 50175
rect 142947 50147 142981 50175
rect 143009 50147 143043 50175
rect 143071 50147 143119 50175
rect 142809 50113 143119 50147
rect 142809 50085 142857 50113
rect 142885 50085 142919 50113
rect 142947 50085 142981 50113
rect 143009 50085 143043 50113
rect 143071 50085 143119 50113
rect 142809 50051 143119 50085
rect 142809 50023 142857 50051
rect 142885 50023 142919 50051
rect 142947 50023 142981 50051
rect 143009 50023 143043 50051
rect 143071 50023 143119 50051
rect 142809 49989 143119 50023
rect 142809 49961 142857 49989
rect 142885 49961 142919 49989
rect 142947 49961 142981 49989
rect 143009 49961 143043 49989
rect 143071 49961 143119 49989
rect 142809 41175 143119 49961
rect 154144 50175 154304 50192
rect 154144 50147 154179 50175
rect 154207 50147 154241 50175
rect 154269 50147 154304 50175
rect 154144 50113 154304 50147
rect 154144 50085 154179 50113
rect 154207 50085 154241 50113
rect 154269 50085 154304 50113
rect 154144 50051 154304 50085
rect 154144 50023 154179 50051
rect 154207 50023 154241 50051
rect 154269 50023 154304 50051
rect 154144 49989 154304 50023
rect 154144 49961 154179 49989
rect 154207 49961 154241 49989
rect 154269 49961 154304 49989
rect 154144 49944 154304 49961
rect 146464 47175 146624 47192
rect 146464 47147 146499 47175
rect 146527 47147 146561 47175
rect 146589 47147 146624 47175
rect 146464 47113 146624 47147
rect 146464 47085 146499 47113
rect 146527 47085 146561 47113
rect 146589 47085 146624 47113
rect 146464 47051 146624 47085
rect 146464 47023 146499 47051
rect 146527 47023 146561 47051
rect 146589 47023 146624 47051
rect 146464 46989 146624 47023
rect 146464 46961 146499 46989
rect 146527 46961 146561 46989
rect 146589 46961 146624 46989
rect 146464 46944 146624 46961
rect 156309 47175 156619 55961
rect 156309 47147 156357 47175
rect 156385 47147 156419 47175
rect 156447 47147 156481 47175
rect 156509 47147 156543 47175
rect 156571 47147 156619 47175
rect 156309 47113 156619 47147
rect 156309 47085 156357 47113
rect 156385 47085 156419 47113
rect 156447 47085 156481 47113
rect 156509 47085 156543 47113
rect 156571 47085 156619 47113
rect 156309 47051 156619 47085
rect 156309 47023 156357 47051
rect 156385 47023 156419 47051
rect 156447 47023 156481 47051
rect 156509 47023 156543 47051
rect 156571 47023 156619 47051
rect 156309 46989 156619 47023
rect 156309 46961 156357 46989
rect 156385 46961 156419 46989
rect 156447 46961 156481 46989
rect 156509 46961 156543 46989
rect 156571 46961 156619 46989
rect 142809 41147 142857 41175
rect 142885 41147 142919 41175
rect 142947 41147 142981 41175
rect 143009 41147 143043 41175
rect 143071 41147 143119 41175
rect 142809 41113 143119 41147
rect 142809 41085 142857 41113
rect 142885 41085 142919 41113
rect 142947 41085 142981 41113
rect 143009 41085 143043 41113
rect 143071 41085 143119 41113
rect 142809 41051 143119 41085
rect 142809 41023 142857 41051
rect 142885 41023 142919 41051
rect 142947 41023 142981 41051
rect 143009 41023 143043 41051
rect 143071 41023 143119 41051
rect 142809 40989 143119 41023
rect 142809 40961 142857 40989
rect 142885 40961 142919 40989
rect 142947 40961 142981 40989
rect 143009 40961 143043 40989
rect 143071 40961 143119 40989
rect 142809 32175 143119 40961
rect 154144 41175 154304 41192
rect 154144 41147 154179 41175
rect 154207 41147 154241 41175
rect 154269 41147 154304 41175
rect 154144 41113 154304 41147
rect 154144 41085 154179 41113
rect 154207 41085 154241 41113
rect 154269 41085 154304 41113
rect 154144 41051 154304 41085
rect 154144 41023 154179 41051
rect 154207 41023 154241 41051
rect 154269 41023 154304 41051
rect 154144 40989 154304 41023
rect 154144 40961 154179 40989
rect 154207 40961 154241 40989
rect 154269 40961 154304 40989
rect 154144 40944 154304 40961
rect 146464 38175 146624 38192
rect 146464 38147 146499 38175
rect 146527 38147 146561 38175
rect 146589 38147 146624 38175
rect 146464 38113 146624 38147
rect 146464 38085 146499 38113
rect 146527 38085 146561 38113
rect 146589 38085 146624 38113
rect 146464 38051 146624 38085
rect 146464 38023 146499 38051
rect 146527 38023 146561 38051
rect 146589 38023 146624 38051
rect 146464 37989 146624 38023
rect 146464 37961 146499 37989
rect 146527 37961 146561 37989
rect 146589 37961 146624 37989
rect 146464 37944 146624 37961
rect 156309 38175 156619 46961
rect 156309 38147 156357 38175
rect 156385 38147 156419 38175
rect 156447 38147 156481 38175
rect 156509 38147 156543 38175
rect 156571 38147 156619 38175
rect 156309 38113 156619 38147
rect 156309 38085 156357 38113
rect 156385 38085 156419 38113
rect 156447 38085 156481 38113
rect 156509 38085 156543 38113
rect 156571 38085 156619 38113
rect 156309 38051 156619 38085
rect 156309 38023 156357 38051
rect 156385 38023 156419 38051
rect 156447 38023 156481 38051
rect 156509 38023 156543 38051
rect 156571 38023 156619 38051
rect 156309 37989 156619 38023
rect 156309 37961 156357 37989
rect 156385 37961 156419 37989
rect 156447 37961 156481 37989
rect 156509 37961 156543 37989
rect 156571 37961 156619 37989
rect 142809 32147 142857 32175
rect 142885 32147 142919 32175
rect 142947 32147 142981 32175
rect 143009 32147 143043 32175
rect 143071 32147 143119 32175
rect 142809 32113 143119 32147
rect 142809 32085 142857 32113
rect 142885 32085 142919 32113
rect 142947 32085 142981 32113
rect 143009 32085 143043 32113
rect 143071 32085 143119 32113
rect 142809 32051 143119 32085
rect 142809 32023 142857 32051
rect 142885 32023 142919 32051
rect 142947 32023 142981 32051
rect 143009 32023 143043 32051
rect 143071 32023 143119 32051
rect 142809 31989 143119 32023
rect 142809 31961 142857 31989
rect 142885 31961 142919 31989
rect 142947 31961 142981 31989
rect 143009 31961 143043 31989
rect 143071 31961 143119 31989
rect 142809 23175 143119 31961
rect 154144 32175 154304 32192
rect 154144 32147 154179 32175
rect 154207 32147 154241 32175
rect 154269 32147 154304 32175
rect 154144 32113 154304 32147
rect 154144 32085 154179 32113
rect 154207 32085 154241 32113
rect 154269 32085 154304 32113
rect 154144 32051 154304 32085
rect 154144 32023 154179 32051
rect 154207 32023 154241 32051
rect 154269 32023 154304 32051
rect 154144 31989 154304 32023
rect 154144 31961 154179 31989
rect 154207 31961 154241 31989
rect 154269 31961 154304 31989
rect 154144 31944 154304 31961
rect 146464 29175 146624 29192
rect 146464 29147 146499 29175
rect 146527 29147 146561 29175
rect 146589 29147 146624 29175
rect 146464 29113 146624 29147
rect 146464 29085 146499 29113
rect 146527 29085 146561 29113
rect 146589 29085 146624 29113
rect 146464 29051 146624 29085
rect 146464 29023 146499 29051
rect 146527 29023 146561 29051
rect 146589 29023 146624 29051
rect 146464 28989 146624 29023
rect 146464 28961 146499 28989
rect 146527 28961 146561 28989
rect 146589 28961 146624 28989
rect 146464 28944 146624 28961
rect 156309 29175 156619 37961
rect 156309 29147 156357 29175
rect 156385 29147 156419 29175
rect 156447 29147 156481 29175
rect 156509 29147 156543 29175
rect 156571 29147 156619 29175
rect 156309 29113 156619 29147
rect 156309 29085 156357 29113
rect 156385 29085 156419 29113
rect 156447 29085 156481 29113
rect 156509 29085 156543 29113
rect 156571 29085 156619 29113
rect 156309 29051 156619 29085
rect 156309 29023 156357 29051
rect 156385 29023 156419 29051
rect 156447 29023 156481 29051
rect 156509 29023 156543 29051
rect 156571 29023 156619 29051
rect 156309 28989 156619 29023
rect 156309 28961 156357 28989
rect 156385 28961 156419 28989
rect 156447 28961 156481 28989
rect 156509 28961 156543 28989
rect 156571 28961 156619 28989
rect 142809 23147 142857 23175
rect 142885 23147 142919 23175
rect 142947 23147 142981 23175
rect 143009 23147 143043 23175
rect 143071 23147 143119 23175
rect 142809 23113 143119 23147
rect 142809 23085 142857 23113
rect 142885 23085 142919 23113
rect 142947 23085 142981 23113
rect 143009 23085 143043 23113
rect 143071 23085 143119 23113
rect 142809 23051 143119 23085
rect 142809 23023 142857 23051
rect 142885 23023 142919 23051
rect 142947 23023 142981 23051
rect 143009 23023 143043 23051
rect 143071 23023 143119 23051
rect 142809 22989 143119 23023
rect 142809 22961 142857 22989
rect 142885 22961 142919 22989
rect 142947 22961 142981 22989
rect 143009 22961 143043 22989
rect 143071 22961 143119 22989
rect 142809 14175 143119 22961
rect 154144 23175 154304 23192
rect 154144 23147 154179 23175
rect 154207 23147 154241 23175
rect 154269 23147 154304 23175
rect 154144 23113 154304 23147
rect 154144 23085 154179 23113
rect 154207 23085 154241 23113
rect 154269 23085 154304 23113
rect 154144 23051 154304 23085
rect 154144 23023 154179 23051
rect 154207 23023 154241 23051
rect 154269 23023 154304 23051
rect 154144 22989 154304 23023
rect 154144 22961 154179 22989
rect 154207 22961 154241 22989
rect 154269 22961 154304 22989
rect 154144 22944 154304 22961
rect 146464 20175 146624 20192
rect 146464 20147 146499 20175
rect 146527 20147 146561 20175
rect 146589 20147 146624 20175
rect 146464 20113 146624 20147
rect 146464 20085 146499 20113
rect 146527 20085 146561 20113
rect 146589 20085 146624 20113
rect 146464 20051 146624 20085
rect 146464 20023 146499 20051
rect 146527 20023 146561 20051
rect 146589 20023 146624 20051
rect 146464 19989 146624 20023
rect 146464 19961 146499 19989
rect 146527 19961 146561 19989
rect 146589 19961 146624 19989
rect 146464 19944 146624 19961
rect 156309 20175 156619 28961
rect 156309 20147 156357 20175
rect 156385 20147 156419 20175
rect 156447 20147 156481 20175
rect 156509 20147 156543 20175
rect 156571 20147 156619 20175
rect 156309 20113 156619 20147
rect 156309 20085 156357 20113
rect 156385 20085 156419 20113
rect 156447 20085 156481 20113
rect 156509 20085 156543 20113
rect 156571 20085 156619 20113
rect 156309 20051 156619 20085
rect 156309 20023 156357 20051
rect 156385 20023 156419 20051
rect 156447 20023 156481 20051
rect 156509 20023 156543 20051
rect 156571 20023 156619 20051
rect 156309 19989 156619 20023
rect 156309 19961 156357 19989
rect 156385 19961 156419 19989
rect 156447 19961 156481 19989
rect 156509 19961 156543 19989
rect 156571 19961 156619 19989
rect 142809 14147 142857 14175
rect 142885 14147 142919 14175
rect 142947 14147 142981 14175
rect 143009 14147 143043 14175
rect 143071 14147 143119 14175
rect 142809 14113 143119 14147
rect 142809 14085 142857 14113
rect 142885 14085 142919 14113
rect 142947 14085 142981 14113
rect 143009 14085 143043 14113
rect 143071 14085 143119 14113
rect 142809 14051 143119 14085
rect 142809 14023 142857 14051
rect 142885 14023 142919 14051
rect 142947 14023 142981 14051
rect 143009 14023 143043 14051
rect 143071 14023 143119 14051
rect 142809 13989 143119 14023
rect 142809 13961 142857 13989
rect 142885 13961 142919 13989
rect 142947 13961 142981 13989
rect 143009 13961 143043 13989
rect 143071 13961 143119 13989
rect 142809 5175 143119 13961
rect 154144 14175 154304 14192
rect 154144 14147 154179 14175
rect 154207 14147 154241 14175
rect 154269 14147 154304 14175
rect 154144 14113 154304 14147
rect 154144 14085 154179 14113
rect 154207 14085 154241 14113
rect 154269 14085 154304 14113
rect 154144 14051 154304 14085
rect 154144 14023 154179 14051
rect 154207 14023 154241 14051
rect 154269 14023 154304 14051
rect 154144 13989 154304 14023
rect 154144 13961 154179 13989
rect 154207 13961 154241 13989
rect 154269 13961 154304 13989
rect 154144 13944 154304 13961
rect 146464 11175 146624 11192
rect 146464 11147 146499 11175
rect 146527 11147 146561 11175
rect 146589 11147 146624 11175
rect 146464 11113 146624 11147
rect 146464 11085 146499 11113
rect 146527 11085 146561 11113
rect 146589 11085 146624 11113
rect 146464 11051 146624 11085
rect 146464 11023 146499 11051
rect 146527 11023 146561 11051
rect 146589 11023 146624 11051
rect 146464 10989 146624 11023
rect 146464 10961 146499 10989
rect 146527 10961 146561 10989
rect 146589 10961 146624 10989
rect 146464 10944 146624 10961
rect 156309 11175 156619 19961
rect 156309 11147 156357 11175
rect 156385 11147 156419 11175
rect 156447 11147 156481 11175
rect 156509 11147 156543 11175
rect 156571 11147 156619 11175
rect 156309 11113 156619 11147
rect 156309 11085 156357 11113
rect 156385 11085 156419 11113
rect 156447 11085 156481 11113
rect 156509 11085 156543 11113
rect 156571 11085 156619 11113
rect 156309 11051 156619 11085
rect 156309 11023 156357 11051
rect 156385 11023 156419 11051
rect 156447 11023 156481 11051
rect 156509 11023 156543 11051
rect 156571 11023 156619 11051
rect 156309 10989 156619 11023
rect 156309 10961 156357 10989
rect 156385 10961 156419 10989
rect 156447 10961 156481 10989
rect 156509 10961 156543 10989
rect 156571 10961 156619 10989
rect 142809 5147 142857 5175
rect 142885 5147 142919 5175
rect 142947 5147 142981 5175
rect 143009 5147 143043 5175
rect 143071 5147 143119 5175
rect 142809 5113 143119 5147
rect 142809 5085 142857 5113
rect 142885 5085 142919 5113
rect 142947 5085 142981 5113
rect 143009 5085 143043 5113
rect 143071 5085 143119 5113
rect 142809 5051 143119 5085
rect 142809 5023 142857 5051
rect 142885 5023 142919 5051
rect 142947 5023 142981 5051
rect 143009 5023 143043 5051
rect 143071 5023 143119 5051
rect 142809 4989 143119 5023
rect 142809 4961 142857 4989
rect 142885 4961 142919 4989
rect 142947 4961 142981 4989
rect 143009 4961 143043 4989
rect 143071 4961 143119 4989
rect 142809 -560 143119 4961
rect 154144 5175 154304 5192
rect 154144 5147 154179 5175
rect 154207 5147 154241 5175
rect 154269 5147 154304 5175
rect 154144 5113 154304 5147
rect 154144 5085 154179 5113
rect 154207 5085 154241 5113
rect 154269 5085 154304 5113
rect 154144 5051 154304 5085
rect 154144 5023 154179 5051
rect 154207 5023 154241 5051
rect 154269 5023 154304 5051
rect 154144 4989 154304 5023
rect 154144 4961 154179 4989
rect 154207 4961 154241 4989
rect 154269 4961 154304 4989
rect 154144 4944 154304 4961
rect 142809 -588 142857 -560
rect 142885 -588 142919 -560
rect 142947 -588 142981 -560
rect 143009 -588 143043 -560
rect 143071 -588 143119 -560
rect 142809 -622 143119 -588
rect 142809 -650 142857 -622
rect 142885 -650 142919 -622
rect 142947 -650 142981 -622
rect 143009 -650 143043 -622
rect 143071 -650 143119 -622
rect 142809 -684 143119 -650
rect 142809 -712 142857 -684
rect 142885 -712 142919 -684
rect 142947 -712 142981 -684
rect 143009 -712 143043 -684
rect 143071 -712 143119 -684
rect 142809 -746 143119 -712
rect 142809 -774 142857 -746
rect 142885 -774 142919 -746
rect 142947 -774 142981 -746
rect 143009 -774 143043 -746
rect 143071 -774 143119 -746
rect 142809 -822 143119 -774
rect 156309 2175 156619 10961
rect 156309 2147 156357 2175
rect 156385 2147 156419 2175
rect 156447 2147 156481 2175
rect 156509 2147 156543 2175
rect 156571 2147 156619 2175
rect 156309 2113 156619 2147
rect 156309 2085 156357 2113
rect 156385 2085 156419 2113
rect 156447 2085 156481 2113
rect 156509 2085 156543 2113
rect 156571 2085 156619 2113
rect 156309 2051 156619 2085
rect 156309 2023 156357 2051
rect 156385 2023 156419 2051
rect 156447 2023 156481 2051
rect 156509 2023 156543 2051
rect 156571 2023 156619 2051
rect 156309 1989 156619 2023
rect 156309 1961 156357 1989
rect 156385 1961 156419 1989
rect 156447 1961 156481 1989
rect 156509 1961 156543 1989
rect 156571 1961 156619 1989
rect 156309 -80 156619 1961
rect 156309 -108 156357 -80
rect 156385 -108 156419 -80
rect 156447 -108 156481 -80
rect 156509 -108 156543 -80
rect 156571 -108 156619 -80
rect 156309 -142 156619 -108
rect 156309 -170 156357 -142
rect 156385 -170 156419 -142
rect 156447 -170 156481 -142
rect 156509 -170 156543 -142
rect 156571 -170 156619 -142
rect 156309 -204 156619 -170
rect 156309 -232 156357 -204
rect 156385 -232 156419 -204
rect 156447 -232 156481 -204
rect 156509 -232 156543 -204
rect 156571 -232 156619 -204
rect 156309 -266 156619 -232
rect 156309 -294 156357 -266
rect 156385 -294 156419 -266
rect 156447 -294 156481 -266
rect 156509 -294 156543 -266
rect 156571 -294 156619 -266
rect 156309 -822 156619 -294
rect 158169 299086 158479 299134
rect 158169 299058 158217 299086
rect 158245 299058 158279 299086
rect 158307 299058 158341 299086
rect 158369 299058 158403 299086
rect 158431 299058 158479 299086
rect 158169 299024 158479 299058
rect 158169 298996 158217 299024
rect 158245 298996 158279 299024
rect 158307 298996 158341 299024
rect 158369 298996 158403 299024
rect 158431 298996 158479 299024
rect 158169 298962 158479 298996
rect 158169 298934 158217 298962
rect 158245 298934 158279 298962
rect 158307 298934 158341 298962
rect 158369 298934 158403 298962
rect 158431 298934 158479 298962
rect 158169 298900 158479 298934
rect 158169 298872 158217 298900
rect 158245 298872 158279 298900
rect 158307 298872 158341 298900
rect 158369 298872 158403 298900
rect 158431 298872 158479 298900
rect 158169 293175 158479 298872
rect 158169 293147 158217 293175
rect 158245 293147 158279 293175
rect 158307 293147 158341 293175
rect 158369 293147 158403 293175
rect 158431 293147 158479 293175
rect 158169 293113 158479 293147
rect 158169 293085 158217 293113
rect 158245 293085 158279 293113
rect 158307 293085 158341 293113
rect 158369 293085 158403 293113
rect 158431 293085 158479 293113
rect 158169 293051 158479 293085
rect 158169 293023 158217 293051
rect 158245 293023 158279 293051
rect 158307 293023 158341 293051
rect 158369 293023 158403 293051
rect 158431 293023 158479 293051
rect 158169 292989 158479 293023
rect 158169 292961 158217 292989
rect 158245 292961 158279 292989
rect 158307 292961 158341 292989
rect 158369 292961 158403 292989
rect 158431 292961 158479 292989
rect 158169 284175 158479 292961
rect 158169 284147 158217 284175
rect 158245 284147 158279 284175
rect 158307 284147 158341 284175
rect 158369 284147 158403 284175
rect 158431 284147 158479 284175
rect 158169 284113 158479 284147
rect 158169 284085 158217 284113
rect 158245 284085 158279 284113
rect 158307 284085 158341 284113
rect 158369 284085 158403 284113
rect 158431 284085 158479 284113
rect 158169 284051 158479 284085
rect 158169 284023 158217 284051
rect 158245 284023 158279 284051
rect 158307 284023 158341 284051
rect 158369 284023 158403 284051
rect 158431 284023 158479 284051
rect 158169 283989 158479 284023
rect 158169 283961 158217 283989
rect 158245 283961 158279 283989
rect 158307 283961 158341 283989
rect 158369 283961 158403 283989
rect 158431 283961 158479 283989
rect 158169 275175 158479 283961
rect 158169 275147 158217 275175
rect 158245 275147 158279 275175
rect 158307 275147 158341 275175
rect 158369 275147 158403 275175
rect 158431 275147 158479 275175
rect 158169 275113 158479 275147
rect 158169 275085 158217 275113
rect 158245 275085 158279 275113
rect 158307 275085 158341 275113
rect 158369 275085 158403 275113
rect 158431 275085 158479 275113
rect 158169 275051 158479 275085
rect 158169 275023 158217 275051
rect 158245 275023 158279 275051
rect 158307 275023 158341 275051
rect 158369 275023 158403 275051
rect 158431 275023 158479 275051
rect 158169 274989 158479 275023
rect 158169 274961 158217 274989
rect 158245 274961 158279 274989
rect 158307 274961 158341 274989
rect 158369 274961 158403 274989
rect 158431 274961 158479 274989
rect 158169 266175 158479 274961
rect 158169 266147 158217 266175
rect 158245 266147 158279 266175
rect 158307 266147 158341 266175
rect 158369 266147 158403 266175
rect 158431 266147 158479 266175
rect 158169 266113 158479 266147
rect 158169 266085 158217 266113
rect 158245 266085 158279 266113
rect 158307 266085 158341 266113
rect 158369 266085 158403 266113
rect 158431 266085 158479 266113
rect 158169 266051 158479 266085
rect 158169 266023 158217 266051
rect 158245 266023 158279 266051
rect 158307 266023 158341 266051
rect 158369 266023 158403 266051
rect 158431 266023 158479 266051
rect 158169 265989 158479 266023
rect 158169 265961 158217 265989
rect 158245 265961 158279 265989
rect 158307 265961 158341 265989
rect 158369 265961 158403 265989
rect 158431 265961 158479 265989
rect 158169 257175 158479 265961
rect 158169 257147 158217 257175
rect 158245 257147 158279 257175
rect 158307 257147 158341 257175
rect 158369 257147 158403 257175
rect 158431 257147 158479 257175
rect 158169 257113 158479 257147
rect 158169 257085 158217 257113
rect 158245 257085 158279 257113
rect 158307 257085 158341 257113
rect 158369 257085 158403 257113
rect 158431 257085 158479 257113
rect 158169 257051 158479 257085
rect 158169 257023 158217 257051
rect 158245 257023 158279 257051
rect 158307 257023 158341 257051
rect 158369 257023 158403 257051
rect 158431 257023 158479 257051
rect 158169 256989 158479 257023
rect 158169 256961 158217 256989
rect 158245 256961 158279 256989
rect 158307 256961 158341 256989
rect 158369 256961 158403 256989
rect 158431 256961 158479 256989
rect 158169 248175 158479 256961
rect 158169 248147 158217 248175
rect 158245 248147 158279 248175
rect 158307 248147 158341 248175
rect 158369 248147 158403 248175
rect 158431 248147 158479 248175
rect 158169 248113 158479 248147
rect 158169 248085 158217 248113
rect 158245 248085 158279 248113
rect 158307 248085 158341 248113
rect 158369 248085 158403 248113
rect 158431 248085 158479 248113
rect 158169 248051 158479 248085
rect 158169 248023 158217 248051
rect 158245 248023 158279 248051
rect 158307 248023 158341 248051
rect 158369 248023 158403 248051
rect 158431 248023 158479 248051
rect 158169 247989 158479 248023
rect 158169 247961 158217 247989
rect 158245 247961 158279 247989
rect 158307 247961 158341 247989
rect 158369 247961 158403 247989
rect 158431 247961 158479 247989
rect 158169 239175 158479 247961
rect 158169 239147 158217 239175
rect 158245 239147 158279 239175
rect 158307 239147 158341 239175
rect 158369 239147 158403 239175
rect 158431 239147 158479 239175
rect 158169 239113 158479 239147
rect 158169 239085 158217 239113
rect 158245 239085 158279 239113
rect 158307 239085 158341 239113
rect 158369 239085 158403 239113
rect 158431 239085 158479 239113
rect 158169 239051 158479 239085
rect 158169 239023 158217 239051
rect 158245 239023 158279 239051
rect 158307 239023 158341 239051
rect 158369 239023 158403 239051
rect 158431 239023 158479 239051
rect 158169 238989 158479 239023
rect 158169 238961 158217 238989
rect 158245 238961 158279 238989
rect 158307 238961 158341 238989
rect 158369 238961 158403 238989
rect 158431 238961 158479 238989
rect 158169 230175 158479 238961
rect 158169 230147 158217 230175
rect 158245 230147 158279 230175
rect 158307 230147 158341 230175
rect 158369 230147 158403 230175
rect 158431 230147 158479 230175
rect 158169 230113 158479 230147
rect 158169 230085 158217 230113
rect 158245 230085 158279 230113
rect 158307 230085 158341 230113
rect 158369 230085 158403 230113
rect 158431 230085 158479 230113
rect 158169 230051 158479 230085
rect 158169 230023 158217 230051
rect 158245 230023 158279 230051
rect 158307 230023 158341 230051
rect 158369 230023 158403 230051
rect 158431 230023 158479 230051
rect 158169 229989 158479 230023
rect 158169 229961 158217 229989
rect 158245 229961 158279 229989
rect 158307 229961 158341 229989
rect 158369 229961 158403 229989
rect 158431 229961 158479 229989
rect 158169 221175 158479 229961
rect 158169 221147 158217 221175
rect 158245 221147 158279 221175
rect 158307 221147 158341 221175
rect 158369 221147 158403 221175
rect 158431 221147 158479 221175
rect 158169 221113 158479 221147
rect 158169 221085 158217 221113
rect 158245 221085 158279 221113
rect 158307 221085 158341 221113
rect 158369 221085 158403 221113
rect 158431 221085 158479 221113
rect 158169 221051 158479 221085
rect 158169 221023 158217 221051
rect 158245 221023 158279 221051
rect 158307 221023 158341 221051
rect 158369 221023 158403 221051
rect 158431 221023 158479 221051
rect 158169 220989 158479 221023
rect 158169 220961 158217 220989
rect 158245 220961 158279 220989
rect 158307 220961 158341 220989
rect 158369 220961 158403 220989
rect 158431 220961 158479 220989
rect 158169 212175 158479 220961
rect 158169 212147 158217 212175
rect 158245 212147 158279 212175
rect 158307 212147 158341 212175
rect 158369 212147 158403 212175
rect 158431 212147 158479 212175
rect 158169 212113 158479 212147
rect 158169 212085 158217 212113
rect 158245 212085 158279 212113
rect 158307 212085 158341 212113
rect 158369 212085 158403 212113
rect 158431 212085 158479 212113
rect 158169 212051 158479 212085
rect 158169 212023 158217 212051
rect 158245 212023 158279 212051
rect 158307 212023 158341 212051
rect 158369 212023 158403 212051
rect 158431 212023 158479 212051
rect 158169 211989 158479 212023
rect 158169 211961 158217 211989
rect 158245 211961 158279 211989
rect 158307 211961 158341 211989
rect 158369 211961 158403 211989
rect 158431 211961 158479 211989
rect 158169 203175 158479 211961
rect 158169 203147 158217 203175
rect 158245 203147 158279 203175
rect 158307 203147 158341 203175
rect 158369 203147 158403 203175
rect 158431 203147 158479 203175
rect 158169 203113 158479 203147
rect 158169 203085 158217 203113
rect 158245 203085 158279 203113
rect 158307 203085 158341 203113
rect 158369 203085 158403 203113
rect 158431 203085 158479 203113
rect 158169 203051 158479 203085
rect 158169 203023 158217 203051
rect 158245 203023 158279 203051
rect 158307 203023 158341 203051
rect 158369 203023 158403 203051
rect 158431 203023 158479 203051
rect 158169 202989 158479 203023
rect 158169 202961 158217 202989
rect 158245 202961 158279 202989
rect 158307 202961 158341 202989
rect 158369 202961 158403 202989
rect 158431 202961 158479 202989
rect 158169 194175 158479 202961
rect 158169 194147 158217 194175
rect 158245 194147 158279 194175
rect 158307 194147 158341 194175
rect 158369 194147 158403 194175
rect 158431 194147 158479 194175
rect 158169 194113 158479 194147
rect 158169 194085 158217 194113
rect 158245 194085 158279 194113
rect 158307 194085 158341 194113
rect 158369 194085 158403 194113
rect 158431 194085 158479 194113
rect 158169 194051 158479 194085
rect 158169 194023 158217 194051
rect 158245 194023 158279 194051
rect 158307 194023 158341 194051
rect 158369 194023 158403 194051
rect 158431 194023 158479 194051
rect 158169 193989 158479 194023
rect 158169 193961 158217 193989
rect 158245 193961 158279 193989
rect 158307 193961 158341 193989
rect 158369 193961 158403 193989
rect 158431 193961 158479 193989
rect 158169 185175 158479 193961
rect 158169 185147 158217 185175
rect 158245 185147 158279 185175
rect 158307 185147 158341 185175
rect 158369 185147 158403 185175
rect 158431 185147 158479 185175
rect 158169 185113 158479 185147
rect 158169 185085 158217 185113
rect 158245 185085 158279 185113
rect 158307 185085 158341 185113
rect 158369 185085 158403 185113
rect 158431 185085 158479 185113
rect 158169 185051 158479 185085
rect 158169 185023 158217 185051
rect 158245 185023 158279 185051
rect 158307 185023 158341 185051
rect 158369 185023 158403 185051
rect 158431 185023 158479 185051
rect 158169 184989 158479 185023
rect 158169 184961 158217 184989
rect 158245 184961 158279 184989
rect 158307 184961 158341 184989
rect 158369 184961 158403 184989
rect 158431 184961 158479 184989
rect 158169 176175 158479 184961
rect 158169 176147 158217 176175
rect 158245 176147 158279 176175
rect 158307 176147 158341 176175
rect 158369 176147 158403 176175
rect 158431 176147 158479 176175
rect 158169 176113 158479 176147
rect 158169 176085 158217 176113
rect 158245 176085 158279 176113
rect 158307 176085 158341 176113
rect 158369 176085 158403 176113
rect 158431 176085 158479 176113
rect 158169 176051 158479 176085
rect 158169 176023 158217 176051
rect 158245 176023 158279 176051
rect 158307 176023 158341 176051
rect 158369 176023 158403 176051
rect 158431 176023 158479 176051
rect 158169 175989 158479 176023
rect 158169 175961 158217 175989
rect 158245 175961 158279 175989
rect 158307 175961 158341 175989
rect 158369 175961 158403 175989
rect 158431 175961 158479 175989
rect 158169 167175 158479 175961
rect 171669 298606 171979 299134
rect 171669 298578 171717 298606
rect 171745 298578 171779 298606
rect 171807 298578 171841 298606
rect 171869 298578 171903 298606
rect 171931 298578 171979 298606
rect 171669 298544 171979 298578
rect 171669 298516 171717 298544
rect 171745 298516 171779 298544
rect 171807 298516 171841 298544
rect 171869 298516 171903 298544
rect 171931 298516 171979 298544
rect 171669 298482 171979 298516
rect 171669 298454 171717 298482
rect 171745 298454 171779 298482
rect 171807 298454 171841 298482
rect 171869 298454 171903 298482
rect 171931 298454 171979 298482
rect 171669 298420 171979 298454
rect 171669 298392 171717 298420
rect 171745 298392 171779 298420
rect 171807 298392 171841 298420
rect 171869 298392 171903 298420
rect 171931 298392 171979 298420
rect 171669 290175 171979 298392
rect 171669 290147 171717 290175
rect 171745 290147 171779 290175
rect 171807 290147 171841 290175
rect 171869 290147 171903 290175
rect 171931 290147 171979 290175
rect 171669 290113 171979 290147
rect 171669 290085 171717 290113
rect 171745 290085 171779 290113
rect 171807 290085 171841 290113
rect 171869 290085 171903 290113
rect 171931 290085 171979 290113
rect 171669 290051 171979 290085
rect 171669 290023 171717 290051
rect 171745 290023 171779 290051
rect 171807 290023 171841 290051
rect 171869 290023 171903 290051
rect 171931 290023 171979 290051
rect 171669 289989 171979 290023
rect 171669 289961 171717 289989
rect 171745 289961 171779 289989
rect 171807 289961 171841 289989
rect 171869 289961 171903 289989
rect 171931 289961 171979 289989
rect 171669 281175 171979 289961
rect 171669 281147 171717 281175
rect 171745 281147 171779 281175
rect 171807 281147 171841 281175
rect 171869 281147 171903 281175
rect 171931 281147 171979 281175
rect 171669 281113 171979 281147
rect 171669 281085 171717 281113
rect 171745 281085 171779 281113
rect 171807 281085 171841 281113
rect 171869 281085 171903 281113
rect 171931 281085 171979 281113
rect 171669 281051 171979 281085
rect 171669 281023 171717 281051
rect 171745 281023 171779 281051
rect 171807 281023 171841 281051
rect 171869 281023 171903 281051
rect 171931 281023 171979 281051
rect 171669 280989 171979 281023
rect 171669 280961 171717 280989
rect 171745 280961 171779 280989
rect 171807 280961 171841 280989
rect 171869 280961 171903 280989
rect 171931 280961 171979 280989
rect 171669 272175 171979 280961
rect 171669 272147 171717 272175
rect 171745 272147 171779 272175
rect 171807 272147 171841 272175
rect 171869 272147 171903 272175
rect 171931 272147 171979 272175
rect 171669 272113 171979 272147
rect 171669 272085 171717 272113
rect 171745 272085 171779 272113
rect 171807 272085 171841 272113
rect 171869 272085 171903 272113
rect 171931 272085 171979 272113
rect 171669 272051 171979 272085
rect 171669 272023 171717 272051
rect 171745 272023 171779 272051
rect 171807 272023 171841 272051
rect 171869 272023 171903 272051
rect 171931 272023 171979 272051
rect 171669 271989 171979 272023
rect 171669 271961 171717 271989
rect 171745 271961 171779 271989
rect 171807 271961 171841 271989
rect 171869 271961 171903 271989
rect 171931 271961 171979 271989
rect 171669 263175 171979 271961
rect 171669 263147 171717 263175
rect 171745 263147 171779 263175
rect 171807 263147 171841 263175
rect 171869 263147 171903 263175
rect 171931 263147 171979 263175
rect 171669 263113 171979 263147
rect 171669 263085 171717 263113
rect 171745 263085 171779 263113
rect 171807 263085 171841 263113
rect 171869 263085 171903 263113
rect 171931 263085 171979 263113
rect 171669 263051 171979 263085
rect 171669 263023 171717 263051
rect 171745 263023 171779 263051
rect 171807 263023 171841 263051
rect 171869 263023 171903 263051
rect 171931 263023 171979 263051
rect 171669 262989 171979 263023
rect 171669 262961 171717 262989
rect 171745 262961 171779 262989
rect 171807 262961 171841 262989
rect 171869 262961 171903 262989
rect 171931 262961 171979 262989
rect 171669 254175 171979 262961
rect 171669 254147 171717 254175
rect 171745 254147 171779 254175
rect 171807 254147 171841 254175
rect 171869 254147 171903 254175
rect 171931 254147 171979 254175
rect 171669 254113 171979 254147
rect 171669 254085 171717 254113
rect 171745 254085 171779 254113
rect 171807 254085 171841 254113
rect 171869 254085 171903 254113
rect 171931 254085 171979 254113
rect 171669 254051 171979 254085
rect 171669 254023 171717 254051
rect 171745 254023 171779 254051
rect 171807 254023 171841 254051
rect 171869 254023 171903 254051
rect 171931 254023 171979 254051
rect 171669 253989 171979 254023
rect 171669 253961 171717 253989
rect 171745 253961 171779 253989
rect 171807 253961 171841 253989
rect 171869 253961 171903 253989
rect 171931 253961 171979 253989
rect 171669 245175 171979 253961
rect 171669 245147 171717 245175
rect 171745 245147 171779 245175
rect 171807 245147 171841 245175
rect 171869 245147 171903 245175
rect 171931 245147 171979 245175
rect 171669 245113 171979 245147
rect 171669 245085 171717 245113
rect 171745 245085 171779 245113
rect 171807 245085 171841 245113
rect 171869 245085 171903 245113
rect 171931 245085 171979 245113
rect 171669 245051 171979 245085
rect 171669 245023 171717 245051
rect 171745 245023 171779 245051
rect 171807 245023 171841 245051
rect 171869 245023 171903 245051
rect 171931 245023 171979 245051
rect 171669 244989 171979 245023
rect 171669 244961 171717 244989
rect 171745 244961 171779 244989
rect 171807 244961 171841 244989
rect 171869 244961 171903 244989
rect 171931 244961 171979 244989
rect 171669 236175 171979 244961
rect 171669 236147 171717 236175
rect 171745 236147 171779 236175
rect 171807 236147 171841 236175
rect 171869 236147 171903 236175
rect 171931 236147 171979 236175
rect 171669 236113 171979 236147
rect 171669 236085 171717 236113
rect 171745 236085 171779 236113
rect 171807 236085 171841 236113
rect 171869 236085 171903 236113
rect 171931 236085 171979 236113
rect 171669 236051 171979 236085
rect 171669 236023 171717 236051
rect 171745 236023 171779 236051
rect 171807 236023 171841 236051
rect 171869 236023 171903 236051
rect 171931 236023 171979 236051
rect 171669 235989 171979 236023
rect 171669 235961 171717 235989
rect 171745 235961 171779 235989
rect 171807 235961 171841 235989
rect 171869 235961 171903 235989
rect 171931 235961 171979 235989
rect 171669 227175 171979 235961
rect 171669 227147 171717 227175
rect 171745 227147 171779 227175
rect 171807 227147 171841 227175
rect 171869 227147 171903 227175
rect 171931 227147 171979 227175
rect 171669 227113 171979 227147
rect 171669 227085 171717 227113
rect 171745 227085 171779 227113
rect 171807 227085 171841 227113
rect 171869 227085 171903 227113
rect 171931 227085 171979 227113
rect 171669 227051 171979 227085
rect 171669 227023 171717 227051
rect 171745 227023 171779 227051
rect 171807 227023 171841 227051
rect 171869 227023 171903 227051
rect 171931 227023 171979 227051
rect 171669 226989 171979 227023
rect 171669 226961 171717 226989
rect 171745 226961 171779 226989
rect 171807 226961 171841 226989
rect 171869 226961 171903 226989
rect 171931 226961 171979 226989
rect 171669 218175 171979 226961
rect 171669 218147 171717 218175
rect 171745 218147 171779 218175
rect 171807 218147 171841 218175
rect 171869 218147 171903 218175
rect 171931 218147 171979 218175
rect 171669 218113 171979 218147
rect 171669 218085 171717 218113
rect 171745 218085 171779 218113
rect 171807 218085 171841 218113
rect 171869 218085 171903 218113
rect 171931 218085 171979 218113
rect 171669 218051 171979 218085
rect 171669 218023 171717 218051
rect 171745 218023 171779 218051
rect 171807 218023 171841 218051
rect 171869 218023 171903 218051
rect 171931 218023 171979 218051
rect 171669 217989 171979 218023
rect 171669 217961 171717 217989
rect 171745 217961 171779 217989
rect 171807 217961 171841 217989
rect 171869 217961 171903 217989
rect 171931 217961 171979 217989
rect 171669 209175 171979 217961
rect 171669 209147 171717 209175
rect 171745 209147 171779 209175
rect 171807 209147 171841 209175
rect 171869 209147 171903 209175
rect 171931 209147 171979 209175
rect 171669 209113 171979 209147
rect 171669 209085 171717 209113
rect 171745 209085 171779 209113
rect 171807 209085 171841 209113
rect 171869 209085 171903 209113
rect 171931 209085 171979 209113
rect 171669 209051 171979 209085
rect 171669 209023 171717 209051
rect 171745 209023 171779 209051
rect 171807 209023 171841 209051
rect 171869 209023 171903 209051
rect 171931 209023 171979 209051
rect 171669 208989 171979 209023
rect 171669 208961 171717 208989
rect 171745 208961 171779 208989
rect 171807 208961 171841 208989
rect 171869 208961 171903 208989
rect 171931 208961 171979 208989
rect 171669 200175 171979 208961
rect 171669 200147 171717 200175
rect 171745 200147 171779 200175
rect 171807 200147 171841 200175
rect 171869 200147 171903 200175
rect 171931 200147 171979 200175
rect 171669 200113 171979 200147
rect 171669 200085 171717 200113
rect 171745 200085 171779 200113
rect 171807 200085 171841 200113
rect 171869 200085 171903 200113
rect 171931 200085 171979 200113
rect 171669 200051 171979 200085
rect 171669 200023 171717 200051
rect 171745 200023 171779 200051
rect 171807 200023 171841 200051
rect 171869 200023 171903 200051
rect 171931 200023 171979 200051
rect 171669 199989 171979 200023
rect 171669 199961 171717 199989
rect 171745 199961 171779 199989
rect 171807 199961 171841 199989
rect 171869 199961 171903 199989
rect 171931 199961 171979 199989
rect 171669 191175 171979 199961
rect 171669 191147 171717 191175
rect 171745 191147 171779 191175
rect 171807 191147 171841 191175
rect 171869 191147 171903 191175
rect 171931 191147 171979 191175
rect 171669 191113 171979 191147
rect 171669 191085 171717 191113
rect 171745 191085 171779 191113
rect 171807 191085 171841 191113
rect 171869 191085 171903 191113
rect 171931 191085 171979 191113
rect 171669 191051 171979 191085
rect 171669 191023 171717 191051
rect 171745 191023 171779 191051
rect 171807 191023 171841 191051
rect 171869 191023 171903 191051
rect 171931 191023 171979 191051
rect 171669 190989 171979 191023
rect 171669 190961 171717 190989
rect 171745 190961 171779 190989
rect 171807 190961 171841 190989
rect 171869 190961 171903 190989
rect 171931 190961 171979 190989
rect 171669 182175 171979 190961
rect 171669 182147 171717 182175
rect 171745 182147 171779 182175
rect 171807 182147 171841 182175
rect 171869 182147 171903 182175
rect 171931 182147 171979 182175
rect 171669 182113 171979 182147
rect 171669 182085 171717 182113
rect 171745 182085 171779 182113
rect 171807 182085 171841 182113
rect 171869 182085 171903 182113
rect 171931 182085 171979 182113
rect 171669 182051 171979 182085
rect 171669 182023 171717 182051
rect 171745 182023 171779 182051
rect 171807 182023 171841 182051
rect 171869 182023 171903 182051
rect 171931 182023 171979 182051
rect 171669 181989 171979 182023
rect 171669 181961 171717 181989
rect 171745 181961 171779 181989
rect 171807 181961 171841 181989
rect 171869 181961 171903 181989
rect 171931 181961 171979 181989
rect 161824 173175 161984 173192
rect 161824 173147 161859 173175
rect 161887 173147 161921 173175
rect 161949 173147 161984 173175
rect 161824 173113 161984 173147
rect 161824 173085 161859 173113
rect 161887 173085 161921 173113
rect 161949 173085 161984 173113
rect 161824 173051 161984 173085
rect 161824 173023 161859 173051
rect 161887 173023 161921 173051
rect 161949 173023 161984 173051
rect 161824 172989 161984 173023
rect 161824 172961 161859 172989
rect 161887 172961 161921 172989
rect 161949 172961 161984 172989
rect 161824 172944 161984 172961
rect 171669 173175 171979 181961
rect 171669 173147 171717 173175
rect 171745 173147 171779 173175
rect 171807 173147 171841 173175
rect 171869 173147 171903 173175
rect 171931 173147 171979 173175
rect 171669 173113 171979 173147
rect 171669 173085 171717 173113
rect 171745 173085 171779 173113
rect 171807 173085 171841 173113
rect 171869 173085 171903 173113
rect 171931 173085 171979 173113
rect 171669 173051 171979 173085
rect 171669 173023 171717 173051
rect 171745 173023 171779 173051
rect 171807 173023 171841 173051
rect 171869 173023 171903 173051
rect 171931 173023 171979 173051
rect 171669 172989 171979 173023
rect 171669 172961 171717 172989
rect 171745 172961 171779 172989
rect 171807 172961 171841 172989
rect 171869 172961 171903 172989
rect 171931 172961 171979 172989
rect 158169 167147 158217 167175
rect 158245 167147 158279 167175
rect 158307 167147 158341 167175
rect 158369 167147 158403 167175
rect 158431 167147 158479 167175
rect 158169 167113 158479 167147
rect 158169 167085 158217 167113
rect 158245 167085 158279 167113
rect 158307 167085 158341 167113
rect 158369 167085 158403 167113
rect 158431 167085 158479 167113
rect 158169 167051 158479 167085
rect 158169 167023 158217 167051
rect 158245 167023 158279 167051
rect 158307 167023 158341 167051
rect 158369 167023 158403 167051
rect 158431 167023 158479 167051
rect 158169 166989 158479 167023
rect 158169 166961 158217 166989
rect 158245 166961 158279 166989
rect 158307 166961 158341 166989
rect 158369 166961 158403 166989
rect 158431 166961 158479 166989
rect 158169 158175 158479 166961
rect 169504 167175 169664 167192
rect 169504 167147 169539 167175
rect 169567 167147 169601 167175
rect 169629 167147 169664 167175
rect 169504 167113 169664 167147
rect 169504 167085 169539 167113
rect 169567 167085 169601 167113
rect 169629 167085 169664 167113
rect 169504 167051 169664 167085
rect 169504 167023 169539 167051
rect 169567 167023 169601 167051
rect 169629 167023 169664 167051
rect 169504 166989 169664 167023
rect 169504 166961 169539 166989
rect 169567 166961 169601 166989
rect 169629 166961 169664 166989
rect 169504 166944 169664 166961
rect 161824 164175 161984 164192
rect 161824 164147 161859 164175
rect 161887 164147 161921 164175
rect 161949 164147 161984 164175
rect 161824 164113 161984 164147
rect 161824 164085 161859 164113
rect 161887 164085 161921 164113
rect 161949 164085 161984 164113
rect 161824 164051 161984 164085
rect 161824 164023 161859 164051
rect 161887 164023 161921 164051
rect 161949 164023 161984 164051
rect 161824 163989 161984 164023
rect 161824 163961 161859 163989
rect 161887 163961 161921 163989
rect 161949 163961 161984 163989
rect 161824 163944 161984 163961
rect 171669 164175 171979 172961
rect 171669 164147 171717 164175
rect 171745 164147 171779 164175
rect 171807 164147 171841 164175
rect 171869 164147 171903 164175
rect 171931 164147 171979 164175
rect 171669 164113 171979 164147
rect 171669 164085 171717 164113
rect 171745 164085 171779 164113
rect 171807 164085 171841 164113
rect 171869 164085 171903 164113
rect 171931 164085 171979 164113
rect 171669 164051 171979 164085
rect 171669 164023 171717 164051
rect 171745 164023 171779 164051
rect 171807 164023 171841 164051
rect 171869 164023 171903 164051
rect 171931 164023 171979 164051
rect 171669 163989 171979 164023
rect 171669 163961 171717 163989
rect 171745 163961 171779 163989
rect 171807 163961 171841 163989
rect 171869 163961 171903 163989
rect 171931 163961 171979 163989
rect 158169 158147 158217 158175
rect 158245 158147 158279 158175
rect 158307 158147 158341 158175
rect 158369 158147 158403 158175
rect 158431 158147 158479 158175
rect 158169 158113 158479 158147
rect 158169 158085 158217 158113
rect 158245 158085 158279 158113
rect 158307 158085 158341 158113
rect 158369 158085 158403 158113
rect 158431 158085 158479 158113
rect 158169 158051 158479 158085
rect 158169 158023 158217 158051
rect 158245 158023 158279 158051
rect 158307 158023 158341 158051
rect 158369 158023 158403 158051
rect 158431 158023 158479 158051
rect 158169 157989 158479 158023
rect 158169 157961 158217 157989
rect 158245 157961 158279 157989
rect 158307 157961 158341 157989
rect 158369 157961 158403 157989
rect 158431 157961 158479 157989
rect 158169 149175 158479 157961
rect 169504 158175 169664 158192
rect 169504 158147 169539 158175
rect 169567 158147 169601 158175
rect 169629 158147 169664 158175
rect 169504 158113 169664 158147
rect 169504 158085 169539 158113
rect 169567 158085 169601 158113
rect 169629 158085 169664 158113
rect 169504 158051 169664 158085
rect 169504 158023 169539 158051
rect 169567 158023 169601 158051
rect 169629 158023 169664 158051
rect 169504 157989 169664 158023
rect 169504 157961 169539 157989
rect 169567 157961 169601 157989
rect 169629 157961 169664 157989
rect 169504 157944 169664 157961
rect 161824 155175 161984 155192
rect 161824 155147 161859 155175
rect 161887 155147 161921 155175
rect 161949 155147 161984 155175
rect 161824 155113 161984 155147
rect 161824 155085 161859 155113
rect 161887 155085 161921 155113
rect 161949 155085 161984 155113
rect 161824 155051 161984 155085
rect 161824 155023 161859 155051
rect 161887 155023 161921 155051
rect 161949 155023 161984 155051
rect 161824 154989 161984 155023
rect 161824 154961 161859 154989
rect 161887 154961 161921 154989
rect 161949 154961 161984 154989
rect 161824 154944 161984 154961
rect 171669 155175 171979 163961
rect 171669 155147 171717 155175
rect 171745 155147 171779 155175
rect 171807 155147 171841 155175
rect 171869 155147 171903 155175
rect 171931 155147 171979 155175
rect 171669 155113 171979 155147
rect 171669 155085 171717 155113
rect 171745 155085 171779 155113
rect 171807 155085 171841 155113
rect 171869 155085 171903 155113
rect 171931 155085 171979 155113
rect 171669 155051 171979 155085
rect 171669 155023 171717 155051
rect 171745 155023 171779 155051
rect 171807 155023 171841 155051
rect 171869 155023 171903 155051
rect 171931 155023 171979 155051
rect 171669 154989 171979 155023
rect 171669 154961 171717 154989
rect 171745 154961 171779 154989
rect 171807 154961 171841 154989
rect 171869 154961 171903 154989
rect 171931 154961 171979 154989
rect 158169 149147 158217 149175
rect 158245 149147 158279 149175
rect 158307 149147 158341 149175
rect 158369 149147 158403 149175
rect 158431 149147 158479 149175
rect 158169 149113 158479 149147
rect 158169 149085 158217 149113
rect 158245 149085 158279 149113
rect 158307 149085 158341 149113
rect 158369 149085 158403 149113
rect 158431 149085 158479 149113
rect 158169 149051 158479 149085
rect 158169 149023 158217 149051
rect 158245 149023 158279 149051
rect 158307 149023 158341 149051
rect 158369 149023 158403 149051
rect 158431 149023 158479 149051
rect 158169 148989 158479 149023
rect 158169 148961 158217 148989
rect 158245 148961 158279 148989
rect 158307 148961 158341 148989
rect 158369 148961 158403 148989
rect 158431 148961 158479 148989
rect 158169 140175 158479 148961
rect 169504 149175 169664 149192
rect 169504 149147 169539 149175
rect 169567 149147 169601 149175
rect 169629 149147 169664 149175
rect 169504 149113 169664 149147
rect 169504 149085 169539 149113
rect 169567 149085 169601 149113
rect 169629 149085 169664 149113
rect 169504 149051 169664 149085
rect 169504 149023 169539 149051
rect 169567 149023 169601 149051
rect 169629 149023 169664 149051
rect 169504 148989 169664 149023
rect 169504 148961 169539 148989
rect 169567 148961 169601 148989
rect 169629 148961 169664 148989
rect 169504 148944 169664 148961
rect 161824 146175 161984 146192
rect 161824 146147 161859 146175
rect 161887 146147 161921 146175
rect 161949 146147 161984 146175
rect 161824 146113 161984 146147
rect 161824 146085 161859 146113
rect 161887 146085 161921 146113
rect 161949 146085 161984 146113
rect 161824 146051 161984 146085
rect 161824 146023 161859 146051
rect 161887 146023 161921 146051
rect 161949 146023 161984 146051
rect 161824 145989 161984 146023
rect 161824 145961 161859 145989
rect 161887 145961 161921 145989
rect 161949 145961 161984 145989
rect 161824 145944 161984 145961
rect 171669 146175 171979 154961
rect 171669 146147 171717 146175
rect 171745 146147 171779 146175
rect 171807 146147 171841 146175
rect 171869 146147 171903 146175
rect 171931 146147 171979 146175
rect 171669 146113 171979 146147
rect 171669 146085 171717 146113
rect 171745 146085 171779 146113
rect 171807 146085 171841 146113
rect 171869 146085 171903 146113
rect 171931 146085 171979 146113
rect 171669 146051 171979 146085
rect 171669 146023 171717 146051
rect 171745 146023 171779 146051
rect 171807 146023 171841 146051
rect 171869 146023 171903 146051
rect 171931 146023 171979 146051
rect 171669 145989 171979 146023
rect 171669 145961 171717 145989
rect 171745 145961 171779 145989
rect 171807 145961 171841 145989
rect 171869 145961 171903 145989
rect 171931 145961 171979 145989
rect 158169 140147 158217 140175
rect 158245 140147 158279 140175
rect 158307 140147 158341 140175
rect 158369 140147 158403 140175
rect 158431 140147 158479 140175
rect 158169 140113 158479 140147
rect 158169 140085 158217 140113
rect 158245 140085 158279 140113
rect 158307 140085 158341 140113
rect 158369 140085 158403 140113
rect 158431 140085 158479 140113
rect 158169 140051 158479 140085
rect 158169 140023 158217 140051
rect 158245 140023 158279 140051
rect 158307 140023 158341 140051
rect 158369 140023 158403 140051
rect 158431 140023 158479 140051
rect 158169 139989 158479 140023
rect 158169 139961 158217 139989
rect 158245 139961 158279 139989
rect 158307 139961 158341 139989
rect 158369 139961 158403 139989
rect 158431 139961 158479 139989
rect 158169 131175 158479 139961
rect 169504 140175 169664 140192
rect 169504 140147 169539 140175
rect 169567 140147 169601 140175
rect 169629 140147 169664 140175
rect 169504 140113 169664 140147
rect 169504 140085 169539 140113
rect 169567 140085 169601 140113
rect 169629 140085 169664 140113
rect 169504 140051 169664 140085
rect 169504 140023 169539 140051
rect 169567 140023 169601 140051
rect 169629 140023 169664 140051
rect 169504 139989 169664 140023
rect 169504 139961 169539 139989
rect 169567 139961 169601 139989
rect 169629 139961 169664 139989
rect 169504 139944 169664 139961
rect 161824 137175 161984 137192
rect 161824 137147 161859 137175
rect 161887 137147 161921 137175
rect 161949 137147 161984 137175
rect 161824 137113 161984 137147
rect 161824 137085 161859 137113
rect 161887 137085 161921 137113
rect 161949 137085 161984 137113
rect 161824 137051 161984 137085
rect 161824 137023 161859 137051
rect 161887 137023 161921 137051
rect 161949 137023 161984 137051
rect 161824 136989 161984 137023
rect 161824 136961 161859 136989
rect 161887 136961 161921 136989
rect 161949 136961 161984 136989
rect 161824 136944 161984 136961
rect 171669 137175 171979 145961
rect 171669 137147 171717 137175
rect 171745 137147 171779 137175
rect 171807 137147 171841 137175
rect 171869 137147 171903 137175
rect 171931 137147 171979 137175
rect 171669 137113 171979 137147
rect 171669 137085 171717 137113
rect 171745 137085 171779 137113
rect 171807 137085 171841 137113
rect 171869 137085 171903 137113
rect 171931 137085 171979 137113
rect 171669 137051 171979 137085
rect 171669 137023 171717 137051
rect 171745 137023 171779 137051
rect 171807 137023 171841 137051
rect 171869 137023 171903 137051
rect 171931 137023 171979 137051
rect 171669 136989 171979 137023
rect 171669 136961 171717 136989
rect 171745 136961 171779 136989
rect 171807 136961 171841 136989
rect 171869 136961 171903 136989
rect 171931 136961 171979 136989
rect 158169 131147 158217 131175
rect 158245 131147 158279 131175
rect 158307 131147 158341 131175
rect 158369 131147 158403 131175
rect 158431 131147 158479 131175
rect 158169 131113 158479 131147
rect 158169 131085 158217 131113
rect 158245 131085 158279 131113
rect 158307 131085 158341 131113
rect 158369 131085 158403 131113
rect 158431 131085 158479 131113
rect 158169 131051 158479 131085
rect 158169 131023 158217 131051
rect 158245 131023 158279 131051
rect 158307 131023 158341 131051
rect 158369 131023 158403 131051
rect 158431 131023 158479 131051
rect 158169 130989 158479 131023
rect 158169 130961 158217 130989
rect 158245 130961 158279 130989
rect 158307 130961 158341 130989
rect 158369 130961 158403 130989
rect 158431 130961 158479 130989
rect 158169 122175 158479 130961
rect 169504 131175 169664 131192
rect 169504 131147 169539 131175
rect 169567 131147 169601 131175
rect 169629 131147 169664 131175
rect 169504 131113 169664 131147
rect 169504 131085 169539 131113
rect 169567 131085 169601 131113
rect 169629 131085 169664 131113
rect 169504 131051 169664 131085
rect 169504 131023 169539 131051
rect 169567 131023 169601 131051
rect 169629 131023 169664 131051
rect 169504 130989 169664 131023
rect 169504 130961 169539 130989
rect 169567 130961 169601 130989
rect 169629 130961 169664 130989
rect 169504 130944 169664 130961
rect 161824 128175 161984 128192
rect 161824 128147 161859 128175
rect 161887 128147 161921 128175
rect 161949 128147 161984 128175
rect 161824 128113 161984 128147
rect 161824 128085 161859 128113
rect 161887 128085 161921 128113
rect 161949 128085 161984 128113
rect 161824 128051 161984 128085
rect 161824 128023 161859 128051
rect 161887 128023 161921 128051
rect 161949 128023 161984 128051
rect 161824 127989 161984 128023
rect 161824 127961 161859 127989
rect 161887 127961 161921 127989
rect 161949 127961 161984 127989
rect 161824 127944 161984 127961
rect 171669 128175 171979 136961
rect 171669 128147 171717 128175
rect 171745 128147 171779 128175
rect 171807 128147 171841 128175
rect 171869 128147 171903 128175
rect 171931 128147 171979 128175
rect 171669 128113 171979 128147
rect 171669 128085 171717 128113
rect 171745 128085 171779 128113
rect 171807 128085 171841 128113
rect 171869 128085 171903 128113
rect 171931 128085 171979 128113
rect 171669 128051 171979 128085
rect 171669 128023 171717 128051
rect 171745 128023 171779 128051
rect 171807 128023 171841 128051
rect 171869 128023 171903 128051
rect 171931 128023 171979 128051
rect 171669 127989 171979 128023
rect 171669 127961 171717 127989
rect 171745 127961 171779 127989
rect 171807 127961 171841 127989
rect 171869 127961 171903 127989
rect 171931 127961 171979 127989
rect 158169 122147 158217 122175
rect 158245 122147 158279 122175
rect 158307 122147 158341 122175
rect 158369 122147 158403 122175
rect 158431 122147 158479 122175
rect 158169 122113 158479 122147
rect 158169 122085 158217 122113
rect 158245 122085 158279 122113
rect 158307 122085 158341 122113
rect 158369 122085 158403 122113
rect 158431 122085 158479 122113
rect 158169 122051 158479 122085
rect 158169 122023 158217 122051
rect 158245 122023 158279 122051
rect 158307 122023 158341 122051
rect 158369 122023 158403 122051
rect 158431 122023 158479 122051
rect 158169 121989 158479 122023
rect 158169 121961 158217 121989
rect 158245 121961 158279 121989
rect 158307 121961 158341 121989
rect 158369 121961 158403 121989
rect 158431 121961 158479 121989
rect 158169 113175 158479 121961
rect 169504 122175 169664 122192
rect 169504 122147 169539 122175
rect 169567 122147 169601 122175
rect 169629 122147 169664 122175
rect 169504 122113 169664 122147
rect 169504 122085 169539 122113
rect 169567 122085 169601 122113
rect 169629 122085 169664 122113
rect 169504 122051 169664 122085
rect 169504 122023 169539 122051
rect 169567 122023 169601 122051
rect 169629 122023 169664 122051
rect 169504 121989 169664 122023
rect 169504 121961 169539 121989
rect 169567 121961 169601 121989
rect 169629 121961 169664 121989
rect 169504 121944 169664 121961
rect 161824 119175 161984 119192
rect 161824 119147 161859 119175
rect 161887 119147 161921 119175
rect 161949 119147 161984 119175
rect 161824 119113 161984 119147
rect 161824 119085 161859 119113
rect 161887 119085 161921 119113
rect 161949 119085 161984 119113
rect 161824 119051 161984 119085
rect 161824 119023 161859 119051
rect 161887 119023 161921 119051
rect 161949 119023 161984 119051
rect 161824 118989 161984 119023
rect 161824 118961 161859 118989
rect 161887 118961 161921 118989
rect 161949 118961 161984 118989
rect 161824 118944 161984 118961
rect 171669 119175 171979 127961
rect 171669 119147 171717 119175
rect 171745 119147 171779 119175
rect 171807 119147 171841 119175
rect 171869 119147 171903 119175
rect 171931 119147 171979 119175
rect 171669 119113 171979 119147
rect 171669 119085 171717 119113
rect 171745 119085 171779 119113
rect 171807 119085 171841 119113
rect 171869 119085 171903 119113
rect 171931 119085 171979 119113
rect 171669 119051 171979 119085
rect 171669 119023 171717 119051
rect 171745 119023 171779 119051
rect 171807 119023 171841 119051
rect 171869 119023 171903 119051
rect 171931 119023 171979 119051
rect 171669 118989 171979 119023
rect 171669 118961 171717 118989
rect 171745 118961 171779 118989
rect 171807 118961 171841 118989
rect 171869 118961 171903 118989
rect 171931 118961 171979 118989
rect 158169 113147 158217 113175
rect 158245 113147 158279 113175
rect 158307 113147 158341 113175
rect 158369 113147 158403 113175
rect 158431 113147 158479 113175
rect 158169 113113 158479 113147
rect 158169 113085 158217 113113
rect 158245 113085 158279 113113
rect 158307 113085 158341 113113
rect 158369 113085 158403 113113
rect 158431 113085 158479 113113
rect 158169 113051 158479 113085
rect 158169 113023 158217 113051
rect 158245 113023 158279 113051
rect 158307 113023 158341 113051
rect 158369 113023 158403 113051
rect 158431 113023 158479 113051
rect 158169 112989 158479 113023
rect 158169 112961 158217 112989
rect 158245 112961 158279 112989
rect 158307 112961 158341 112989
rect 158369 112961 158403 112989
rect 158431 112961 158479 112989
rect 158169 104175 158479 112961
rect 169504 113175 169664 113192
rect 169504 113147 169539 113175
rect 169567 113147 169601 113175
rect 169629 113147 169664 113175
rect 169504 113113 169664 113147
rect 169504 113085 169539 113113
rect 169567 113085 169601 113113
rect 169629 113085 169664 113113
rect 169504 113051 169664 113085
rect 169504 113023 169539 113051
rect 169567 113023 169601 113051
rect 169629 113023 169664 113051
rect 169504 112989 169664 113023
rect 169504 112961 169539 112989
rect 169567 112961 169601 112989
rect 169629 112961 169664 112989
rect 169504 112944 169664 112961
rect 161824 110175 161984 110192
rect 161824 110147 161859 110175
rect 161887 110147 161921 110175
rect 161949 110147 161984 110175
rect 161824 110113 161984 110147
rect 161824 110085 161859 110113
rect 161887 110085 161921 110113
rect 161949 110085 161984 110113
rect 161824 110051 161984 110085
rect 161824 110023 161859 110051
rect 161887 110023 161921 110051
rect 161949 110023 161984 110051
rect 161824 109989 161984 110023
rect 161824 109961 161859 109989
rect 161887 109961 161921 109989
rect 161949 109961 161984 109989
rect 161824 109944 161984 109961
rect 171669 110175 171979 118961
rect 171669 110147 171717 110175
rect 171745 110147 171779 110175
rect 171807 110147 171841 110175
rect 171869 110147 171903 110175
rect 171931 110147 171979 110175
rect 171669 110113 171979 110147
rect 171669 110085 171717 110113
rect 171745 110085 171779 110113
rect 171807 110085 171841 110113
rect 171869 110085 171903 110113
rect 171931 110085 171979 110113
rect 171669 110051 171979 110085
rect 171669 110023 171717 110051
rect 171745 110023 171779 110051
rect 171807 110023 171841 110051
rect 171869 110023 171903 110051
rect 171931 110023 171979 110051
rect 171669 109989 171979 110023
rect 171669 109961 171717 109989
rect 171745 109961 171779 109989
rect 171807 109961 171841 109989
rect 171869 109961 171903 109989
rect 171931 109961 171979 109989
rect 158169 104147 158217 104175
rect 158245 104147 158279 104175
rect 158307 104147 158341 104175
rect 158369 104147 158403 104175
rect 158431 104147 158479 104175
rect 158169 104113 158479 104147
rect 158169 104085 158217 104113
rect 158245 104085 158279 104113
rect 158307 104085 158341 104113
rect 158369 104085 158403 104113
rect 158431 104085 158479 104113
rect 158169 104051 158479 104085
rect 158169 104023 158217 104051
rect 158245 104023 158279 104051
rect 158307 104023 158341 104051
rect 158369 104023 158403 104051
rect 158431 104023 158479 104051
rect 158169 103989 158479 104023
rect 158169 103961 158217 103989
rect 158245 103961 158279 103989
rect 158307 103961 158341 103989
rect 158369 103961 158403 103989
rect 158431 103961 158479 103989
rect 158169 95175 158479 103961
rect 169504 104175 169664 104192
rect 169504 104147 169539 104175
rect 169567 104147 169601 104175
rect 169629 104147 169664 104175
rect 169504 104113 169664 104147
rect 169504 104085 169539 104113
rect 169567 104085 169601 104113
rect 169629 104085 169664 104113
rect 169504 104051 169664 104085
rect 169504 104023 169539 104051
rect 169567 104023 169601 104051
rect 169629 104023 169664 104051
rect 169504 103989 169664 104023
rect 169504 103961 169539 103989
rect 169567 103961 169601 103989
rect 169629 103961 169664 103989
rect 169504 103944 169664 103961
rect 161824 101175 161984 101192
rect 161824 101147 161859 101175
rect 161887 101147 161921 101175
rect 161949 101147 161984 101175
rect 161824 101113 161984 101147
rect 161824 101085 161859 101113
rect 161887 101085 161921 101113
rect 161949 101085 161984 101113
rect 161824 101051 161984 101085
rect 161824 101023 161859 101051
rect 161887 101023 161921 101051
rect 161949 101023 161984 101051
rect 161824 100989 161984 101023
rect 161824 100961 161859 100989
rect 161887 100961 161921 100989
rect 161949 100961 161984 100989
rect 161824 100944 161984 100961
rect 171669 101175 171979 109961
rect 171669 101147 171717 101175
rect 171745 101147 171779 101175
rect 171807 101147 171841 101175
rect 171869 101147 171903 101175
rect 171931 101147 171979 101175
rect 171669 101113 171979 101147
rect 171669 101085 171717 101113
rect 171745 101085 171779 101113
rect 171807 101085 171841 101113
rect 171869 101085 171903 101113
rect 171931 101085 171979 101113
rect 171669 101051 171979 101085
rect 171669 101023 171717 101051
rect 171745 101023 171779 101051
rect 171807 101023 171841 101051
rect 171869 101023 171903 101051
rect 171931 101023 171979 101051
rect 171669 100989 171979 101023
rect 171669 100961 171717 100989
rect 171745 100961 171779 100989
rect 171807 100961 171841 100989
rect 171869 100961 171903 100989
rect 171931 100961 171979 100989
rect 158169 95147 158217 95175
rect 158245 95147 158279 95175
rect 158307 95147 158341 95175
rect 158369 95147 158403 95175
rect 158431 95147 158479 95175
rect 158169 95113 158479 95147
rect 158169 95085 158217 95113
rect 158245 95085 158279 95113
rect 158307 95085 158341 95113
rect 158369 95085 158403 95113
rect 158431 95085 158479 95113
rect 158169 95051 158479 95085
rect 158169 95023 158217 95051
rect 158245 95023 158279 95051
rect 158307 95023 158341 95051
rect 158369 95023 158403 95051
rect 158431 95023 158479 95051
rect 158169 94989 158479 95023
rect 158169 94961 158217 94989
rect 158245 94961 158279 94989
rect 158307 94961 158341 94989
rect 158369 94961 158403 94989
rect 158431 94961 158479 94989
rect 158169 86175 158479 94961
rect 169504 95175 169664 95192
rect 169504 95147 169539 95175
rect 169567 95147 169601 95175
rect 169629 95147 169664 95175
rect 169504 95113 169664 95147
rect 169504 95085 169539 95113
rect 169567 95085 169601 95113
rect 169629 95085 169664 95113
rect 169504 95051 169664 95085
rect 169504 95023 169539 95051
rect 169567 95023 169601 95051
rect 169629 95023 169664 95051
rect 169504 94989 169664 95023
rect 169504 94961 169539 94989
rect 169567 94961 169601 94989
rect 169629 94961 169664 94989
rect 169504 94944 169664 94961
rect 161824 92175 161984 92192
rect 161824 92147 161859 92175
rect 161887 92147 161921 92175
rect 161949 92147 161984 92175
rect 161824 92113 161984 92147
rect 161824 92085 161859 92113
rect 161887 92085 161921 92113
rect 161949 92085 161984 92113
rect 161824 92051 161984 92085
rect 161824 92023 161859 92051
rect 161887 92023 161921 92051
rect 161949 92023 161984 92051
rect 161824 91989 161984 92023
rect 161824 91961 161859 91989
rect 161887 91961 161921 91989
rect 161949 91961 161984 91989
rect 161824 91944 161984 91961
rect 171669 92175 171979 100961
rect 171669 92147 171717 92175
rect 171745 92147 171779 92175
rect 171807 92147 171841 92175
rect 171869 92147 171903 92175
rect 171931 92147 171979 92175
rect 171669 92113 171979 92147
rect 171669 92085 171717 92113
rect 171745 92085 171779 92113
rect 171807 92085 171841 92113
rect 171869 92085 171903 92113
rect 171931 92085 171979 92113
rect 171669 92051 171979 92085
rect 171669 92023 171717 92051
rect 171745 92023 171779 92051
rect 171807 92023 171841 92051
rect 171869 92023 171903 92051
rect 171931 92023 171979 92051
rect 171669 91989 171979 92023
rect 171669 91961 171717 91989
rect 171745 91961 171779 91989
rect 171807 91961 171841 91989
rect 171869 91961 171903 91989
rect 171931 91961 171979 91989
rect 158169 86147 158217 86175
rect 158245 86147 158279 86175
rect 158307 86147 158341 86175
rect 158369 86147 158403 86175
rect 158431 86147 158479 86175
rect 158169 86113 158479 86147
rect 158169 86085 158217 86113
rect 158245 86085 158279 86113
rect 158307 86085 158341 86113
rect 158369 86085 158403 86113
rect 158431 86085 158479 86113
rect 158169 86051 158479 86085
rect 158169 86023 158217 86051
rect 158245 86023 158279 86051
rect 158307 86023 158341 86051
rect 158369 86023 158403 86051
rect 158431 86023 158479 86051
rect 158169 85989 158479 86023
rect 158169 85961 158217 85989
rect 158245 85961 158279 85989
rect 158307 85961 158341 85989
rect 158369 85961 158403 85989
rect 158431 85961 158479 85989
rect 158169 77175 158479 85961
rect 169504 86175 169664 86192
rect 169504 86147 169539 86175
rect 169567 86147 169601 86175
rect 169629 86147 169664 86175
rect 169504 86113 169664 86147
rect 169504 86085 169539 86113
rect 169567 86085 169601 86113
rect 169629 86085 169664 86113
rect 169504 86051 169664 86085
rect 169504 86023 169539 86051
rect 169567 86023 169601 86051
rect 169629 86023 169664 86051
rect 169504 85989 169664 86023
rect 169504 85961 169539 85989
rect 169567 85961 169601 85989
rect 169629 85961 169664 85989
rect 169504 85944 169664 85961
rect 161824 83175 161984 83192
rect 161824 83147 161859 83175
rect 161887 83147 161921 83175
rect 161949 83147 161984 83175
rect 161824 83113 161984 83147
rect 161824 83085 161859 83113
rect 161887 83085 161921 83113
rect 161949 83085 161984 83113
rect 161824 83051 161984 83085
rect 161824 83023 161859 83051
rect 161887 83023 161921 83051
rect 161949 83023 161984 83051
rect 161824 82989 161984 83023
rect 161824 82961 161859 82989
rect 161887 82961 161921 82989
rect 161949 82961 161984 82989
rect 161824 82944 161984 82961
rect 171669 83175 171979 91961
rect 171669 83147 171717 83175
rect 171745 83147 171779 83175
rect 171807 83147 171841 83175
rect 171869 83147 171903 83175
rect 171931 83147 171979 83175
rect 171669 83113 171979 83147
rect 171669 83085 171717 83113
rect 171745 83085 171779 83113
rect 171807 83085 171841 83113
rect 171869 83085 171903 83113
rect 171931 83085 171979 83113
rect 171669 83051 171979 83085
rect 171669 83023 171717 83051
rect 171745 83023 171779 83051
rect 171807 83023 171841 83051
rect 171869 83023 171903 83051
rect 171931 83023 171979 83051
rect 171669 82989 171979 83023
rect 171669 82961 171717 82989
rect 171745 82961 171779 82989
rect 171807 82961 171841 82989
rect 171869 82961 171903 82989
rect 171931 82961 171979 82989
rect 158169 77147 158217 77175
rect 158245 77147 158279 77175
rect 158307 77147 158341 77175
rect 158369 77147 158403 77175
rect 158431 77147 158479 77175
rect 158169 77113 158479 77147
rect 158169 77085 158217 77113
rect 158245 77085 158279 77113
rect 158307 77085 158341 77113
rect 158369 77085 158403 77113
rect 158431 77085 158479 77113
rect 158169 77051 158479 77085
rect 158169 77023 158217 77051
rect 158245 77023 158279 77051
rect 158307 77023 158341 77051
rect 158369 77023 158403 77051
rect 158431 77023 158479 77051
rect 158169 76989 158479 77023
rect 158169 76961 158217 76989
rect 158245 76961 158279 76989
rect 158307 76961 158341 76989
rect 158369 76961 158403 76989
rect 158431 76961 158479 76989
rect 158169 68175 158479 76961
rect 169504 77175 169664 77192
rect 169504 77147 169539 77175
rect 169567 77147 169601 77175
rect 169629 77147 169664 77175
rect 169504 77113 169664 77147
rect 169504 77085 169539 77113
rect 169567 77085 169601 77113
rect 169629 77085 169664 77113
rect 169504 77051 169664 77085
rect 169504 77023 169539 77051
rect 169567 77023 169601 77051
rect 169629 77023 169664 77051
rect 169504 76989 169664 77023
rect 169504 76961 169539 76989
rect 169567 76961 169601 76989
rect 169629 76961 169664 76989
rect 169504 76944 169664 76961
rect 161824 74175 161984 74192
rect 161824 74147 161859 74175
rect 161887 74147 161921 74175
rect 161949 74147 161984 74175
rect 161824 74113 161984 74147
rect 161824 74085 161859 74113
rect 161887 74085 161921 74113
rect 161949 74085 161984 74113
rect 161824 74051 161984 74085
rect 161824 74023 161859 74051
rect 161887 74023 161921 74051
rect 161949 74023 161984 74051
rect 161824 73989 161984 74023
rect 161824 73961 161859 73989
rect 161887 73961 161921 73989
rect 161949 73961 161984 73989
rect 161824 73944 161984 73961
rect 171669 74175 171979 82961
rect 171669 74147 171717 74175
rect 171745 74147 171779 74175
rect 171807 74147 171841 74175
rect 171869 74147 171903 74175
rect 171931 74147 171979 74175
rect 171669 74113 171979 74147
rect 171669 74085 171717 74113
rect 171745 74085 171779 74113
rect 171807 74085 171841 74113
rect 171869 74085 171903 74113
rect 171931 74085 171979 74113
rect 171669 74051 171979 74085
rect 171669 74023 171717 74051
rect 171745 74023 171779 74051
rect 171807 74023 171841 74051
rect 171869 74023 171903 74051
rect 171931 74023 171979 74051
rect 171669 73989 171979 74023
rect 171669 73961 171717 73989
rect 171745 73961 171779 73989
rect 171807 73961 171841 73989
rect 171869 73961 171903 73989
rect 171931 73961 171979 73989
rect 158169 68147 158217 68175
rect 158245 68147 158279 68175
rect 158307 68147 158341 68175
rect 158369 68147 158403 68175
rect 158431 68147 158479 68175
rect 158169 68113 158479 68147
rect 158169 68085 158217 68113
rect 158245 68085 158279 68113
rect 158307 68085 158341 68113
rect 158369 68085 158403 68113
rect 158431 68085 158479 68113
rect 158169 68051 158479 68085
rect 158169 68023 158217 68051
rect 158245 68023 158279 68051
rect 158307 68023 158341 68051
rect 158369 68023 158403 68051
rect 158431 68023 158479 68051
rect 158169 67989 158479 68023
rect 158169 67961 158217 67989
rect 158245 67961 158279 67989
rect 158307 67961 158341 67989
rect 158369 67961 158403 67989
rect 158431 67961 158479 67989
rect 158169 59175 158479 67961
rect 169504 68175 169664 68192
rect 169504 68147 169539 68175
rect 169567 68147 169601 68175
rect 169629 68147 169664 68175
rect 169504 68113 169664 68147
rect 169504 68085 169539 68113
rect 169567 68085 169601 68113
rect 169629 68085 169664 68113
rect 169504 68051 169664 68085
rect 169504 68023 169539 68051
rect 169567 68023 169601 68051
rect 169629 68023 169664 68051
rect 169504 67989 169664 68023
rect 169504 67961 169539 67989
rect 169567 67961 169601 67989
rect 169629 67961 169664 67989
rect 169504 67944 169664 67961
rect 161824 65175 161984 65192
rect 161824 65147 161859 65175
rect 161887 65147 161921 65175
rect 161949 65147 161984 65175
rect 161824 65113 161984 65147
rect 161824 65085 161859 65113
rect 161887 65085 161921 65113
rect 161949 65085 161984 65113
rect 161824 65051 161984 65085
rect 161824 65023 161859 65051
rect 161887 65023 161921 65051
rect 161949 65023 161984 65051
rect 161824 64989 161984 65023
rect 161824 64961 161859 64989
rect 161887 64961 161921 64989
rect 161949 64961 161984 64989
rect 161824 64944 161984 64961
rect 171669 65175 171979 73961
rect 171669 65147 171717 65175
rect 171745 65147 171779 65175
rect 171807 65147 171841 65175
rect 171869 65147 171903 65175
rect 171931 65147 171979 65175
rect 171669 65113 171979 65147
rect 171669 65085 171717 65113
rect 171745 65085 171779 65113
rect 171807 65085 171841 65113
rect 171869 65085 171903 65113
rect 171931 65085 171979 65113
rect 171669 65051 171979 65085
rect 171669 65023 171717 65051
rect 171745 65023 171779 65051
rect 171807 65023 171841 65051
rect 171869 65023 171903 65051
rect 171931 65023 171979 65051
rect 171669 64989 171979 65023
rect 171669 64961 171717 64989
rect 171745 64961 171779 64989
rect 171807 64961 171841 64989
rect 171869 64961 171903 64989
rect 171931 64961 171979 64989
rect 158169 59147 158217 59175
rect 158245 59147 158279 59175
rect 158307 59147 158341 59175
rect 158369 59147 158403 59175
rect 158431 59147 158479 59175
rect 158169 59113 158479 59147
rect 158169 59085 158217 59113
rect 158245 59085 158279 59113
rect 158307 59085 158341 59113
rect 158369 59085 158403 59113
rect 158431 59085 158479 59113
rect 158169 59051 158479 59085
rect 158169 59023 158217 59051
rect 158245 59023 158279 59051
rect 158307 59023 158341 59051
rect 158369 59023 158403 59051
rect 158431 59023 158479 59051
rect 158169 58989 158479 59023
rect 158169 58961 158217 58989
rect 158245 58961 158279 58989
rect 158307 58961 158341 58989
rect 158369 58961 158403 58989
rect 158431 58961 158479 58989
rect 158169 50175 158479 58961
rect 169504 59175 169664 59192
rect 169504 59147 169539 59175
rect 169567 59147 169601 59175
rect 169629 59147 169664 59175
rect 169504 59113 169664 59147
rect 169504 59085 169539 59113
rect 169567 59085 169601 59113
rect 169629 59085 169664 59113
rect 169504 59051 169664 59085
rect 169504 59023 169539 59051
rect 169567 59023 169601 59051
rect 169629 59023 169664 59051
rect 169504 58989 169664 59023
rect 169504 58961 169539 58989
rect 169567 58961 169601 58989
rect 169629 58961 169664 58989
rect 169504 58944 169664 58961
rect 161824 56175 161984 56192
rect 161824 56147 161859 56175
rect 161887 56147 161921 56175
rect 161949 56147 161984 56175
rect 161824 56113 161984 56147
rect 161824 56085 161859 56113
rect 161887 56085 161921 56113
rect 161949 56085 161984 56113
rect 161824 56051 161984 56085
rect 161824 56023 161859 56051
rect 161887 56023 161921 56051
rect 161949 56023 161984 56051
rect 161824 55989 161984 56023
rect 161824 55961 161859 55989
rect 161887 55961 161921 55989
rect 161949 55961 161984 55989
rect 161824 55944 161984 55961
rect 171669 56175 171979 64961
rect 171669 56147 171717 56175
rect 171745 56147 171779 56175
rect 171807 56147 171841 56175
rect 171869 56147 171903 56175
rect 171931 56147 171979 56175
rect 171669 56113 171979 56147
rect 171669 56085 171717 56113
rect 171745 56085 171779 56113
rect 171807 56085 171841 56113
rect 171869 56085 171903 56113
rect 171931 56085 171979 56113
rect 171669 56051 171979 56085
rect 171669 56023 171717 56051
rect 171745 56023 171779 56051
rect 171807 56023 171841 56051
rect 171869 56023 171903 56051
rect 171931 56023 171979 56051
rect 171669 55989 171979 56023
rect 171669 55961 171717 55989
rect 171745 55961 171779 55989
rect 171807 55961 171841 55989
rect 171869 55961 171903 55989
rect 171931 55961 171979 55989
rect 158169 50147 158217 50175
rect 158245 50147 158279 50175
rect 158307 50147 158341 50175
rect 158369 50147 158403 50175
rect 158431 50147 158479 50175
rect 158169 50113 158479 50147
rect 158169 50085 158217 50113
rect 158245 50085 158279 50113
rect 158307 50085 158341 50113
rect 158369 50085 158403 50113
rect 158431 50085 158479 50113
rect 158169 50051 158479 50085
rect 158169 50023 158217 50051
rect 158245 50023 158279 50051
rect 158307 50023 158341 50051
rect 158369 50023 158403 50051
rect 158431 50023 158479 50051
rect 158169 49989 158479 50023
rect 158169 49961 158217 49989
rect 158245 49961 158279 49989
rect 158307 49961 158341 49989
rect 158369 49961 158403 49989
rect 158431 49961 158479 49989
rect 158169 41175 158479 49961
rect 169504 50175 169664 50192
rect 169504 50147 169539 50175
rect 169567 50147 169601 50175
rect 169629 50147 169664 50175
rect 169504 50113 169664 50147
rect 169504 50085 169539 50113
rect 169567 50085 169601 50113
rect 169629 50085 169664 50113
rect 169504 50051 169664 50085
rect 169504 50023 169539 50051
rect 169567 50023 169601 50051
rect 169629 50023 169664 50051
rect 169504 49989 169664 50023
rect 169504 49961 169539 49989
rect 169567 49961 169601 49989
rect 169629 49961 169664 49989
rect 169504 49944 169664 49961
rect 161824 47175 161984 47192
rect 161824 47147 161859 47175
rect 161887 47147 161921 47175
rect 161949 47147 161984 47175
rect 161824 47113 161984 47147
rect 161824 47085 161859 47113
rect 161887 47085 161921 47113
rect 161949 47085 161984 47113
rect 161824 47051 161984 47085
rect 161824 47023 161859 47051
rect 161887 47023 161921 47051
rect 161949 47023 161984 47051
rect 161824 46989 161984 47023
rect 161824 46961 161859 46989
rect 161887 46961 161921 46989
rect 161949 46961 161984 46989
rect 161824 46944 161984 46961
rect 171669 47175 171979 55961
rect 171669 47147 171717 47175
rect 171745 47147 171779 47175
rect 171807 47147 171841 47175
rect 171869 47147 171903 47175
rect 171931 47147 171979 47175
rect 171669 47113 171979 47147
rect 171669 47085 171717 47113
rect 171745 47085 171779 47113
rect 171807 47085 171841 47113
rect 171869 47085 171903 47113
rect 171931 47085 171979 47113
rect 171669 47051 171979 47085
rect 171669 47023 171717 47051
rect 171745 47023 171779 47051
rect 171807 47023 171841 47051
rect 171869 47023 171903 47051
rect 171931 47023 171979 47051
rect 171669 46989 171979 47023
rect 171669 46961 171717 46989
rect 171745 46961 171779 46989
rect 171807 46961 171841 46989
rect 171869 46961 171903 46989
rect 171931 46961 171979 46989
rect 158169 41147 158217 41175
rect 158245 41147 158279 41175
rect 158307 41147 158341 41175
rect 158369 41147 158403 41175
rect 158431 41147 158479 41175
rect 158169 41113 158479 41147
rect 158169 41085 158217 41113
rect 158245 41085 158279 41113
rect 158307 41085 158341 41113
rect 158369 41085 158403 41113
rect 158431 41085 158479 41113
rect 158169 41051 158479 41085
rect 158169 41023 158217 41051
rect 158245 41023 158279 41051
rect 158307 41023 158341 41051
rect 158369 41023 158403 41051
rect 158431 41023 158479 41051
rect 158169 40989 158479 41023
rect 158169 40961 158217 40989
rect 158245 40961 158279 40989
rect 158307 40961 158341 40989
rect 158369 40961 158403 40989
rect 158431 40961 158479 40989
rect 158169 32175 158479 40961
rect 169504 41175 169664 41192
rect 169504 41147 169539 41175
rect 169567 41147 169601 41175
rect 169629 41147 169664 41175
rect 169504 41113 169664 41147
rect 169504 41085 169539 41113
rect 169567 41085 169601 41113
rect 169629 41085 169664 41113
rect 169504 41051 169664 41085
rect 169504 41023 169539 41051
rect 169567 41023 169601 41051
rect 169629 41023 169664 41051
rect 169504 40989 169664 41023
rect 169504 40961 169539 40989
rect 169567 40961 169601 40989
rect 169629 40961 169664 40989
rect 169504 40944 169664 40961
rect 161824 38175 161984 38192
rect 161824 38147 161859 38175
rect 161887 38147 161921 38175
rect 161949 38147 161984 38175
rect 161824 38113 161984 38147
rect 161824 38085 161859 38113
rect 161887 38085 161921 38113
rect 161949 38085 161984 38113
rect 161824 38051 161984 38085
rect 161824 38023 161859 38051
rect 161887 38023 161921 38051
rect 161949 38023 161984 38051
rect 161824 37989 161984 38023
rect 161824 37961 161859 37989
rect 161887 37961 161921 37989
rect 161949 37961 161984 37989
rect 161824 37944 161984 37961
rect 171669 38175 171979 46961
rect 171669 38147 171717 38175
rect 171745 38147 171779 38175
rect 171807 38147 171841 38175
rect 171869 38147 171903 38175
rect 171931 38147 171979 38175
rect 171669 38113 171979 38147
rect 171669 38085 171717 38113
rect 171745 38085 171779 38113
rect 171807 38085 171841 38113
rect 171869 38085 171903 38113
rect 171931 38085 171979 38113
rect 171669 38051 171979 38085
rect 171669 38023 171717 38051
rect 171745 38023 171779 38051
rect 171807 38023 171841 38051
rect 171869 38023 171903 38051
rect 171931 38023 171979 38051
rect 171669 37989 171979 38023
rect 171669 37961 171717 37989
rect 171745 37961 171779 37989
rect 171807 37961 171841 37989
rect 171869 37961 171903 37989
rect 171931 37961 171979 37989
rect 158169 32147 158217 32175
rect 158245 32147 158279 32175
rect 158307 32147 158341 32175
rect 158369 32147 158403 32175
rect 158431 32147 158479 32175
rect 158169 32113 158479 32147
rect 158169 32085 158217 32113
rect 158245 32085 158279 32113
rect 158307 32085 158341 32113
rect 158369 32085 158403 32113
rect 158431 32085 158479 32113
rect 158169 32051 158479 32085
rect 158169 32023 158217 32051
rect 158245 32023 158279 32051
rect 158307 32023 158341 32051
rect 158369 32023 158403 32051
rect 158431 32023 158479 32051
rect 158169 31989 158479 32023
rect 158169 31961 158217 31989
rect 158245 31961 158279 31989
rect 158307 31961 158341 31989
rect 158369 31961 158403 31989
rect 158431 31961 158479 31989
rect 158169 23175 158479 31961
rect 169504 32175 169664 32192
rect 169504 32147 169539 32175
rect 169567 32147 169601 32175
rect 169629 32147 169664 32175
rect 169504 32113 169664 32147
rect 169504 32085 169539 32113
rect 169567 32085 169601 32113
rect 169629 32085 169664 32113
rect 169504 32051 169664 32085
rect 169504 32023 169539 32051
rect 169567 32023 169601 32051
rect 169629 32023 169664 32051
rect 169504 31989 169664 32023
rect 169504 31961 169539 31989
rect 169567 31961 169601 31989
rect 169629 31961 169664 31989
rect 169504 31944 169664 31961
rect 161824 29175 161984 29192
rect 161824 29147 161859 29175
rect 161887 29147 161921 29175
rect 161949 29147 161984 29175
rect 161824 29113 161984 29147
rect 161824 29085 161859 29113
rect 161887 29085 161921 29113
rect 161949 29085 161984 29113
rect 161824 29051 161984 29085
rect 161824 29023 161859 29051
rect 161887 29023 161921 29051
rect 161949 29023 161984 29051
rect 161824 28989 161984 29023
rect 161824 28961 161859 28989
rect 161887 28961 161921 28989
rect 161949 28961 161984 28989
rect 161824 28944 161984 28961
rect 171669 29175 171979 37961
rect 171669 29147 171717 29175
rect 171745 29147 171779 29175
rect 171807 29147 171841 29175
rect 171869 29147 171903 29175
rect 171931 29147 171979 29175
rect 171669 29113 171979 29147
rect 171669 29085 171717 29113
rect 171745 29085 171779 29113
rect 171807 29085 171841 29113
rect 171869 29085 171903 29113
rect 171931 29085 171979 29113
rect 171669 29051 171979 29085
rect 171669 29023 171717 29051
rect 171745 29023 171779 29051
rect 171807 29023 171841 29051
rect 171869 29023 171903 29051
rect 171931 29023 171979 29051
rect 171669 28989 171979 29023
rect 171669 28961 171717 28989
rect 171745 28961 171779 28989
rect 171807 28961 171841 28989
rect 171869 28961 171903 28989
rect 171931 28961 171979 28989
rect 158169 23147 158217 23175
rect 158245 23147 158279 23175
rect 158307 23147 158341 23175
rect 158369 23147 158403 23175
rect 158431 23147 158479 23175
rect 158169 23113 158479 23147
rect 158169 23085 158217 23113
rect 158245 23085 158279 23113
rect 158307 23085 158341 23113
rect 158369 23085 158403 23113
rect 158431 23085 158479 23113
rect 158169 23051 158479 23085
rect 158169 23023 158217 23051
rect 158245 23023 158279 23051
rect 158307 23023 158341 23051
rect 158369 23023 158403 23051
rect 158431 23023 158479 23051
rect 158169 22989 158479 23023
rect 158169 22961 158217 22989
rect 158245 22961 158279 22989
rect 158307 22961 158341 22989
rect 158369 22961 158403 22989
rect 158431 22961 158479 22989
rect 158169 14175 158479 22961
rect 169504 23175 169664 23192
rect 169504 23147 169539 23175
rect 169567 23147 169601 23175
rect 169629 23147 169664 23175
rect 169504 23113 169664 23147
rect 169504 23085 169539 23113
rect 169567 23085 169601 23113
rect 169629 23085 169664 23113
rect 169504 23051 169664 23085
rect 169504 23023 169539 23051
rect 169567 23023 169601 23051
rect 169629 23023 169664 23051
rect 169504 22989 169664 23023
rect 169504 22961 169539 22989
rect 169567 22961 169601 22989
rect 169629 22961 169664 22989
rect 169504 22944 169664 22961
rect 161824 20175 161984 20192
rect 161824 20147 161859 20175
rect 161887 20147 161921 20175
rect 161949 20147 161984 20175
rect 161824 20113 161984 20147
rect 161824 20085 161859 20113
rect 161887 20085 161921 20113
rect 161949 20085 161984 20113
rect 161824 20051 161984 20085
rect 161824 20023 161859 20051
rect 161887 20023 161921 20051
rect 161949 20023 161984 20051
rect 161824 19989 161984 20023
rect 161824 19961 161859 19989
rect 161887 19961 161921 19989
rect 161949 19961 161984 19989
rect 161824 19944 161984 19961
rect 171669 20175 171979 28961
rect 171669 20147 171717 20175
rect 171745 20147 171779 20175
rect 171807 20147 171841 20175
rect 171869 20147 171903 20175
rect 171931 20147 171979 20175
rect 171669 20113 171979 20147
rect 171669 20085 171717 20113
rect 171745 20085 171779 20113
rect 171807 20085 171841 20113
rect 171869 20085 171903 20113
rect 171931 20085 171979 20113
rect 171669 20051 171979 20085
rect 171669 20023 171717 20051
rect 171745 20023 171779 20051
rect 171807 20023 171841 20051
rect 171869 20023 171903 20051
rect 171931 20023 171979 20051
rect 171669 19989 171979 20023
rect 171669 19961 171717 19989
rect 171745 19961 171779 19989
rect 171807 19961 171841 19989
rect 171869 19961 171903 19989
rect 171931 19961 171979 19989
rect 158169 14147 158217 14175
rect 158245 14147 158279 14175
rect 158307 14147 158341 14175
rect 158369 14147 158403 14175
rect 158431 14147 158479 14175
rect 158169 14113 158479 14147
rect 158169 14085 158217 14113
rect 158245 14085 158279 14113
rect 158307 14085 158341 14113
rect 158369 14085 158403 14113
rect 158431 14085 158479 14113
rect 158169 14051 158479 14085
rect 158169 14023 158217 14051
rect 158245 14023 158279 14051
rect 158307 14023 158341 14051
rect 158369 14023 158403 14051
rect 158431 14023 158479 14051
rect 158169 13989 158479 14023
rect 158169 13961 158217 13989
rect 158245 13961 158279 13989
rect 158307 13961 158341 13989
rect 158369 13961 158403 13989
rect 158431 13961 158479 13989
rect 158169 5175 158479 13961
rect 169504 14175 169664 14192
rect 169504 14147 169539 14175
rect 169567 14147 169601 14175
rect 169629 14147 169664 14175
rect 169504 14113 169664 14147
rect 169504 14085 169539 14113
rect 169567 14085 169601 14113
rect 169629 14085 169664 14113
rect 169504 14051 169664 14085
rect 169504 14023 169539 14051
rect 169567 14023 169601 14051
rect 169629 14023 169664 14051
rect 169504 13989 169664 14023
rect 169504 13961 169539 13989
rect 169567 13961 169601 13989
rect 169629 13961 169664 13989
rect 169504 13944 169664 13961
rect 161824 11175 161984 11192
rect 161824 11147 161859 11175
rect 161887 11147 161921 11175
rect 161949 11147 161984 11175
rect 161824 11113 161984 11147
rect 161824 11085 161859 11113
rect 161887 11085 161921 11113
rect 161949 11085 161984 11113
rect 161824 11051 161984 11085
rect 161824 11023 161859 11051
rect 161887 11023 161921 11051
rect 161949 11023 161984 11051
rect 161824 10989 161984 11023
rect 161824 10961 161859 10989
rect 161887 10961 161921 10989
rect 161949 10961 161984 10989
rect 161824 10944 161984 10961
rect 171669 11175 171979 19961
rect 171669 11147 171717 11175
rect 171745 11147 171779 11175
rect 171807 11147 171841 11175
rect 171869 11147 171903 11175
rect 171931 11147 171979 11175
rect 171669 11113 171979 11147
rect 171669 11085 171717 11113
rect 171745 11085 171779 11113
rect 171807 11085 171841 11113
rect 171869 11085 171903 11113
rect 171931 11085 171979 11113
rect 171669 11051 171979 11085
rect 171669 11023 171717 11051
rect 171745 11023 171779 11051
rect 171807 11023 171841 11051
rect 171869 11023 171903 11051
rect 171931 11023 171979 11051
rect 171669 10989 171979 11023
rect 171669 10961 171717 10989
rect 171745 10961 171779 10989
rect 171807 10961 171841 10989
rect 171869 10961 171903 10989
rect 171931 10961 171979 10989
rect 158169 5147 158217 5175
rect 158245 5147 158279 5175
rect 158307 5147 158341 5175
rect 158369 5147 158403 5175
rect 158431 5147 158479 5175
rect 158169 5113 158479 5147
rect 158169 5085 158217 5113
rect 158245 5085 158279 5113
rect 158307 5085 158341 5113
rect 158369 5085 158403 5113
rect 158431 5085 158479 5113
rect 158169 5051 158479 5085
rect 158169 5023 158217 5051
rect 158245 5023 158279 5051
rect 158307 5023 158341 5051
rect 158369 5023 158403 5051
rect 158431 5023 158479 5051
rect 158169 4989 158479 5023
rect 158169 4961 158217 4989
rect 158245 4961 158279 4989
rect 158307 4961 158341 4989
rect 158369 4961 158403 4989
rect 158431 4961 158479 4989
rect 158169 -560 158479 4961
rect 169504 5175 169664 5192
rect 169504 5147 169539 5175
rect 169567 5147 169601 5175
rect 169629 5147 169664 5175
rect 169504 5113 169664 5147
rect 169504 5085 169539 5113
rect 169567 5085 169601 5113
rect 169629 5085 169664 5113
rect 169504 5051 169664 5085
rect 169504 5023 169539 5051
rect 169567 5023 169601 5051
rect 169629 5023 169664 5051
rect 169504 4989 169664 5023
rect 169504 4961 169539 4989
rect 169567 4961 169601 4989
rect 169629 4961 169664 4989
rect 169504 4944 169664 4961
rect 158169 -588 158217 -560
rect 158245 -588 158279 -560
rect 158307 -588 158341 -560
rect 158369 -588 158403 -560
rect 158431 -588 158479 -560
rect 158169 -622 158479 -588
rect 158169 -650 158217 -622
rect 158245 -650 158279 -622
rect 158307 -650 158341 -622
rect 158369 -650 158403 -622
rect 158431 -650 158479 -622
rect 158169 -684 158479 -650
rect 158169 -712 158217 -684
rect 158245 -712 158279 -684
rect 158307 -712 158341 -684
rect 158369 -712 158403 -684
rect 158431 -712 158479 -684
rect 158169 -746 158479 -712
rect 158169 -774 158217 -746
rect 158245 -774 158279 -746
rect 158307 -774 158341 -746
rect 158369 -774 158403 -746
rect 158431 -774 158479 -746
rect 158169 -822 158479 -774
rect 171669 2175 171979 10961
rect 171669 2147 171717 2175
rect 171745 2147 171779 2175
rect 171807 2147 171841 2175
rect 171869 2147 171903 2175
rect 171931 2147 171979 2175
rect 171669 2113 171979 2147
rect 171669 2085 171717 2113
rect 171745 2085 171779 2113
rect 171807 2085 171841 2113
rect 171869 2085 171903 2113
rect 171931 2085 171979 2113
rect 171669 2051 171979 2085
rect 171669 2023 171717 2051
rect 171745 2023 171779 2051
rect 171807 2023 171841 2051
rect 171869 2023 171903 2051
rect 171931 2023 171979 2051
rect 171669 1989 171979 2023
rect 171669 1961 171717 1989
rect 171745 1961 171779 1989
rect 171807 1961 171841 1989
rect 171869 1961 171903 1989
rect 171931 1961 171979 1989
rect 171669 -80 171979 1961
rect 171669 -108 171717 -80
rect 171745 -108 171779 -80
rect 171807 -108 171841 -80
rect 171869 -108 171903 -80
rect 171931 -108 171979 -80
rect 171669 -142 171979 -108
rect 171669 -170 171717 -142
rect 171745 -170 171779 -142
rect 171807 -170 171841 -142
rect 171869 -170 171903 -142
rect 171931 -170 171979 -142
rect 171669 -204 171979 -170
rect 171669 -232 171717 -204
rect 171745 -232 171779 -204
rect 171807 -232 171841 -204
rect 171869 -232 171903 -204
rect 171931 -232 171979 -204
rect 171669 -266 171979 -232
rect 171669 -294 171717 -266
rect 171745 -294 171779 -266
rect 171807 -294 171841 -266
rect 171869 -294 171903 -266
rect 171931 -294 171979 -266
rect 171669 -822 171979 -294
rect 173529 299086 173839 299134
rect 173529 299058 173577 299086
rect 173605 299058 173639 299086
rect 173667 299058 173701 299086
rect 173729 299058 173763 299086
rect 173791 299058 173839 299086
rect 173529 299024 173839 299058
rect 173529 298996 173577 299024
rect 173605 298996 173639 299024
rect 173667 298996 173701 299024
rect 173729 298996 173763 299024
rect 173791 298996 173839 299024
rect 173529 298962 173839 298996
rect 173529 298934 173577 298962
rect 173605 298934 173639 298962
rect 173667 298934 173701 298962
rect 173729 298934 173763 298962
rect 173791 298934 173839 298962
rect 173529 298900 173839 298934
rect 173529 298872 173577 298900
rect 173605 298872 173639 298900
rect 173667 298872 173701 298900
rect 173729 298872 173763 298900
rect 173791 298872 173839 298900
rect 173529 293175 173839 298872
rect 173529 293147 173577 293175
rect 173605 293147 173639 293175
rect 173667 293147 173701 293175
rect 173729 293147 173763 293175
rect 173791 293147 173839 293175
rect 173529 293113 173839 293147
rect 173529 293085 173577 293113
rect 173605 293085 173639 293113
rect 173667 293085 173701 293113
rect 173729 293085 173763 293113
rect 173791 293085 173839 293113
rect 173529 293051 173839 293085
rect 173529 293023 173577 293051
rect 173605 293023 173639 293051
rect 173667 293023 173701 293051
rect 173729 293023 173763 293051
rect 173791 293023 173839 293051
rect 173529 292989 173839 293023
rect 173529 292961 173577 292989
rect 173605 292961 173639 292989
rect 173667 292961 173701 292989
rect 173729 292961 173763 292989
rect 173791 292961 173839 292989
rect 173529 284175 173839 292961
rect 173529 284147 173577 284175
rect 173605 284147 173639 284175
rect 173667 284147 173701 284175
rect 173729 284147 173763 284175
rect 173791 284147 173839 284175
rect 173529 284113 173839 284147
rect 173529 284085 173577 284113
rect 173605 284085 173639 284113
rect 173667 284085 173701 284113
rect 173729 284085 173763 284113
rect 173791 284085 173839 284113
rect 173529 284051 173839 284085
rect 173529 284023 173577 284051
rect 173605 284023 173639 284051
rect 173667 284023 173701 284051
rect 173729 284023 173763 284051
rect 173791 284023 173839 284051
rect 173529 283989 173839 284023
rect 173529 283961 173577 283989
rect 173605 283961 173639 283989
rect 173667 283961 173701 283989
rect 173729 283961 173763 283989
rect 173791 283961 173839 283989
rect 173529 275175 173839 283961
rect 173529 275147 173577 275175
rect 173605 275147 173639 275175
rect 173667 275147 173701 275175
rect 173729 275147 173763 275175
rect 173791 275147 173839 275175
rect 173529 275113 173839 275147
rect 173529 275085 173577 275113
rect 173605 275085 173639 275113
rect 173667 275085 173701 275113
rect 173729 275085 173763 275113
rect 173791 275085 173839 275113
rect 173529 275051 173839 275085
rect 173529 275023 173577 275051
rect 173605 275023 173639 275051
rect 173667 275023 173701 275051
rect 173729 275023 173763 275051
rect 173791 275023 173839 275051
rect 173529 274989 173839 275023
rect 173529 274961 173577 274989
rect 173605 274961 173639 274989
rect 173667 274961 173701 274989
rect 173729 274961 173763 274989
rect 173791 274961 173839 274989
rect 173529 266175 173839 274961
rect 173529 266147 173577 266175
rect 173605 266147 173639 266175
rect 173667 266147 173701 266175
rect 173729 266147 173763 266175
rect 173791 266147 173839 266175
rect 173529 266113 173839 266147
rect 173529 266085 173577 266113
rect 173605 266085 173639 266113
rect 173667 266085 173701 266113
rect 173729 266085 173763 266113
rect 173791 266085 173839 266113
rect 173529 266051 173839 266085
rect 173529 266023 173577 266051
rect 173605 266023 173639 266051
rect 173667 266023 173701 266051
rect 173729 266023 173763 266051
rect 173791 266023 173839 266051
rect 173529 265989 173839 266023
rect 173529 265961 173577 265989
rect 173605 265961 173639 265989
rect 173667 265961 173701 265989
rect 173729 265961 173763 265989
rect 173791 265961 173839 265989
rect 173529 257175 173839 265961
rect 173529 257147 173577 257175
rect 173605 257147 173639 257175
rect 173667 257147 173701 257175
rect 173729 257147 173763 257175
rect 173791 257147 173839 257175
rect 173529 257113 173839 257147
rect 173529 257085 173577 257113
rect 173605 257085 173639 257113
rect 173667 257085 173701 257113
rect 173729 257085 173763 257113
rect 173791 257085 173839 257113
rect 173529 257051 173839 257085
rect 173529 257023 173577 257051
rect 173605 257023 173639 257051
rect 173667 257023 173701 257051
rect 173729 257023 173763 257051
rect 173791 257023 173839 257051
rect 173529 256989 173839 257023
rect 173529 256961 173577 256989
rect 173605 256961 173639 256989
rect 173667 256961 173701 256989
rect 173729 256961 173763 256989
rect 173791 256961 173839 256989
rect 173529 248175 173839 256961
rect 173529 248147 173577 248175
rect 173605 248147 173639 248175
rect 173667 248147 173701 248175
rect 173729 248147 173763 248175
rect 173791 248147 173839 248175
rect 173529 248113 173839 248147
rect 173529 248085 173577 248113
rect 173605 248085 173639 248113
rect 173667 248085 173701 248113
rect 173729 248085 173763 248113
rect 173791 248085 173839 248113
rect 173529 248051 173839 248085
rect 173529 248023 173577 248051
rect 173605 248023 173639 248051
rect 173667 248023 173701 248051
rect 173729 248023 173763 248051
rect 173791 248023 173839 248051
rect 173529 247989 173839 248023
rect 173529 247961 173577 247989
rect 173605 247961 173639 247989
rect 173667 247961 173701 247989
rect 173729 247961 173763 247989
rect 173791 247961 173839 247989
rect 173529 239175 173839 247961
rect 173529 239147 173577 239175
rect 173605 239147 173639 239175
rect 173667 239147 173701 239175
rect 173729 239147 173763 239175
rect 173791 239147 173839 239175
rect 173529 239113 173839 239147
rect 173529 239085 173577 239113
rect 173605 239085 173639 239113
rect 173667 239085 173701 239113
rect 173729 239085 173763 239113
rect 173791 239085 173839 239113
rect 173529 239051 173839 239085
rect 173529 239023 173577 239051
rect 173605 239023 173639 239051
rect 173667 239023 173701 239051
rect 173729 239023 173763 239051
rect 173791 239023 173839 239051
rect 173529 238989 173839 239023
rect 173529 238961 173577 238989
rect 173605 238961 173639 238989
rect 173667 238961 173701 238989
rect 173729 238961 173763 238989
rect 173791 238961 173839 238989
rect 173529 230175 173839 238961
rect 173529 230147 173577 230175
rect 173605 230147 173639 230175
rect 173667 230147 173701 230175
rect 173729 230147 173763 230175
rect 173791 230147 173839 230175
rect 173529 230113 173839 230147
rect 173529 230085 173577 230113
rect 173605 230085 173639 230113
rect 173667 230085 173701 230113
rect 173729 230085 173763 230113
rect 173791 230085 173839 230113
rect 173529 230051 173839 230085
rect 173529 230023 173577 230051
rect 173605 230023 173639 230051
rect 173667 230023 173701 230051
rect 173729 230023 173763 230051
rect 173791 230023 173839 230051
rect 173529 229989 173839 230023
rect 173529 229961 173577 229989
rect 173605 229961 173639 229989
rect 173667 229961 173701 229989
rect 173729 229961 173763 229989
rect 173791 229961 173839 229989
rect 173529 221175 173839 229961
rect 173529 221147 173577 221175
rect 173605 221147 173639 221175
rect 173667 221147 173701 221175
rect 173729 221147 173763 221175
rect 173791 221147 173839 221175
rect 173529 221113 173839 221147
rect 173529 221085 173577 221113
rect 173605 221085 173639 221113
rect 173667 221085 173701 221113
rect 173729 221085 173763 221113
rect 173791 221085 173839 221113
rect 173529 221051 173839 221085
rect 173529 221023 173577 221051
rect 173605 221023 173639 221051
rect 173667 221023 173701 221051
rect 173729 221023 173763 221051
rect 173791 221023 173839 221051
rect 173529 220989 173839 221023
rect 173529 220961 173577 220989
rect 173605 220961 173639 220989
rect 173667 220961 173701 220989
rect 173729 220961 173763 220989
rect 173791 220961 173839 220989
rect 173529 212175 173839 220961
rect 173529 212147 173577 212175
rect 173605 212147 173639 212175
rect 173667 212147 173701 212175
rect 173729 212147 173763 212175
rect 173791 212147 173839 212175
rect 173529 212113 173839 212147
rect 173529 212085 173577 212113
rect 173605 212085 173639 212113
rect 173667 212085 173701 212113
rect 173729 212085 173763 212113
rect 173791 212085 173839 212113
rect 173529 212051 173839 212085
rect 173529 212023 173577 212051
rect 173605 212023 173639 212051
rect 173667 212023 173701 212051
rect 173729 212023 173763 212051
rect 173791 212023 173839 212051
rect 173529 211989 173839 212023
rect 173529 211961 173577 211989
rect 173605 211961 173639 211989
rect 173667 211961 173701 211989
rect 173729 211961 173763 211989
rect 173791 211961 173839 211989
rect 173529 203175 173839 211961
rect 173529 203147 173577 203175
rect 173605 203147 173639 203175
rect 173667 203147 173701 203175
rect 173729 203147 173763 203175
rect 173791 203147 173839 203175
rect 173529 203113 173839 203147
rect 173529 203085 173577 203113
rect 173605 203085 173639 203113
rect 173667 203085 173701 203113
rect 173729 203085 173763 203113
rect 173791 203085 173839 203113
rect 173529 203051 173839 203085
rect 173529 203023 173577 203051
rect 173605 203023 173639 203051
rect 173667 203023 173701 203051
rect 173729 203023 173763 203051
rect 173791 203023 173839 203051
rect 173529 202989 173839 203023
rect 173529 202961 173577 202989
rect 173605 202961 173639 202989
rect 173667 202961 173701 202989
rect 173729 202961 173763 202989
rect 173791 202961 173839 202989
rect 173529 194175 173839 202961
rect 173529 194147 173577 194175
rect 173605 194147 173639 194175
rect 173667 194147 173701 194175
rect 173729 194147 173763 194175
rect 173791 194147 173839 194175
rect 173529 194113 173839 194147
rect 173529 194085 173577 194113
rect 173605 194085 173639 194113
rect 173667 194085 173701 194113
rect 173729 194085 173763 194113
rect 173791 194085 173839 194113
rect 173529 194051 173839 194085
rect 173529 194023 173577 194051
rect 173605 194023 173639 194051
rect 173667 194023 173701 194051
rect 173729 194023 173763 194051
rect 173791 194023 173839 194051
rect 173529 193989 173839 194023
rect 173529 193961 173577 193989
rect 173605 193961 173639 193989
rect 173667 193961 173701 193989
rect 173729 193961 173763 193989
rect 173791 193961 173839 193989
rect 173529 185175 173839 193961
rect 173529 185147 173577 185175
rect 173605 185147 173639 185175
rect 173667 185147 173701 185175
rect 173729 185147 173763 185175
rect 173791 185147 173839 185175
rect 173529 185113 173839 185147
rect 173529 185085 173577 185113
rect 173605 185085 173639 185113
rect 173667 185085 173701 185113
rect 173729 185085 173763 185113
rect 173791 185085 173839 185113
rect 173529 185051 173839 185085
rect 173529 185023 173577 185051
rect 173605 185023 173639 185051
rect 173667 185023 173701 185051
rect 173729 185023 173763 185051
rect 173791 185023 173839 185051
rect 173529 184989 173839 185023
rect 173529 184961 173577 184989
rect 173605 184961 173639 184989
rect 173667 184961 173701 184989
rect 173729 184961 173763 184989
rect 173791 184961 173839 184989
rect 173529 176175 173839 184961
rect 173529 176147 173577 176175
rect 173605 176147 173639 176175
rect 173667 176147 173701 176175
rect 173729 176147 173763 176175
rect 173791 176147 173839 176175
rect 173529 176113 173839 176147
rect 173529 176085 173577 176113
rect 173605 176085 173639 176113
rect 173667 176085 173701 176113
rect 173729 176085 173763 176113
rect 173791 176085 173839 176113
rect 173529 176051 173839 176085
rect 173529 176023 173577 176051
rect 173605 176023 173639 176051
rect 173667 176023 173701 176051
rect 173729 176023 173763 176051
rect 173791 176023 173839 176051
rect 173529 175989 173839 176023
rect 173529 175961 173577 175989
rect 173605 175961 173639 175989
rect 173667 175961 173701 175989
rect 173729 175961 173763 175989
rect 173791 175961 173839 175989
rect 173529 167175 173839 175961
rect 187029 298606 187339 299134
rect 187029 298578 187077 298606
rect 187105 298578 187139 298606
rect 187167 298578 187201 298606
rect 187229 298578 187263 298606
rect 187291 298578 187339 298606
rect 187029 298544 187339 298578
rect 187029 298516 187077 298544
rect 187105 298516 187139 298544
rect 187167 298516 187201 298544
rect 187229 298516 187263 298544
rect 187291 298516 187339 298544
rect 187029 298482 187339 298516
rect 187029 298454 187077 298482
rect 187105 298454 187139 298482
rect 187167 298454 187201 298482
rect 187229 298454 187263 298482
rect 187291 298454 187339 298482
rect 187029 298420 187339 298454
rect 187029 298392 187077 298420
rect 187105 298392 187139 298420
rect 187167 298392 187201 298420
rect 187229 298392 187263 298420
rect 187291 298392 187339 298420
rect 187029 290175 187339 298392
rect 187029 290147 187077 290175
rect 187105 290147 187139 290175
rect 187167 290147 187201 290175
rect 187229 290147 187263 290175
rect 187291 290147 187339 290175
rect 187029 290113 187339 290147
rect 187029 290085 187077 290113
rect 187105 290085 187139 290113
rect 187167 290085 187201 290113
rect 187229 290085 187263 290113
rect 187291 290085 187339 290113
rect 187029 290051 187339 290085
rect 187029 290023 187077 290051
rect 187105 290023 187139 290051
rect 187167 290023 187201 290051
rect 187229 290023 187263 290051
rect 187291 290023 187339 290051
rect 187029 289989 187339 290023
rect 187029 289961 187077 289989
rect 187105 289961 187139 289989
rect 187167 289961 187201 289989
rect 187229 289961 187263 289989
rect 187291 289961 187339 289989
rect 187029 281175 187339 289961
rect 187029 281147 187077 281175
rect 187105 281147 187139 281175
rect 187167 281147 187201 281175
rect 187229 281147 187263 281175
rect 187291 281147 187339 281175
rect 187029 281113 187339 281147
rect 187029 281085 187077 281113
rect 187105 281085 187139 281113
rect 187167 281085 187201 281113
rect 187229 281085 187263 281113
rect 187291 281085 187339 281113
rect 187029 281051 187339 281085
rect 187029 281023 187077 281051
rect 187105 281023 187139 281051
rect 187167 281023 187201 281051
rect 187229 281023 187263 281051
rect 187291 281023 187339 281051
rect 187029 280989 187339 281023
rect 187029 280961 187077 280989
rect 187105 280961 187139 280989
rect 187167 280961 187201 280989
rect 187229 280961 187263 280989
rect 187291 280961 187339 280989
rect 187029 272175 187339 280961
rect 187029 272147 187077 272175
rect 187105 272147 187139 272175
rect 187167 272147 187201 272175
rect 187229 272147 187263 272175
rect 187291 272147 187339 272175
rect 187029 272113 187339 272147
rect 187029 272085 187077 272113
rect 187105 272085 187139 272113
rect 187167 272085 187201 272113
rect 187229 272085 187263 272113
rect 187291 272085 187339 272113
rect 187029 272051 187339 272085
rect 187029 272023 187077 272051
rect 187105 272023 187139 272051
rect 187167 272023 187201 272051
rect 187229 272023 187263 272051
rect 187291 272023 187339 272051
rect 187029 271989 187339 272023
rect 187029 271961 187077 271989
rect 187105 271961 187139 271989
rect 187167 271961 187201 271989
rect 187229 271961 187263 271989
rect 187291 271961 187339 271989
rect 187029 263175 187339 271961
rect 187029 263147 187077 263175
rect 187105 263147 187139 263175
rect 187167 263147 187201 263175
rect 187229 263147 187263 263175
rect 187291 263147 187339 263175
rect 187029 263113 187339 263147
rect 187029 263085 187077 263113
rect 187105 263085 187139 263113
rect 187167 263085 187201 263113
rect 187229 263085 187263 263113
rect 187291 263085 187339 263113
rect 187029 263051 187339 263085
rect 187029 263023 187077 263051
rect 187105 263023 187139 263051
rect 187167 263023 187201 263051
rect 187229 263023 187263 263051
rect 187291 263023 187339 263051
rect 187029 262989 187339 263023
rect 187029 262961 187077 262989
rect 187105 262961 187139 262989
rect 187167 262961 187201 262989
rect 187229 262961 187263 262989
rect 187291 262961 187339 262989
rect 187029 254175 187339 262961
rect 187029 254147 187077 254175
rect 187105 254147 187139 254175
rect 187167 254147 187201 254175
rect 187229 254147 187263 254175
rect 187291 254147 187339 254175
rect 187029 254113 187339 254147
rect 187029 254085 187077 254113
rect 187105 254085 187139 254113
rect 187167 254085 187201 254113
rect 187229 254085 187263 254113
rect 187291 254085 187339 254113
rect 187029 254051 187339 254085
rect 187029 254023 187077 254051
rect 187105 254023 187139 254051
rect 187167 254023 187201 254051
rect 187229 254023 187263 254051
rect 187291 254023 187339 254051
rect 187029 253989 187339 254023
rect 187029 253961 187077 253989
rect 187105 253961 187139 253989
rect 187167 253961 187201 253989
rect 187229 253961 187263 253989
rect 187291 253961 187339 253989
rect 187029 245175 187339 253961
rect 187029 245147 187077 245175
rect 187105 245147 187139 245175
rect 187167 245147 187201 245175
rect 187229 245147 187263 245175
rect 187291 245147 187339 245175
rect 187029 245113 187339 245147
rect 187029 245085 187077 245113
rect 187105 245085 187139 245113
rect 187167 245085 187201 245113
rect 187229 245085 187263 245113
rect 187291 245085 187339 245113
rect 187029 245051 187339 245085
rect 187029 245023 187077 245051
rect 187105 245023 187139 245051
rect 187167 245023 187201 245051
rect 187229 245023 187263 245051
rect 187291 245023 187339 245051
rect 187029 244989 187339 245023
rect 187029 244961 187077 244989
rect 187105 244961 187139 244989
rect 187167 244961 187201 244989
rect 187229 244961 187263 244989
rect 187291 244961 187339 244989
rect 187029 236175 187339 244961
rect 187029 236147 187077 236175
rect 187105 236147 187139 236175
rect 187167 236147 187201 236175
rect 187229 236147 187263 236175
rect 187291 236147 187339 236175
rect 187029 236113 187339 236147
rect 187029 236085 187077 236113
rect 187105 236085 187139 236113
rect 187167 236085 187201 236113
rect 187229 236085 187263 236113
rect 187291 236085 187339 236113
rect 187029 236051 187339 236085
rect 187029 236023 187077 236051
rect 187105 236023 187139 236051
rect 187167 236023 187201 236051
rect 187229 236023 187263 236051
rect 187291 236023 187339 236051
rect 187029 235989 187339 236023
rect 187029 235961 187077 235989
rect 187105 235961 187139 235989
rect 187167 235961 187201 235989
rect 187229 235961 187263 235989
rect 187291 235961 187339 235989
rect 187029 227175 187339 235961
rect 187029 227147 187077 227175
rect 187105 227147 187139 227175
rect 187167 227147 187201 227175
rect 187229 227147 187263 227175
rect 187291 227147 187339 227175
rect 187029 227113 187339 227147
rect 187029 227085 187077 227113
rect 187105 227085 187139 227113
rect 187167 227085 187201 227113
rect 187229 227085 187263 227113
rect 187291 227085 187339 227113
rect 187029 227051 187339 227085
rect 187029 227023 187077 227051
rect 187105 227023 187139 227051
rect 187167 227023 187201 227051
rect 187229 227023 187263 227051
rect 187291 227023 187339 227051
rect 187029 226989 187339 227023
rect 187029 226961 187077 226989
rect 187105 226961 187139 226989
rect 187167 226961 187201 226989
rect 187229 226961 187263 226989
rect 187291 226961 187339 226989
rect 187029 218175 187339 226961
rect 187029 218147 187077 218175
rect 187105 218147 187139 218175
rect 187167 218147 187201 218175
rect 187229 218147 187263 218175
rect 187291 218147 187339 218175
rect 187029 218113 187339 218147
rect 187029 218085 187077 218113
rect 187105 218085 187139 218113
rect 187167 218085 187201 218113
rect 187229 218085 187263 218113
rect 187291 218085 187339 218113
rect 187029 218051 187339 218085
rect 187029 218023 187077 218051
rect 187105 218023 187139 218051
rect 187167 218023 187201 218051
rect 187229 218023 187263 218051
rect 187291 218023 187339 218051
rect 187029 217989 187339 218023
rect 187029 217961 187077 217989
rect 187105 217961 187139 217989
rect 187167 217961 187201 217989
rect 187229 217961 187263 217989
rect 187291 217961 187339 217989
rect 187029 209175 187339 217961
rect 187029 209147 187077 209175
rect 187105 209147 187139 209175
rect 187167 209147 187201 209175
rect 187229 209147 187263 209175
rect 187291 209147 187339 209175
rect 187029 209113 187339 209147
rect 187029 209085 187077 209113
rect 187105 209085 187139 209113
rect 187167 209085 187201 209113
rect 187229 209085 187263 209113
rect 187291 209085 187339 209113
rect 187029 209051 187339 209085
rect 187029 209023 187077 209051
rect 187105 209023 187139 209051
rect 187167 209023 187201 209051
rect 187229 209023 187263 209051
rect 187291 209023 187339 209051
rect 187029 208989 187339 209023
rect 187029 208961 187077 208989
rect 187105 208961 187139 208989
rect 187167 208961 187201 208989
rect 187229 208961 187263 208989
rect 187291 208961 187339 208989
rect 187029 200175 187339 208961
rect 187029 200147 187077 200175
rect 187105 200147 187139 200175
rect 187167 200147 187201 200175
rect 187229 200147 187263 200175
rect 187291 200147 187339 200175
rect 187029 200113 187339 200147
rect 187029 200085 187077 200113
rect 187105 200085 187139 200113
rect 187167 200085 187201 200113
rect 187229 200085 187263 200113
rect 187291 200085 187339 200113
rect 187029 200051 187339 200085
rect 187029 200023 187077 200051
rect 187105 200023 187139 200051
rect 187167 200023 187201 200051
rect 187229 200023 187263 200051
rect 187291 200023 187339 200051
rect 187029 199989 187339 200023
rect 187029 199961 187077 199989
rect 187105 199961 187139 199989
rect 187167 199961 187201 199989
rect 187229 199961 187263 199989
rect 187291 199961 187339 199989
rect 187029 191175 187339 199961
rect 187029 191147 187077 191175
rect 187105 191147 187139 191175
rect 187167 191147 187201 191175
rect 187229 191147 187263 191175
rect 187291 191147 187339 191175
rect 187029 191113 187339 191147
rect 187029 191085 187077 191113
rect 187105 191085 187139 191113
rect 187167 191085 187201 191113
rect 187229 191085 187263 191113
rect 187291 191085 187339 191113
rect 187029 191051 187339 191085
rect 187029 191023 187077 191051
rect 187105 191023 187139 191051
rect 187167 191023 187201 191051
rect 187229 191023 187263 191051
rect 187291 191023 187339 191051
rect 187029 190989 187339 191023
rect 187029 190961 187077 190989
rect 187105 190961 187139 190989
rect 187167 190961 187201 190989
rect 187229 190961 187263 190989
rect 187291 190961 187339 190989
rect 187029 182175 187339 190961
rect 187029 182147 187077 182175
rect 187105 182147 187139 182175
rect 187167 182147 187201 182175
rect 187229 182147 187263 182175
rect 187291 182147 187339 182175
rect 187029 182113 187339 182147
rect 187029 182085 187077 182113
rect 187105 182085 187139 182113
rect 187167 182085 187201 182113
rect 187229 182085 187263 182113
rect 187291 182085 187339 182113
rect 187029 182051 187339 182085
rect 187029 182023 187077 182051
rect 187105 182023 187139 182051
rect 187167 182023 187201 182051
rect 187229 182023 187263 182051
rect 187291 182023 187339 182051
rect 187029 181989 187339 182023
rect 187029 181961 187077 181989
rect 187105 181961 187139 181989
rect 187167 181961 187201 181989
rect 187229 181961 187263 181989
rect 187291 181961 187339 181989
rect 177184 173175 177344 173192
rect 177184 173147 177219 173175
rect 177247 173147 177281 173175
rect 177309 173147 177344 173175
rect 177184 173113 177344 173147
rect 177184 173085 177219 173113
rect 177247 173085 177281 173113
rect 177309 173085 177344 173113
rect 177184 173051 177344 173085
rect 177184 173023 177219 173051
rect 177247 173023 177281 173051
rect 177309 173023 177344 173051
rect 177184 172989 177344 173023
rect 177184 172961 177219 172989
rect 177247 172961 177281 172989
rect 177309 172961 177344 172989
rect 177184 172944 177344 172961
rect 187029 173175 187339 181961
rect 187029 173147 187077 173175
rect 187105 173147 187139 173175
rect 187167 173147 187201 173175
rect 187229 173147 187263 173175
rect 187291 173147 187339 173175
rect 187029 173113 187339 173147
rect 187029 173085 187077 173113
rect 187105 173085 187139 173113
rect 187167 173085 187201 173113
rect 187229 173085 187263 173113
rect 187291 173085 187339 173113
rect 187029 173051 187339 173085
rect 187029 173023 187077 173051
rect 187105 173023 187139 173051
rect 187167 173023 187201 173051
rect 187229 173023 187263 173051
rect 187291 173023 187339 173051
rect 187029 172989 187339 173023
rect 187029 172961 187077 172989
rect 187105 172961 187139 172989
rect 187167 172961 187201 172989
rect 187229 172961 187263 172989
rect 187291 172961 187339 172989
rect 173529 167147 173577 167175
rect 173605 167147 173639 167175
rect 173667 167147 173701 167175
rect 173729 167147 173763 167175
rect 173791 167147 173839 167175
rect 173529 167113 173839 167147
rect 173529 167085 173577 167113
rect 173605 167085 173639 167113
rect 173667 167085 173701 167113
rect 173729 167085 173763 167113
rect 173791 167085 173839 167113
rect 173529 167051 173839 167085
rect 173529 167023 173577 167051
rect 173605 167023 173639 167051
rect 173667 167023 173701 167051
rect 173729 167023 173763 167051
rect 173791 167023 173839 167051
rect 173529 166989 173839 167023
rect 173529 166961 173577 166989
rect 173605 166961 173639 166989
rect 173667 166961 173701 166989
rect 173729 166961 173763 166989
rect 173791 166961 173839 166989
rect 173529 158175 173839 166961
rect 184864 167175 185024 167192
rect 184864 167147 184899 167175
rect 184927 167147 184961 167175
rect 184989 167147 185024 167175
rect 184864 167113 185024 167147
rect 184864 167085 184899 167113
rect 184927 167085 184961 167113
rect 184989 167085 185024 167113
rect 184864 167051 185024 167085
rect 184864 167023 184899 167051
rect 184927 167023 184961 167051
rect 184989 167023 185024 167051
rect 184864 166989 185024 167023
rect 184864 166961 184899 166989
rect 184927 166961 184961 166989
rect 184989 166961 185024 166989
rect 184864 166944 185024 166961
rect 177184 164175 177344 164192
rect 177184 164147 177219 164175
rect 177247 164147 177281 164175
rect 177309 164147 177344 164175
rect 177184 164113 177344 164147
rect 177184 164085 177219 164113
rect 177247 164085 177281 164113
rect 177309 164085 177344 164113
rect 177184 164051 177344 164085
rect 177184 164023 177219 164051
rect 177247 164023 177281 164051
rect 177309 164023 177344 164051
rect 177184 163989 177344 164023
rect 177184 163961 177219 163989
rect 177247 163961 177281 163989
rect 177309 163961 177344 163989
rect 177184 163944 177344 163961
rect 187029 164175 187339 172961
rect 187029 164147 187077 164175
rect 187105 164147 187139 164175
rect 187167 164147 187201 164175
rect 187229 164147 187263 164175
rect 187291 164147 187339 164175
rect 187029 164113 187339 164147
rect 187029 164085 187077 164113
rect 187105 164085 187139 164113
rect 187167 164085 187201 164113
rect 187229 164085 187263 164113
rect 187291 164085 187339 164113
rect 187029 164051 187339 164085
rect 187029 164023 187077 164051
rect 187105 164023 187139 164051
rect 187167 164023 187201 164051
rect 187229 164023 187263 164051
rect 187291 164023 187339 164051
rect 187029 163989 187339 164023
rect 187029 163961 187077 163989
rect 187105 163961 187139 163989
rect 187167 163961 187201 163989
rect 187229 163961 187263 163989
rect 187291 163961 187339 163989
rect 173529 158147 173577 158175
rect 173605 158147 173639 158175
rect 173667 158147 173701 158175
rect 173729 158147 173763 158175
rect 173791 158147 173839 158175
rect 173529 158113 173839 158147
rect 173529 158085 173577 158113
rect 173605 158085 173639 158113
rect 173667 158085 173701 158113
rect 173729 158085 173763 158113
rect 173791 158085 173839 158113
rect 173529 158051 173839 158085
rect 173529 158023 173577 158051
rect 173605 158023 173639 158051
rect 173667 158023 173701 158051
rect 173729 158023 173763 158051
rect 173791 158023 173839 158051
rect 173529 157989 173839 158023
rect 173529 157961 173577 157989
rect 173605 157961 173639 157989
rect 173667 157961 173701 157989
rect 173729 157961 173763 157989
rect 173791 157961 173839 157989
rect 173529 149175 173839 157961
rect 184864 158175 185024 158192
rect 184864 158147 184899 158175
rect 184927 158147 184961 158175
rect 184989 158147 185024 158175
rect 184864 158113 185024 158147
rect 184864 158085 184899 158113
rect 184927 158085 184961 158113
rect 184989 158085 185024 158113
rect 184864 158051 185024 158085
rect 184864 158023 184899 158051
rect 184927 158023 184961 158051
rect 184989 158023 185024 158051
rect 184864 157989 185024 158023
rect 184864 157961 184899 157989
rect 184927 157961 184961 157989
rect 184989 157961 185024 157989
rect 184864 157944 185024 157961
rect 177184 155175 177344 155192
rect 177184 155147 177219 155175
rect 177247 155147 177281 155175
rect 177309 155147 177344 155175
rect 177184 155113 177344 155147
rect 177184 155085 177219 155113
rect 177247 155085 177281 155113
rect 177309 155085 177344 155113
rect 177184 155051 177344 155085
rect 177184 155023 177219 155051
rect 177247 155023 177281 155051
rect 177309 155023 177344 155051
rect 177184 154989 177344 155023
rect 177184 154961 177219 154989
rect 177247 154961 177281 154989
rect 177309 154961 177344 154989
rect 177184 154944 177344 154961
rect 187029 155175 187339 163961
rect 187029 155147 187077 155175
rect 187105 155147 187139 155175
rect 187167 155147 187201 155175
rect 187229 155147 187263 155175
rect 187291 155147 187339 155175
rect 187029 155113 187339 155147
rect 187029 155085 187077 155113
rect 187105 155085 187139 155113
rect 187167 155085 187201 155113
rect 187229 155085 187263 155113
rect 187291 155085 187339 155113
rect 187029 155051 187339 155085
rect 187029 155023 187077 155051
rect 187105 155023 187139 155051
rect 187167 155023 187201 155051
rect 187229 155023 187263 155051
rect 187291 155023 187339 155051
rect 187029 154989 187339 155023
rect 187029 154961 187077 154989
rect 187105 154961 187139 154989
rect 187167 154961 187201 154989
rect 187229 154961 187263 154989
rect 187291 154961 187339 154989
rect 173529 149147 173577 149175
rect 173605 149147 173639 149175
rect 173667 149147 173701 149175
rect 173729 149147 173763 149175
rect 173791 149147 173839 149175
rect 173529 149113 173839 149147
rect 173529 149085 173577 149113
rect 173605 149085 173639 149113
rect 173667 149085 173701 149113
rect 173729 149085 173763 149113
rect 173791 149085 173839 149113
rect 173529 149051 173839 149085
rect 173529 149023 173577 149051
rect 173605 149023 173639 149051
rect 173667 149023 173701 149051
rect 173729 149023 173763 149051
rect 173791 149023 173839 149051
rect 173529 148989 173839 149023
rect 173529 148961 173577 148989
rect 173605 148961 173639 148989
rect 173667 148961 173701 148989
rect 173729 148961 173763 148989
rect 173791 148961 173839 148989
rect 173529 140175 173839 148961
rect 184864 149175 185024 149192
rect 184864 149147 184899 149175
rect 184927 149147 184961 149175
rect 184989 149147 185024 149175
rect 184864 149113 185024 149147
rect 184864 149085 184899 149113
rect 184927 149085 184961 149113
rect 184989 149085 185024 149113
rect 184864 149051 185024 149085
rect 184864 149023 184899 149051
rect 184927 149023 184961 149051
rect 184989 149023 185024 149051
rect 184864 148989 185024 149023
rect 184864 148961 184899 148989
rect 184927 148961 184961 148989
rect 184989 148961 185024 148989
rect 184864 148944 185024 148961
rect 177184 146175 177344 146192
rect 177184 146147 177219 146175
rect 177247 146147 177281 146175
rect 177309 146147 177344 146175
rect 177184 146113 177344 146147
rect 177184 146085 177219 146113
rect 177247 146085 177281 146113
rect 177309 146085 177344 146113
rect 177184 146051 177344 146085
rect 177184 146023 177219 146051
rect 177247 146023 177281 146051
rect 177309 146023 177344 146051
rect 177184 145989 177344 146023
rect 177184 145961 177219 145989
rect 177247 145961 177281 145989
rect 177309 145961 177344 145989
rect 177184 145944 177344 145961
rect 187029 146175 187339 154961
rect 187029 146147 187077 146175
rect 187105 146147 187139 146175
rect 187167 146147 187201 146175
rect 187229 146147 187263 146175
rect 187291 146147 187339 146175
rect 187029 146113 187339 146147
rect 187029 146085 187077 146113
rect 187105 146085 187139 146113
rect 187167 146085 187201 146113
rect 187229 146085 187263 146113
rect 187291 146085 187339 146113
rect 187029 146051 187339 146085
rect 187029 146023 187077 146051
rect 187105 146023 187139 146051
rect 187167 146023 187201 146051
rect 187229 146023 187263 146051
rect 187291 146023 187339 146051
rect 187029 145989 187339 146023
rect 187029 145961 187077 145989
rect 187105 145961 187139 145989
rect 187167 145961 187201 145989
rect 187229 145961 187263 145989
rect 187291 145961 187339 145989
rect 173529 140147 173577 140175
rect 173605 140147 173639 140175
rect 173667 140147 173701 140175
rect 173729 140147 173763 140175
rect 173791 140147 173839 140175
rect 173529 140113 173839 140147
rect 173529 140085 173577 140113
rect 173605 140085 173639 140113
rect 173667 140085 173701 140113
rect 173729 140085 173763 140113
rect 173791 140085 173839 140113
rect 173529 140051 173839 140085
rect 173529 140023 173577 140051
rect 173605 140023 173639 140051
rect 173667 140023 173701 140051
rect 173729 140023 173763 140051
rect 173791 140023 173839 140051
rect 173529 139989 173839 140023
rect 173529 139961 173577 139989
rect 173605 139961 173639 139989
rect 173667 139961 173701 139989
rect 173729 139961 173763 139989
rect 173791 139961 173839 139989
rect 173529 131175 173839 139961
rect 184864 140175 185024 140192
rect 184864 140147 184899 140175
rect 184927 140147 184961 140175
rect 184989 140147 185024 140175
rect 184864 140113 185024 140147
rect 184864 140085 184899 140113
rect 184927 140085 184961 140113
rect 184989 140085 185024 140113
rect 184864 140051 185024 140085
rect 184864 140023 184899 140051
rect 184927 140023 184961 140051
rect 184989 140023 185024 140051
rect 184864 139989 185024 140023
rect 184864 139961 184899 139989
rect 184927 139961 184961 139989
rect 184989 139961 185024 139989
rect 184864 139944 185024 139961
rect 177184 137175 177344 137192
rect 177184 137147 177219 137175
rect 177247 137147 177281 137175
rect 177309 137147 177344 137175
rect 177184 137113 177344 137147
rect 177184 137085 177219 137113
rect 177247 137085 177281 137113
rect 177309 137085 177344 137113
rect 177184 137051 177344 137085
rect 177184 137023 177219 137051
rect 177247 137023 177281 137051
rect 177309 137023 177344 137051
rect 177184 136989 177344 137023
rect 177184 136961 177219 136989
rect 177247 136961 177281 136989
rect 177309 136961 177344 136989
rect 177184 136944 177344 136961
rect 187029 137175 187339 145961
rect 187029 137147 187077 137175
rect 187105 137147 187139 137175
rect 187167 137147 187201 137175
rect 187229 137147 187263 137175
rect 187291 137147 187339 137175
rect 187029 137113 187339 137147
rect 187029 137085 187077 137113
rect 187105 137085 187139 137113
rect 187167 137085 187201 137113
rect 187229 137085 187263 137113
rect 187291 137085 187339 137113
rect 187029 137051 187339 137085
rect 187029 137023 187077 137051
rect 187105 137023 187139 137051
rect 187167 137023 187201 137051
rect 187229 137023 187263 137051
rect 187291 137023 187339 137051
rect 187029 136989 187339 137023
rect 187029 136961 187077 136989
rect 187105 136961 187139 136989
rect 187167 136961 187201 136989
rect 187229 136961 187263 136989
rect 187291 136961 187339 136989
rect 173529 131147 173577 131175
rect 173605 131147 173639 131175
rect 173667 131147 173701 131175
rect 173729 131147 173763 131175
rect 173791 131147 173839 131175
rect 173529 131113 173839 131147
rect 173529 131085 173577 131113
rect 173605 131085 173639 131113
rect 173667 131085 173701 131113
rect 173729 131085 173763 131113
rect 173791 131085 173839 131113
rect 173529 131051 173839 131085
rect 173529 131023 173577 131051
rect 173605 131023 173639 131051
rect 173667 131023 173701 131051
rect 173729 131023 173763 131051
rect 173791 131023 173839 131051
rect 173529 130989 173839 131023
rect 173529 130961 173577 130989
rect 173605 130961 173639 130989
rect 173667 130961 173701 130989
rect 173729 130961 173763 130989
rect 173791 130961 173839 130989
rect 173529 122175 173839 130961
rect 184864 131175 185024 131192
rect 184864 131147 184899 131175
rect 184927 131147 184961 131175
rect 184989 131147 185024 131175
rect 184864 131113 185024 131147
rect 184864 131085 184899 131113
rect 184927 131085 184961 131113
rect 184989 131085 185024 131113
rect 184864 131051 185024 131085
rect 184864 131023 184899 131051
rect 184927 131023 184961 131051
rect 184989 131023 185024 131051
rect 184864 130989 185024 131023
rect 184864 130961 184899 130989
rect 184927 130961 184961 130989
rect 184989 130961 185024 130989
rect 184864 130944 185024 130961
rect 177184 128175 177344 128192
rect 177184 128147 177219 128175
rect 177247 128147 177281 128175
rect 177309 128147 177344 128175
rect 177184 128113 177344 128147
rect 177184 128085 177219 128113
rect 177247 128085 177281 128113
rect 177309 128085 177344 128113
rect 177184 128051 177344 128085
rect 177184 128023 177219 128051
rect 177247 128023 177281 128051
rect 177309 128023 177344 128051
rect 177184 127989 177344 128023
rect 177184 127961 177219 127989
rect 177247 127961 177281 127989
rect 177309 127961 177344 127989
rect 177184 127944 177344 127961
rect 187029 128175 187339 136961
rect 187029 128147 187077 128175
rect 187105 128147 187139 128175
rect 187167 128147 187201 128175
rect 187229 128147 187263 128175
rect 187291 128147 187339 128175
rect 187029 128113 187339 128147
rect 187029 128085 187077 128113
rect 187105 128085 187139 128113
rect 187167 128085 187201 128113
rect 187229 128085 187263 128113
rect 187291 128085 187339 128113
rect 187029 128051 187339 128085
rect 187029 128023 187077 128051
rect 187105 128023 187139 128051
rect 187167 128023 187201 128051
rect 187229 128023 187263 128051
rect 187291 128023 187339 128051
rect 187029 127989 187339 128023
rect 187029 127961 187077 127989
rect 187105 127961 187139 127989
rect 187167 127961 187201 127989
rect 187229 127961 187263 127989
rect 187291 127961 187339 127989
rect 173529 122147 173577 122175
rect 173605 122147 173639 122175
rect 173667 122147 173701 122175
rect 173729 122147 173763 122175
rect 173791 122147 173839 122175
rect 173529 122113 173839 122147
rect 173529 122085 173577 122113
rect 173605 122085 173639 122113
rect 173667 122085 173701 122113
rect 173729 122085 173763 122113
rect 173791 122085 173839 122113
rect 173529 122051 173839 122085
rect 173529 122023 173577 122051
rect 173605 122023 173639 122051
rect 173667 122023 173701 122051
rect 173729 122023 173763 122051
rect 173791 122023 173839 122051
rect 173529 121989 173839 122023
rect 173529 121961 173577 121989
rect 173605 121961 173639 121989
rect 173667 121961 173701 121989
rect 173729 121961 173763 121989
rect 173791 121961 173839 121989
rect 173529 113175 173839 121961
rect 184864 122175 185024 122192
rect 184864 122147 184899 122175
rect 184927 122147 184961 122175
rect 184989 122147 185024 122175
rect 184864 122113 185024 122147
rect 184864 122085 184899 122113
rect 184927 122085 184961 122113
rect 184989 122085 185024 122113
rect 184864 122051 185024 122085
rect 184864 122023 184899 122051
rect 184927 122023 184961 122051
rect 184989 122023 185024 122051
rect 184864 121989 185024 122023
rect 184864 121961 184899 121989
rect 184927 121961 184961 121989
rect 184989 121961 185024 121989
rect 184864 121944 185024 121961
rect 177184 119175 177344 119192
rect 177184 119147 177219 119175
rect 177247 119147 177281 119175
rect 177309 119147 177344 119175
rect 177184 119113 177344 119147
rect 177184 119085 177219 119113
rect 177247 119085 177281 119113
rect 177309 119085 177344 119113
rect 177184 119051 177344 119085
rect 177184 119023 177219 119051
rect 177247 119023 177281 119051
rect 177309 119023 177344 119051
rect 177184 118989 177344 119023
rect 177184 118961 177219 118989
rect 177247 118961 177281 118989
rect 177309 118961 177344 118989
rect 177184 118944 177344 118961
rect 187029 119175 187339 127961
rect 187029 119147 187077 119175
rect 187105 119147 187139 119175
rect 187167 119147 187201 119175
rect 187229 119147 187263 119175
rect 187291 119147 187339 119175
rect 187029 119113 187339 119147
rect 187029 119085 187077 119113
rect 187105 119085 187139 119113
rect 187167 119085 187201 119113
rect 187229 119085 187263 119113
rect 187291 119085 187339 119113
rect 187029 119051 187339 119085
rect 187029 119023 187077 119051
rect 187105 119023 187139 119051
rect 187167 119023 187201 119051
rect 187229 119023 187263 119051
rect 187291 119023 187339 119051
rect 187029 118989 187339 119023
rect 187029 118961 187077 118989
rect 187105 118961 187139 118989
rect 187167 118961 187201 118989
rect 187229 118961 187263 118989
rect 187291 118961 187339 118989
rect 173529 113147 173577 113175
rect 173605 113147 173639 113175
rect 173667 113147 173701 113175
rect 173729 113147 173763 113175
rect 173791 113147 173839 113175
rect 173529 113113 173839 113147
rect 173529 113085 173577 113113
rect 173605 113085 173639 113113
rect 173667 113085 173701 113113
rect 173729 113085 173763 113113
rect 173791 113085 173839 113113
rect 173529 113051 173839 113085
rect 173529 113023 173577 113051
rect 173605 113023 173639 113051
rect 173667 113023 173701 113051
rect 173729 113023 173763 113051
rect 173791 113023 173839 113051
rect 173529 112989 173839 113023
rect 173529 112961 173577 112989
rect 173605 112961 173639 112989
rect 173667 112961 173701 112989
rect 173729 112961 173763 112989
rect 173791 112961 173839 112989
rect 173529 104175 173839 112961
rect 184864 113175 185024 113192
rect 184864 113147 184899 113175
rect 184927 113147 184961 113175
rect 184989 113147 185024 113175
rect 184864 113113 185024 113147
rect 184864 113085 184899 113113
rect 184927 113085 184961 113113
rect 184989 113085 185024 113113
rect 184864 113051 185024 113085
rect 184864 113023 184899 113051
rect 184927 113023 184961 113051
rect 184989 113023 185024 113051
rect 184864 112989 185024 113023
rect 184864 112961 184899 112989
rect 184927 112961 184961 112989
rect 184989 112961 185024 112989
rect 184864 112944 185024 112961
rect 177184 110175 177344 110192
rect 177184 110147 177219 110175
rect 177247 110147 177281 110175
rect 177309 110147 177344 110175
rect 177184 110113 177344 110147
rect 177184 110085 177219 110113
rect 177247 110085 177281 110113
rect 177309 110085 177344 110113
rect 177184 110051 177344 110085
rect 177184 110023 177219 110051
rect 177247 110023 177281 110051
rect 177309 110023 177344 110051
rect 177184 109989 177344 110023
rect 177184 109961 177219 109989
rect 177247 109961 177281 109989
rect 177309 109961 177344 109989
rect 177184 109944 177344 109961
rect 187029 110175 187339 118961
rect 187029 110147 187077 110175
rect 187105 110147 187139 110175
rect 187167 110147 187201 110175
rect 187229 110147 187263 110175
rect 187291 110147 187339 110175
rect 187029 110113 187339 110147
rect 187029 110085 187077 110113
rect 187105 110085 187139 110113
rect 187167 110085 187201 110113
rect 187229 110085 187263 110113
rect 187291 110085 187339 110113
rect 187029 110051 187339 110085
rect 187029 110023 187077 110051
rect 187105 110023 187139 110051
rect 187167 110023 187201 110051
rect 187229 110023 187263 110051
rect 187291 110023 187339 110051
rect 187029 109989 187339 110023
rect 187029 109961 187077 109989
rect 187105 109961 187139 109989
rect 187167 109961 187201 109989
rect 187229 109961 187263 109989
rect 187291 109961 187339 109989
rect 173529 104147 173577 104175
rect 173605 104147 173639 104175
rect 173667 104147 173701 104175
rect 173729 104147 173763 104175
rect 173791 104147 173839 104175
rect 173529 104113 173839 104147
rect 173529 104085 173577 104113
rect 173605 104085 173639 104113
rect 173667 104085 173701 104113
rect 173729 104085 173763 104113
rect 173791 104085 173839 104113
rect 173529 104051 173839 104085
rect 173529 104023 173577 104051
rect 173605 104023 173639 104051
rect 173667 104023 173701 104051
rect 173729 104023 173763 104051
rect 173791 104023 173839 104051
rect 173529 103989 173839 104023
rect 173529 103961 173577 103989
rect 173605 103961 173639 103989
rect 173667 103961 173701 103989
rect 173729 103961 173763 103989
rect 173791 103961 173839 103989
rect 173529 95175 173839 103961
rect 184864 104175 185024 104192
rect 184864 104147 184899 104175
rect 184927 104147 184961 104175
rect 184989 104147 185024 104175
rect 184864 104113 185024 104147
rect 184864 104085 184899 104113
rect 184927 104085 184961 104113
rect 184989 104085 185024 104113
rect 184864 104051 185024 104085
rect 184864 104023 184899 104051
rect 184927 104023 184961 104051
rect 184989 104023 185024 104051
rect 184864 103989 185024 104023
rect 184864 103961 184899 103989
rect 184927 103961 184961 103989
rect 184989 103961 185024 103989
rect 184864 103944 185024 103961
rect 177184 101175 177344 101192
rect 177184 101147 177219 101175
rect 177247 101147 177281 101175
rect 177309 101147 177344 101175
rect 177184 101113 177344 101147
rect 177184 101085 177219 101113
rect 177247 101085 177281 101113
rect 177309 101085 177344 101113
rect 177184 101051 177344 101085
rect 177184 101023 177219 101051
rect 177247 101023 177281 101051
rect 177309 101023 177344 101051
rect 177184 100989 177344 101023
rect 177184 100961 177219 100989
rect 177247 100961 177281 100989
rect 177309 100961 177344 100989
rect 177184 100944 177344 100961
rect 187029 101175 187339 109961
rect 187029 101147 187077 101175
rect 187105 101147 187139 101175
rect 187167 101147 187201 101175
rect 187229 101147 187263 101175
rect 187291 101147 187339 101175
rect 187029 101113 187339 101147
rect 187029 101085 187077 101113
rect 187105 101085 187139 101113
rect 187167 101085 187201 101113
rect 187229 101085 187263 101113
rect 187291 101085 187339 101113
rect 187029 101051 187339 101085
rect 187029 101023 187077 101051
rect 187105 101023 187139 101051
rect 187167 101023 187201 101051
rect 187229 101023 187263 101051
rect 187291 101023 187339 101051
rect 187029 100989 187339 101023
rect 187029 100961 187077 100989
rect 187105 100961 187139 100989
rect 187167 100961 187201 100989
rect 187229 100961 187263 100989
rect 187291 100961 187339 100989
rect 173529 95147 173577 95175
rect 173605 95147 173639 95175
rect 173667 95147 173701 95175
rect 173729 95147 173763 95175
rect 173791 95147 173839 95175
rect 173529 95113 173839 95147
rect 173529 95085 173577 95113
rect 173605 95085 173639 95113
rect 173667 95085 173701 95113
rect 173729 95085 173763 95113
rect 173791 95085 173839 95113
rect 173529 95051 173839 95085
rect 173529 95023 173577 95051
rect 173605 95023 173639 95051
rect 173667 95023 173701 95051
rect 173729 95023 173763 95051
rect 173791 95023 173839 95051
rect 173529 94989 173839 95023
rect 173529 94961 173577 94989
rect 173605 94961 173639 94989
rect 173667 94961 173701 94989
rect 173729 94961 173763 94989
rect 173791 94961 173839 94989
rect 173529 86175 173839 94961
rect 184864 95175 185024 95192
rect 184864 95147 184899 95175
rect 184927 95147 184961 95175
rect 184989 95147 185024 95175
rect 184864 95113 185024 95147
rect 184864 95085 184899 95113
rect 184927 95085 184961 95113
rect 184989 95085 185024 95113
rect 184864 95051 185024 95085
rect 184864 95023 184899 95051
rect 184927 95023 184961 95051
rect 184989 95023 185024 95051
rect 184864 94989 185024 95023
rect 184864 94961 184899 94989
rect 184927 94961 184961 94989
rect 184989 94961 185024 94989
rect 184864 94944 185024 94961
rect 177184 92175 177344 92192
rect 177184 92147 177219 92175
rect 177247 92147 177281 92175
rect 177309 92147 177344 92175
rect 177184 92113 177344 92147
rect 177184 92085 177219 92113
rect 177247 92085 177281 92113
rect 177309 92085 177344 92113
rect 177184 92051 177344 92085
rect 177184 92023 177219 92051
rect 177247 92023 177281 92051
rect 177309 92023 177344 92051
rect 177184 91989 177344 92023
rect 177184 91961 177219 91989
rect 177247 91961 177281 91989
rect 177309 91961 177344 91989
rect 177184 91944 177344 91961
rect 187029 92175 187339 100961
rect 187029 92147 187077 92175
rect 187105 92147 187139 92175
rect 187167 92147 187201 92175
rect 187229 92147 187263 92175
rect 187291 92147 187339 92175
rect 187029 92113 187339 92147
rect 187029 92085 187077 92113
rect 187105 92085 187139 92113
rect 187167 92085 187201 92113
rect 187229 92085 187263 92113
rect 187291 92085 187339 92113
rect 187029 92051 187339 92085
rect 187029 92023 187077 92051
rect 187105 92023 187139 92051
rect 187167 92023 187201 92051
rect 187229 92023 187263 92051
rect 187291 92023 187339 92051
rect 187029 91989 187339 92023
rect 187029 91961 187077 91989
rect 187105 91961 187139 91989
rect 187167 91961 187201 91989
rect 187229 91961 187263 91989
rect 187291 91961 187339 91989
rect 173529 86147 173577 86175
rect 173605 86147 173639 86175
rect 173667 86147 173701 86175
rect 173729 86147 173763 86175
rect 173791 86147 173839 86175
rect 173529 86113 173839 86147
rect 173529 86085 173577 86113
rect 173605 86085 173639 86113
rect 173667 86085 173701 86113
rect 173729 86085 173763 86113
rect 173791 86085 173839 86113
rect 173529 86051 173839 86085
rect 173529 86023 173577 86051
rect 173605 86023 173639 86051
rect 173667 86023 173701 86051
rect 173729 86023 173763 86051
rect 173791 86023 173839 86051
rect 173529 85989 173839 86023
rect 173529 85961 173577 85989
rect 173605 85961 173639 85989
rect 173667 85961 173701 85989
rect 173729 85961 173763 85989
rect 173791 85961 173839 85989
rect 173529 77175 173839 85961
rect 184864 86175 185024 86192
rect 184864 86147 184899 86175
rect 184927 86147 184961 86175
rect 184989 86147 185024 86175
rect 184864 86113 185024 86147
rect 184864 86085 184899 86113
rect 184927 86085 184961 86113
rect 184989 86085 185024 86113
rect 184864 86051 185024 86085
rect 184864 86023 184899 86051
rect 184927 86023 184961 86051
rect 184989 86023 185024 86051
rect 184864 85989 185024 86023
rect 184864 85961 184899 85989
rect 184927 85961 184961 85989
rect 184989 85961 185024 85989
rect 184864 85944 185024 85961
rect 177184 83175 177344 83192
rect 177184 83147 177219 83175
rect 177247 83147 177281 83175
rect 177309 83147 177344 83175
rect 177184 83113 177344 83147
rect 177184 83085 177219 83113
rect 177247 83085 177281 83113
rect 177309 83085 177344 83113
rect 177184 83051 177344 83085
rect 177184 83023 177219 83051
rect 177247 83023 177281 83051
rect 177309 83023 177344 83051
rect 177184 82989 177344 83023
rect 177184 82961 177219 82989
rect 177247 82961 177281 82989
rect 177309 82961 177344 82989
rect 177184 82944 177344 82961
rect 187029 83175 187339 91961
rect 187029 83147 187077 83175
rect 187105 83147 187139 83175
rect 187167 83147 187201 83175
rect 187229 83147 187263 83175
rect 187291 83147 187339 83175
rect 187029 83113 187339 83147
rect 187029 83085 187077 83113
rect 187105 83085 187139 83113
rect 187167 83085 187201 83113
rect 187229 83085 187263 83113
rect 187291 83085 187339 83113
rect 187029 83051 187339 83085
rect 187029 83023 187077 83051
rect 187105 83023 187139 83051
rect 187167 83023 187201 83051
rect 187229 83023 187263 83051
rect 187291 83023 187339 83051
rect 187029 82989 187339 83023
rect 187029 82961 187077 82989
rect 187105 82961 187139 82989
rect 187167 82961 187201 82989
rect 187229 82961 187263 82989
rect 187291 82961 187339 82989
rect 173529 77147 173577 77175
rect 173605 77147 173639 77175
rect 173667 77147 173701 77175
rect 173729 77147 173763 77175
rect 173791 77147 173839 77175
rect 173529 77113 173839 77147
rect 173529 77085 173577 77113
rect 173605 77085 173639 77113
rect 173667 77085 173701 77113
rect 173729 77085 173763 77113
rect 173791 77085 173839 77113
rect 173529 77051 173839 77085
rect 173529 77023 173577 77051
rect 173605 77023 173639 77051
rect 173667 77023 173701 77051
rect 173729 77023 173763 77051
rect 173791 77023 173839 77051
rect 173529 76989 173839 77023
rect 173529 76961 173577 76989
rect 173605 76961 173639 76989
rect 173667 76961 173701 76989
rect 173729 76961 173763 76989
rect 173791 76961 173839 76989
rect 173529 68175 173839 76961
rect 184864 77175 185024 77192
rect 184864 77147 184899 77175
rect 184927 77147 184961 77175
rect 184989 77147 185024 77175
rect 184864 77113 185024 77147
rect 184864 77085 184899 77113
rect 184927 77085 184961 77113
rect 184989 77085 185024 77113
rect 184864 77051 185024 77085
rect 184864 77023 184899 77051
rect 184927 77023 184961 77051
rect 184989 77023 185024 77051
rect 184864 76989 185024 77023
rect 184864 76961 184899 76989
rect 184927 76961 184961 76989
rect 184989 76961 185024 76989
rect 184864 76944 185024 76961
rect 177184 74175 177344 74192
rect 177184 74147 177219 74175
rect 177247 74147 177281 74175
rect 177309 74147 177344 74175
rect 177184 74113 177344 74147
rect 177184 74085 177219 74113
rect 177247 74085 177281 74113
rect 177309 74085 177344 74113
rect 177184 74051 177344 74085
rect 177184 74023 177219 74051
rect 177247 74023 177281 74051
rect 177309 74023 177344 74051
rect 177184 73989 177344 74023
rect 177184 73961 177219 73989
rect 177247 73961 177281 73989
rect 177309 73961 177344 73989
rect 177184 73944 177344 73961
rect 187029 74175 187339 82961
rect 187029 74147 187077 74175
rect 187105 74147 187139 74175
rect 187167 74147 187201 74175
rect 187229 74147 187263 74175
rect 187291 74147 187339 74175
rect 187029 74113 187339 74147
rect 187029 74085 187077 74113
rect 187105 74085 187139 74113
rect 187167 74085 187201 74113
rect 187229 74085 187263 74113
rect 187291 74085 187339 74113
rect 187029 74051 187339 74085
rect 187029 74023 187077 74051
rect 187105 74023 187139 74051
rect 187167 74023 187201 74051
rect 187229 74023 187263 74051
rect 187291 74023 187339 74051
rect 187029 73989 187339 74023
rect 187029 73961 187077 73989
rect 187105 73961 187139 73989
rect 187167 73961 187201 73989
rect 187229 73961 187263 73989
rect 187291 73961 187339 73989
rect 173529 68147 173577 68175
rect 173605 68147 173639 68175
rect 173667 68147 173701 68175
rect 173729 68147 173763 68175
rect 173791 68147 173839 68175
rect 173529 68113 173839 68147
rect 173529 68085 173577 68113
rect 173605 68085 173639 68113
rect 173667 68085 173701 68113
rect 173729 68085 173763 68113
rect 173791 68085 173839 68113
rect 173529 68051 173839 68085
rect 173529 68023 173577 68051
rect 173605 68023 173639 68051
rect 173667 68023 173701 68051
rect 173729 68023 173763 68051
rect 173791 68023 173839 68051
rect 173529 67989 173839 68023
rect 173529 67961 173577 67989
rect 173605 67961 173639 67989
rect 173667 67961 173701 67989
rect 173729 67961 173763 67989
rect 173791 67961 173839 67989
rect 173529 59175 173839 67961
rect 184864 68175 185024 68192
rect 184864 68147 184899 68175
rect 184927 68147 184961 68175
rect 184989 68147 185024 68175
rect 184864 68113 185024 68147
rect 184864 68085 184899 68113
rect 184927 68085 184961 68113
rect 184989 68085 185024 68113
rect 184864 68051 185024 68085
rect 184864 68023 184899 68051
rect 184927 68023 184961 68051
rect 184989 68023 185024 68051
rect 184864 67989 185024 68023
rect 184864 67961 184899 67989
rect 184927 67961 184961 67989
rect 184989 67961 185024 67989
rect 184864 67944 185024 67961
rect 177184 65175 177344 65192
rect 177184 65147 177219 65175
rect 177247 65147 177281 65175
rect 177309 65147 177344 65175
rect 177184 65113 177344 65147
rect 177184 65085 177219 65113
rect 177247 65085 177281 65113
rect 177309 65085 177344 65113
rect 177184 65051 177344 65085
rect 177184 65023 177219 65051
rect 177247 65023 177281 65051
rect 177309 65023 177344 65051
rect 177184 64989 177344 65023
rect 177184 64961 177219 64989
rect 177247 64961 177281 64989
rect 177309 64961 177344 64989
rect 177184 64944 177344 64961
rect 187029 65175 187339 73961
rect 187029 65147 187077 65175
rect 187105 65147 187139 65175
rect 187167 65147 187201 65175
rect 187229 65147 187263 65175
rect 187291 65147 187339 65175
rect 187029 65113 187339 65147
rect 187029 65085 187077 65113
rect 187105 65085 187139 65113
rect 187167 65085 187201 65113
rect 187229 65085 187263 65113
rect 187291 65085 187339 65113
rect 187029 65051 187339 65085
rect 187029 65023 187077 65051
rect 187105 65023 187139 65051
rect 187167 65023 187201 65051
rect 187229 65023 187263 65051
rect 187291 65023 187339 65051
rect 187029 64989 187339 65023
rect 187029 64961 187077 64989
rect 187105 64961 187139 64989
rect 187167 64961 187201 64989
rect 187229 64961 187263 64989
rect 187291 64961 187339 64989
rect 173529 59147 173577 59175
rect 173605 59147 173639 59175
rect 173667 59147 173701 59175
rect 173729 59147 173763 59175
rect 173791 59147 173839 59175
rect 173529 59113 173839 59147
rect 173529 59085 173577 59113
rect 173605 59085 173639 59113
rect 173667 59085 173701 59113
rect 173729 59085 173763 59113
rect 173791 59085 173839 59113
rect 173529 59051 173839 59085
rect 173529 59023 173577 59051
rect 173605 59023 173639 59051
rect 173667 59023 173701 59051
rect 173729 59023 173763 59051
rect 173791 59023 173839 59051
rect 173529 58989 173839 59023
rect 173529 58961 173577 58989
rect 173605 58961 173639 58989
rect 173667 58961 173701 58989
rect 173729 58961 173763 58989
rect 173791 58961 173839 58989
rect 173529 50175 173839 58961
rect 184864 59175 185024 59192
rect 184864 59147 184899 59175
rect 184927 59147 184961 59175
rect 184989 59147 185024 59175
rect 184864 59113 185024 59147
rect 184864 59085 184899 59113
rect 184927 59085 184961 59113
rect 184989 59085 185024 59113
rect 184864 59051 185024 59085
rect 184864 59023 184899 59051
rect 184927 59023 184961 59051
rect 184989 59023 185024 59051
rect 184864 58989 185024 59023
rect 184864 58961 184899 58989
rect 184927 58961 184961 58989
rect 184989 58961 185024 58989
rect 184864 58944 185024 58961
rect 177184 56175 177344 56192
rect 177184 56147 177219 56175
rect 177247 56147 177281 56175
rect 177309 56147 177344 56175
rect 177184 56113 177344 56147
rect 177184 56085 177219 56113
rect 177247 56085 177281 56113
rect 177309 56085 177344 56113
rect 177184 56051 177344 56085
rect 177184 56023 177219 56051
rect 177247 56023 177281 56051
rect 177309 56023 177344 56051
rect 177184 55989 177344 56023
rect 177184 55961 177219 55989
rect 177247 55961 177281 55989
rect 177309 55961 177344 55989
rect 177184 55944 177344 55961
rect 187029 56175 187339 64961
rect 187029 56147 187077 56175
rect 187105 56147 187139 56175
rect 187167 56147 187201 56175
rect 187229 56147 187263 56175
rect 187291 56147 187339 56175
rect 187029 56113 187339 56147
rect 187029 56085 187077 56113
rect 187105 56085 187139 56113
rect 187167 56085 187201 56113
rect 187229 56085 187263 56113
rect 187291 56085 187339 56113
rect 187029 56051 187339 56085
rect 187029 56023 187077 56051
rect 187105 56023 187139 56051
rect 187167 56023 187201 56051
rect 187229 56023 187263 56051
rect 187291 56023 187339 56051
rect 187029 55989 187339 56023
rect 187029 55961 187077 55989
rect 187105 55961 187139 55989
rect 187167 55961 187201 55989
rect 187229 55961 187263 55989
rect 187291 55961 187339 55989
rect 173529 50147 173577 50175
rect 173605 50147 173639 50175
rect 173667 50147 173701 50175
rect 173729 50147 173763 50175
rect 173791 50147 173839 50175
rect 173529 50113 173839 50147
rect 173529 50085 173577 50113
rect 173605 50085 173639 50113
rect 173667 50085 173701 50113
rect 173729 50085 173763 50113
rect 173791 50085 173839 50113
rect 173529 50051 173839 50085
rect 173529 50023 173577 50051
rect 173605 50023 173639 50051
rect 173667 50023 173701 50051
rect 173729 50023 173763 50051
rect 173791 50023 173839 50051
rect 173529 49989 173839 50023
rect 173529 49961 173577 49989
rect 173605 49961 173639 49989
rect 173667 49961 173701 49989
rect 173729 49961 173763 49989
rect 173791 49961 173839 49989
rect 173529 41175 173839 49961
rect 184864 50175 185024 50192
rect 184864 50147 184899 50175
rect 184927 50147 184961 50175
rect 184989 50147 185024 50175
rect 184864 50113 185024 50147
rect 184864 50085 184899 50113
rect 184927 50085 184961 50113
rect 184989 50085 185024 50113
rect 184864 50051 185024 50085
rect 184864 50023 184899 50051
rect 184927 50023 184961 50051
rect 184989 50023 185024 50051
rect 184864 49989 185024 50023
rect 184864 49961 184899 49989
rect 184927 49961 184961 49989
rect 184989 49961 185024 49989
rect 184864 49944 185024 49961
rect 177184 47175 177344 47192
rect 177184 47147 177219 47175
rect 177247 47147 177281 47175
rect 177309 47147 177344 47175
rect 177184 47113 177344 47147
rect 177184 47085 177219 47113
rect 177247 47085 177281 47113
rect 177309 47085 177344 47113
rect 177184 47051 177344 47085
rect 177184 47023 177219 47051
rect 177247 47023 177281 47051
rect 177309 47023 177344 47051
rect 177184 46989 177344 47023
rect 177184 46961 177219 46989
rect 177247 46961 177281 46989
rect 177309 46961 177344 46989
rect 177184 46944 177344 46961
rect 187029 47175 187339 55961
rect 187029 47147 187077 47175
rect 187105 47147 187139 47175
rect 187167 47147 187201 47175
rect 187229 47147 187263 47175
rect 187291 47147 187339 47175
rect 187029 47113 187339 47147
rect 187029 47085 187077 47113
rect 187105 47085 187139 47113
rect 187167 47085 187201 47113
rect 187229 47085 187263 47113
rect 187291 47085 187339 47113
rect 187029 47051 187339 47085
rect 187029 47023 187077 47051
rect 187105 47023 187139 47051
rect 187167 47023 187201 47051
rect 187229 47023 187263 47051
rect 187291 47023 187339 47051
rect 187029 46989 187339 47023
rect 187029 46961 187077 46989
rect 187105 46961 187139 46989
rect 187167 46961 187201 46989
rect 187229 46961 187263 46989
rect 187291 46961 187339 46989
rect 173529 41147 173577 41175
rect 173605 41147 173639 41175
rect 173667 41147 173701 41175
rect 173729 41147 173763 41175
rect 173791 41147 173839 41175
rect 173529 41113 173839 41147
rect 173529 41085 173577 41113
rect 173605 41085 173639 41113
rect 173667 41085 173701 41113
rect 173729 41085 173763 41113
rect 173791 41085 173839 41113
rect 173529 41051 173839 41085
rect 173529 41023 173577 41051
rect 173605 41023 173639 41051
rect 173667 41023 173701 41051
rect 173729 41023 173763 41051
rect 173791 41023 173839 41051
rect 173529 40989 173839 41023
rect 173529 40961 173577 40989
rect 173605 40961 173639 40989
rect 173667 40961 173701 40989
rect 173729 40961 173763 40989
rect 173791 40961 173839 40989
rect 173529 32175 173839 40961
rect 184864 41175 185024 41192
rect 184864 41147 184899 41175
rect 184927 41147 184961 41175
rect 184989 41147 185024 41175
rect 184864 41113 185024 41147
rect 184864 41085 184899 41113
rect 184927 41085 184961 41113
rect 184989 41085 185024 41113
rect 184864 41051 185024 41085
rect 184864 41023 184899 41051
rect 184927 41023 184961 41051
rect 184989 41023 185024 41051
rect 184864 40989 185024 41023
rect 184864 40961 184899 40989
rect 184927 40961 184961 40989
rect 184989 40961 185024 40989
rect 184864 40944 185024 40961
rect 177184 38175 177344 38192
rect 177184 38147 177219 38175
rect 177247 38147 177281 38175
rect 177309 38147 177344 38175
rect 177184 38113 177344 38147
rect 177184 38085 177219 38113
rect 177247 38085 177281 38113
rect 177309 38085 177344 38113
rect 177184 38051 177344 38085
rect 177184 38023 177219 38051
rect 177247 38023 177281 38051
rect 177309 38023 177344 38051
rect 177184 37989 177344 38023
rect 177184 37961 177219 37989
rect 177247 37961 177281 37989
rect 177309 37961 177344 37989
rect 177184 37944 177344 37961
rect 187029 38175 187339 46961
rect 187029 38147 187077 38175
rect 187105 38147 187139 38175
rect 187167 38147 187201 38175
rect 187229 38147 187263 38175
rect 187291 38147 187339 38175
rect 187029 38113 187339 38147
rect 187029 38085 187077 38113
rect 187105 38085 187139 38113
rect 187167 38085 187201 38113
rect 187229 38085 187263 38113
rect 187291 38085 187339 38113
rect 187029 38051 187339 38085
rect 187029 38023 187077 38051
rect 187105 38023 187139 38051
rect 187167 38023 187201 38051
rect 187229 38023 187263 38051
rect 187291 38023 187339 38051
rect 187029 37989 187339 38023
rect 187029 37961 187077 37989
rect 187105 37961 187139 37989
rect 187167 37961 187201 37989
rect 187229 37961 187263 37989
rect 187291 37961 187339 37989
rect 173529 32147 173577 32175
rect 173605 32147 173639 32175
rect 173667 32147 173701 32175
rect 173729 32147 173763 32175
rect 173791 32147 173839 32175
rect 173529 32113 173839 32147
rect 173529 32085 173577 32113
rect 173605 32085 173639 32113
rect 173667 32085 173701 32113
rect 173729 32085 173763 32113
rect 173791 32085 173839 32113
rect 173529 32051 173839 32085
rect 173529 32023 173577 32051
rect 173605 32023 173639 32051
rect 173667 32023 173701 32051
rect 173729 32023 173763 32051
rect 173791 32023 173839 32051
rect 173529 31989 173839 32023
rect 173529 31961 173577 31989
rect 173605 31961 173639 31989
rect 173667 31961 173701 31989
rect 173729 31961 173763 31989
rect 173791 31961 173839 31989
rect 173529 23175 173839 31961
rect 184864 32175 185024 32192
rect 184864 32147 184899 32175
rect 184927 32147 184961 32175
rect 184989 32147 185024 32175
rect 184864 32113 185024 32147
rect 184864 32085 184899 32113
rect 184927 32085 184961 32113
rect 184989 32085 185024 32113
rect 184864 32051 185024 32085
rect 184864 32023 184899 32051
rect 184927 32023 184961 32051
rect 184989 32023 185024 32051
rect 184864 31989 185024 32023
rect 184864 31961 184899 31989
rect 184927 31961 184961 31989
rect 184989 31961 185024 31989
rect 184864 31944 185024 31961
rect 177184 29175 177344 29192
rect 177184 29147 177219 29175
rect 177247 29147 177281 29175
rect 177309 29147 177344 29175
rect 177184 29113 177344 29147
rect 177184 29085 177219 29113
rect 177247 29085 177281 29113
rect 177309 29085 177344 29113
rect 177184 29051 177344 29085
rect 177184 29023 177219 29051
rect 177247 29023 177281 29051
rect 177309 29023 177344 29051
rect 177184 28989 177344 29023
rect 177184 28961 177219 28989
rect 177247 28961 177281 28989
rect 177309 28961 177344 28989
rect 177184 28944 177344 28961
rect 187029 29175 187339 37961
rect 187029 29147 187077 29175
rect 187105 29147 187139 29175
rect 187167 29147 187201 29175
rect 187229 29147 187263 29175
rect 187291 29147 187339 29175
rect 187029 29113 187339 29147
rect 187029 29085 187077 29113
rect 187105 29085 187139 29113
rect 187167 29085 187201 29113
rect 187229 29085 187263 29113
rect 187291 29085 187339 29113
rect 187029 29051 187339 29085
rect 187029 29023 187077 29051
rect 187105 29023 187139 29051
rect 187167 29023 187201 29051
rect 187229 29023 187263 29051
rect 187291 29023 187339 29051
rect 187029 28989 187339 29023
rect 187029 28961 187077 28989
rect 187105 28961 187139 28989
rect 187167 28961 187201 28989
rect 187229 28961 187263 28989
rect 187291 28961 187339 28989
rect 173529 23147 173577 23175
rect 173605 23147 173639 23175
rect 173667 23147 173701 23175
rect 173729 23147 173763 23175
rect 173791 23147 173839 23175
rect 173529 23113 173839 23147
rect 173529 23085 173577 23113
rect 173605 23085 173639 23113
rect 173667 23085 173701 23113
rect 173729 23085 173763 23113
rect 173791 23085 173839 23113
rect 173529 23051 173839 23085
rect 173529 23023 173577 23051
rect 173605 23023 173639 23051
rect 173667 23023 173701 23051
rect 173729 23023 173763 23051
rect 173791 23023 173839 23051
rect 173529 22989 173839 23023
rect 173529 22961 173577 22989
rect 173605 22961 173639 22989
rect 173667 22961 173701 22989
rect 173729 22961 173763 22989
rect 173791 22961 173839 22989
rect 173529 14175 173839 22961
rect 184864 23175 185024 23192
rect 184864 23147 184899 23175
rect 184927 23147 184961 23175
rect 184989 23147 185024 23175
rect 184864 23113 185024 23147
rect 184864 23085 184899 23113
rect 184927 23085 184961 23113
rect 184989 23085 185024 23113
rect 184864 23051 185024 23085
rect 184864 23023 184899 23051
rect 184927 23023 184961 23051
rect 184989 23023 185024 23051
rect 184864 22989 185024 23023
rect 184864 22961 184899 22989
rect 184927 22961 184961 22989
rect 184989 22961 185024 22989
rect 184864 22944 185024 22961
rect 177184 20175 177344 20192
rect 177184 20147 177219 20175
rect 177247 20147 177281 20175
rect 177309 20147 177344 20175
rect 177184 20113 177344 20147
rect 177184 20085 177219 20113
rect 177247 20085 177281 20113
rect 177309 20085 177344 20113
rect 177184 20051 177344 20085
rect 177184 20023 177219 20051
rect 177247 20023 177281 20051
rect 177309 20023 177344 20051
rect 177184 19989 177344 20023
rect 177184 19961 177219 19989
rect 177247 19961 177281 19989
rect 177309 19961 177344 19989
rect 177184 19944 177344 19961
rect 187029 20175 187339 28961
rect 187029 20147 187077 20175
rect 187105 20147 187139 20175
rect 187167 20147 187201 20175
rect 187229 20147 187263 20175
rect 187291 20147 187339 20175
rect 187029 20113 187339 20147
rect 187029 20085 187077 20113
rect 187105 20085 187139 20113
rect 187167 20085 187201 20113
rect 187229 20085 187263 20113
rect 187291 20085 187339 20113
rect 187029 20051 187339 20085
rect 187029 20023 187077 20051
rect 187105 20023 187139 20051
rect 187167 20023 187201 20051
rect 187229 20023 187263 20051
rect 187291 20023 187339 20051
rect 187029 19989 187339 20023
rect 187029 19961 187077 19989
rect 187105 19961 187139 19989
rect 187167 19961 187201 19989
rect 187229 19961 187263 19989
rect 187291 19961 187339 19989
rect 173529 14147 173577 14175
rect 173605 14147 173639 14175
rect 173667 14147 173701 14175
rect 173729 14147 173763 14175
rect 173791 14147 173839 14175
rect 173529 14113 173839 14147
rect 173529 14085 173577 14113
rect 173605 14085 173639 14113
rect 173667 14085 173701 14113
rect 173729 14085 173763 14113
rect 173791 14085 173839 14113
rect 173529 14051 173839 14085
rect 173529 14023 173577 14051
rect 173605 14023 173639 14051
rect 173667 14023 173701 14051
rect 173729 14023 173763 14051
rect 173791 14023 173839 14051
rect 173529 13989 173839 14023
rect 173529 13961 173577 13989
rect 173605 13961 173639 13989
rect 173667 13961 173701 13989
rect 173729 13961 173763 13989
rect 173791 13961 173839 13989
rect 173529 5175 173839 13961
rect 184864 14175 185024 14192
rect 184864 14147 184899 14175
rect 184927 14147 184961 14175
rect 184989 14147 185024 14175
rect 184864 14113 185024 14147
rect 184864 14085 184899 14113
rect 184927 14085 184961 14113
rect 184989 14085 185024 14113
rect 184864 14051 185024 14085
rect 184864 14023 184899 14051
rect 184927 14023 184961 14051
rect 184989 14023 185024 14051
rect 184864 13989 185024 14023
rect 184864 13961 184899 13989
rect 184927 13961 184961 13989
rect 184989 13961 185024 13989
rect 184864 13944 185024 13961
rect 177184 11175 177344 11192
rect 177184 11147 177219 11175
rect 177247 11147 177281 11175
rect 177309 11147 177344 11175
rect 177184 11113 177344 11147
rect 177184 11085 177219 11113
rect 177247 11085 177281 11113
rect 177309 11085 177344 11113
rect 177184 11051 177344 11085
rect 177184 11023 177219 11051
rect 177247 11023 177281 11051
rect 177309 11023 177344 11051
rect 177184 10989 177344 11023
rect 177184 10961 177219 10989
rect 177247 10961 177281 10989
rect 177309 10961 177344 10989
rect 177184 10944 177344 10961
rect 187029 11175 187339 19961
rect 187029 11147 187077 11175
rect 187105 11147 187139 11175
rect 187167 11147 187201 11175
rect 187229 11147 187263 11175
rect 187291 11147 187339 11175
rect 187029 11113 187339 11147
rect 187029 11085 187077 11113
rect 187105 11085 187139 11113
rect 187167 11085 187201 11113
rect 187229 11085 187263 11113
rect 187291 11085 187339 11113
rect 187029 11051 187339 11085
rect 187029 11023 187077 11051
rect 187105 11023 187139 11051
rect 187167 11023 187201 11051
rect 187229 11023 187263 11051
rect 187291 11023 187339 11051
rect 187029 10989 187339 11023
rect 187029 10961 187077 10989
rect 187105 10961 187139 10989
rect 187167 10961 187201 10989
rect 187229 10961 187263 10989
rect 187291 10961 187339 10989
rect 173529 5147 173577 5175
rect 173605 5147 173639 5175
rect 173667 5147 173701 5175
rect 173729 5147 173763 5175
rect 173791 5147 173839 5175
rect 173529 5113 173839 5147
rect 173529 5085 173577 5113
rect 173605 5085 173639 5113
rect 173667 5085 173701 5113
rect 173729 5085 173763 5113
rect 173791 5085 173839 5113
rect 173529 5051 173839 5085
rect 173529 5023 173577 5051
rect 173605 5023 173639 5051
rect 173667 5023 173701 5051
rect 173729 5023 173763 5051
rect 173791 5023 173839 5051
rect 173529 4989 173839 5023
rect 173529 4961 173577 4989
rect 173605 4961 173639 4989
rect 173667 4961 173701 4989
rect 173729 4961 173763 4989
rect 173791 4961 173839 4989
rect 173529 -560 173839 4961
rect 184864 5175 185024 5192
rect 184864 5147 184899 5175
rect 184927 5147 184961 5175
rect 184989 5147 185024 5175
rect 184864 5113 185024 5147
rect 184864 5085 184899 5113
rect 184927 5085 184961 5113
rect 184989 5085 185024 5113
rect 184864 5051 185024 5085
rect 184864 5023 184899 5051
rect 184927 5023 184961 5051
rect 184989 5023 185024 5051
rect 184864 4989 185024 5023
rect 184864 4961 184899 4989
rect 184927 4961 184961 4989
rect 184989 4961 185024 4989
rect 184864 4944 185024 4961
rect 173529 -588 173577 -560
rect 173605 -588 173639 -560
rect 173667 -588 173701 -560
rect 173729 -588 173763 -560
rect 173791 -588 173839 -560
rect 173529 -622 173839 -588
rect 173529 -650 173577 -622
rect 173605 -650 173639 -622
rect 173667 -650 173701 -622
rect 173729 -650 173763 -622
rect 173791 -650 173839 -622
rect 173529 -684 173839 -650
rect 173529 -712 173577 -684
rect 173605 -712 173639 -684
rect 173667 -712 173701 -684
rect 173729 -712 173763 -684
rect 173791 -712 173839 -684
rect 173529 -746 173839 -712
rect 173529 -774 173577 -746
rect 173605 -774 173639 -746
rect 173667 -774 173701 -746
rect 173729 -774 173763 -746
rect 173791 -774 173839 -746
rect 173529 -822 173839 -774
rect 187029 2175 187339 10961
rect 187029 2147 187077 2175
rect 187105 2147 187139 2175
rect 187167 2147 187201 2175
rect 187229 2147 187263 2175
rect 187291 2147 187339 2175
rect 187029 2113 187339 2147
rect 187029 2085 187077 2113
rect 187105 2085 187139 2113
rect 187167 2085 187201 2113
rect 187229 2085 187263 2113
rect 187291 2085 187339 2113
rect 187029 2051 187339 2085
rect 187029 2023 187077 2051
rect 187105 2023 187139 2051
rect 187167 2023 187201 2051
rect 187229 2023 187263 2051
rect 187291 2023 187339 2051
rect 187029 1989 187339 2023
rect 187029 1961 187077 1989
rect 187105 1961 187139 1989
rect 187167 1961 187201 1989
rect 187229 1961 187263 1989
rect 187291 1961 187339 1989
rect 187029 -80 187339 1961
rect 187029 -108 187077 -80
rect 187105 -108 187139 -80
rect 187167 -108 187201 -80
rect 187229 -108 187263 -80
rect 187291 -108 187339 -80
rect 187029 -142 187339 -108
rect 187029 -170 187077 -142
rect 187105 -170 187139 -142
rect 187167 -170 187201 -142
rect 187229 -170 187263 -142
rect 187291 -170 187339 -142
rect 187029 -204 187339 -170
rect 187029 -232 187077 -204
rect 187105 -232 187139 -204
rect 187167 -232 187201 -204
rect 187229 -232 187263 -204
rect 187291 -232 187339 -204
rect 187029 -266 187339 -232
rect 187029 -294 187077 -266
rect 187105 -294 187139 -266
rect 187167 -294 187201 -266
rect 187229 -294 187263 -266
rect 187291 -294 187339 -266
rect 187029 -822 187339 -294
rect 188889 299086 189199 299134
rect 188889 299058 188937 299086
rect 188965 299058 188999 299086
rect 189027 299058 189061 299086
rect 189089 299058 189123 299086
rect 189151 299058 189199 299086
rect 188889 299024 189199 299058
rect 188889 298996 188937 299024
rect 188965 298996 188999 299024
rect 189027 298996 189061 299024
rect 189089 298996 189123 299024
rect 189151 298996 189199 299024
rect 188889 298962 189199 298996
rect 188889 298934 188937 298962
rect 188965 298934 188999 298962
rect 189027 298934 189061 298962
rect 189089 298934 189123 298962
rect 189151 298934 189199 298962
rect 188889 298900 189199 298934
rect 188889 298872 188937 298900
rect 188965 298872 188999 298900
rect 189027 298872 189061 298900
rect 189089 298872 189123 298900
rect 189151 298872 189199 298900
rect 188889 293175 189199 298872
rect 188889 293147 188937 293175
rect 188965 293147 188999 293175
rect 189027 293147 189061 293175
rect 189089 293147 189123 293175
rect 189151 293147 189199 293175
rect 188889 293113 189199 293147
rect 188889 293085 188937 293113
rect 188965 293085 188999 293113
rect 189027 293085 189061 293113
rect 189089 293085 189123 293113
rect 189151 293085 189199 293113
rect 188889 293051 189199 293085
rect 188889 293023 188937 293051
rect 188965 293023 188999 293051
rect 189027 293023 189061 293051
rect 189089 293023 189123 293051
rect 189151 293023 189199 293051
rect 188889 292989 189199 293023
rect 188889 292961 188937 292989
rect 188965 292961 188999 292989
rect 189027 292961 189061 292989
rect 189089 292961 189123 292989
rect 189151 292961 189199 292989
rect 188889 284175 189199 292961
rect 188889 284147 188937 284175
rect 188965 284147 188999 284175
rect 189027 284147 189061 284175
rect 189089 284147 189123 284175
rect 189151 284147 189199 284175
rect 188889 284113 189199 284147
rect 188889 284085 188937 284113
rect 188965 284085 188999 284113
rect 189027 284085 189061 284113
rect 189089 284085 189123 284113
rect 189151 284085 189199 284113
rect 188889 284051 189199 284085
rect 188889 284023 188937 284051
rect 188965 284023 188999 284051
rect 189027 284023 189061 284051
rect 189089 284023 189123 284051
rect 189151 284023 189199 284051
rect 188889 283989 189199 284023
rect 188889 283961 188937 283989
rect 188965 283961 188999 283989
rect 189027 283961 189061 283989
rect 189089 283961 189123 283989
rect 189151 283961 189199 283989
rect 188889 275175 189199 283961
rect 188889 275147 188937 275175
rect 188965 275147 188999 275175
rect 189027 275147 189061 275175
rect 189089 275147 189123 275175
rect 189151 275147 189199 275175
rect 188889 275113 189199 275147
rect 188889 275085 188937 275113
rect 188965 275085 188999 275113
rect 189027 275085 189061 275113
rect 189089 275085 189123 275113
rect 189151 275085 189199 275113
rect 188889 275051 189199 275085
rect 188889 275023 188937 275051
rect 188965 275023 188999 275051
rect 189027 275023 189061 275051
rect 189089 275023 189123 275051
rect 189151 275023 189199 275051
rect 188889 274989 189199 275023
rect 188889 274961 188937 274989
rect 188965 274961 188999 274989
rect 189027 274961 189061 274989
rect 189089 274961 189123 274989
rect 189151 274961 189199 274989
rect 188889 266175 189199 274961
rect 188889 266147 188937 266175
rect 188965 266147 188999 266175
rect 189027 266147 189061 266175
rect 189089 266147 189123 266175
rect 189151 266147 189199 266175
rect 188889 266113 189199 266147
rect 188889 266085 188937 266113
rect 188965 266085 188999 266113
rect 189027 266085 189061 266113
rect 189089 266085 189123 266113
rect 189151 266085 189199 266113
rect 188889 266051 189199 266085
rect 188889 266023 188937 266051
rect 188965 266023 188999 266051
rect 189027 266023 189061 266051
rect 189089 266023 189123 266051
rect 189151 266023 189199 266051
rect 188889 265989 189199 266023
rect 188889 265961 188937 265989
rect 188965 265961 188999 265989
rect 189027 265961 189061 265989
rect 189089 265961 189123 265989
rect 189151 265961 189199 265989
rect 188889 257175 189199 265961
rect 188889 257147 188937 257175
rect 188965 257147 188999 257175
rect 189027 257147 189061 257175
rect 189089 257147 189123 257175
rect 189151 257147 189199 257175
rect 188889 257113 189199 257147
rect 188889 257085 188937 257113
rect 188965 257085 188999 257113
rect 189027 257085 189061 257113
rect 189089 257085 189123 257113
rect 189151 257085 189199 257113
rect 188889 257051 189199 257085
rect 188889 257023 188937 257051
rect 188965 257023 188999 257051
rect 189027 257023 189061 257051
rect 189089 257023 189123 257051
rect 189151 257023 189199 257051
rect 188889 256989 189199 257023
rect 188889 256961 188937 256989
rect 188965 256961 188999 256989
rect 189027 256961 189061 256989
rect 189089 256961 189123 256989
rect 189151 256961 189199 256989
rect 188889 248175 189199 256961
rect 188889 248147 188937 248175
rect 188965 248147 188999 248175
rect 189027 248147 189061 248175
rect 189089 248147 189123 248175
rect 189151 248147 189199 248175
rect 188889 248113 189199 248147
rect 188889 248085 188937 248113
rect 188965 248085 188999 248113
rect 189027 248085 189061 248113
rect 189089 248085 189123 248113
rect 189151 248085 189199 248113
rect 188889 248051 189199 248085
rect 188889 248023 188937 248051
rect 188965 248023 188999 248051
rect 189027 248023 189061 248051
rect 189089 248023 189123 248051
rect 189151 248023 189199 248051
rect 188889 247989 189199 248023
rect 188889 247961 188937 247989
rect 188965 247961 188999 247989
rect 189027 247961 189061 247989
rect 189089 247961 189123 247989
rect 189151 247961 189199 247989
rect 188889 239175 189199 247961
rect 188889 239147 188937 239175
rect 188965 239147 188999 239175
rect 189027 239147 189061 239175
rect 189089 239147 189123 239175
rect 189151 239147 189199 239175
rect 188889 239113 189199 239147
rect 188889 239085 188937 239113
rect 188965 239085 188999 239113
rect 189027 239085 189061 239113
rect 189089 239085 189123 239113
rect 189151 239085 189199 239113
rect 188889 239051 189199 239085
rect 188889 239023 188937 239051
rect 188965 239023 188999 239051
rect 189027 239023 189061 239051
rect 189089 239023 189123 239051
rect 189151 239023 189199 239051
rect 188889 238989 189199 239023
rect 188889 238961 188937 238989
rect 188965 238961 188999 238989
rect 189027 238961 189061 238989
rect 189089 238961 189123 238989
rect 189151 238961 189199 238989
rect 188889 230175 189199 238961
rect 188889 230147 188937 230175
rect 188965 230147 188999 230175
rect 189027 230147 189061 230175
rect 189089 230147 189123 230175
rect 189151 230147 189199 230175
rect 188889 230113 189199 230147
rect 188889 230085 188937 230113
rect 188965 230085 188999 230113
rect 189027 230085 189061 230113
rect 189089 230085 189123 230113
rect 189151 230085 189199 230113
rect 188889 230051 189199 230085
rect 188889 230023 188937 230051
rect 188965 230023 188999 230051
rect 189027 230023 189061 230051
rect 189089 230023 189123 230051
rect 189151 230023 189199 230051
rect 188889 229989 189199 230023
rect 188889 229961 188937 229989
rect 188965 229961 188999 229989
rect 189027 229961 189061 229989
rect 189089 229961 189123 229989
rect 189151 229961 189199 229989
rect 188889 221175 189199 229961
rect 188889 221147 188937 221175
rect 188965 221147 188999 221175
rect 189027 221147 189061 221175
rect 189089 221147 189123 221175
rect 189151 221147 189199 221175
rect 188889 221113 189199 221147
rect 188889 221085 188937 221113
rect 188965 221085 188999 221113
rect 189027 221085 189061 221113
rect 189089 221085 189123 221113
rect 189151 221085 189199 221113
rect 188889 221051 189199 221085
rect 188889 221023 188937 221051
rect 188965 221023 188999 221051
rect 189027 221023 189061 221051
rect 189089 221023 189123 221051
rect 189151 221023 189199 221051
rect 188889 220989 189199 221023
rect 188889 220961 188937 220989
rect 188965 220961 188999 220989
rect 189027 220961 189061 220989
rect 189089 220961 189123 220989
rect 189151 220961 189199 220989
rect 188889 212175 189199 220961
rect 188889 212147 188937 212175
rect 188965 212147 188999 212175
rect 189027 212147 189061 212175
rect 189089 212147 189123 212175
rect 189151 212147 189199 212175
rect 188889 212113 189199 212147
rect 188889 212085 188937 212113
rect 188965 212085 188999 212113
rect 189027 212085 189061 212113
rect 189089 212085 189123 212113
rect 189151 212085 189199 212113
rect 188889 212051 189199 212085
rect 188889 212023 188937 212051
rect 188965 212023 188999 212051
rect 189027 212023 189061 212051
rect 189089 212023 189123 212051
rect 189151 212023 189199 212051
rect 188889 211989 189199 212023
rect 188889 211961 188937 211989
rect 188965 211961 188999 211989
rect 189027 211961 189061 211989
rect 189089 211961 189123 211989
rect 189151 211961 189199 211989
rect 188889 203175 189199 211961
rect 188889 203147 188937 203175
rect 188965 203147 188999 203175
rect 189027 203147 189061 203175
rect 189089 203147 189123 203175
rect 189151 203147 189199 203175
rect 188889 203113 189199 203147
rect 188889 203085 188937 203113
rect 188965 203085 188999 203113
rect 189027 203085 189061 203113
rect 189089 203085 189123 203113
rect 189151 203085 189199 203113
rect 188889 203051 189199 203085
rect 188889 203023 188937 203051
rect 188965 203023 188999 203051
rect 189027 203023 189061 203051
rect 189089 203023 189123 203051
rect 189151 203023 189199 203051
rect 188889 202989 189199 203023
rect 188889 202961 188937 202989
rect 188965 202961 188999 202989
rect 189027 202961 189061 202989
rect 189089 202961 189123 202989
rect 189151 202961 189199 202989
rect 188889 194175 189199 202961
rect 188889 194147 188937 194175
rect 188965 194147 188999 194175
rect 189027 194147 189061 194175
rect 189089 194147 189123 194175
rect 189151 194147 189199 194175
rect 188889 194113 189199 194147
rect 188889 194085 188937 194113
rect 188965 194085 188999 194113
rect 189027 194085 189061 194113
rect 189089 194085 189123 194113
rect 189151 194085 189199 194113
rect 188889 194051 189199 194085
rect 188889 194023 188937 194051
rect 188965 194023 188999 194051
rect 189027 194023 189061 194051
rect 189089 194023 189123 194051
rect 189151 194023 189199 194051
rect 188889 193989 189199 194023
rect 188889 193961 188937 193989
rect 188965 193961 188999 193989
rect 189027 193961 189061 193989
rect 189089 193961 189123 193989
rect 189151 193961 189199 193989
rect 188889 185175 189199 193961
rect 188889 185147 188937 185175
rect 188965 185147 188999 185175
rect 189027 185147 189061 185175
rect 189089 185147 189123 185175
rect 189151 185147 189199 185175
rect 188889 185113 189199 185147
rect 188889 185085 188937 185113
rect 188965 185085 188999 185113
rect 189027 185085 189061 185113
rect 189089 185085 189123 185113
rect 189151 185085 189199 185113
rect 188889 185051 189199 185085
rect 188889 185023 188937 185051
rect 188965 185023 188999 185051
rect 189027 185023 189061 185051
rect 189089 185023 189123 185051
rect 189151 185023 189199 185051
rect 188889 184989 189199 185023
rect 188889 184961 188937 184989
rect 188965 184961 188999 184989
rect 189027 184961 189061 184989
rect 189089 184961 189123 184989
rect 189151 184961 189199 184989
rect 188889 176175 189199 184961
rect 188889 176147 188937 176175
rect 188965 176147 188999 176175
rect 189027 176147 189061 176175
rect 189089 176147 189123 176175
rect 189151 176147 189199 176175
rect 188889 176113 189199 176147
rect 188889 176085 188937 176113
rect 188965 176085 188999 176113
rect 189027 176085 189061 176113
rect 189089 176085 189123 176113
rect 189151 176085 189199 176113
rect 188889 176051 189199 176085
rect 188889 176023 188937 176051
rect 188965 176023 188999 176051
rect 189027 176023 189061 176051
rect 189089 176023 189123 176051
rect 189151 176023 189199 176051
rect 188889 175989 189199 176023
rect 188889 175961 188937 175989
rect 188965 175961 188999 175989
rect 189027 175961 189061 175989
rect 189089 175961 189123 175989
rect 189151 175961 189199 175989
rect 188889 167175 189199 175961
rect 202389 298606 202699 299134
rect 202389 298578 202437 298606
rect 202465 298578 202499 298606
rect 202527 298578 202561 298606
rect 202589 298578 202623 298606
rect 202651 298578 202699 298606
rect 202389 298544 202699 298578
rect 202389 298516 202437 298544
rect 202465 298516 202499 298544
rect 202527 298516 202561 298544
rect 202589 298516 202623 298544
rect 202651 298516 202699 298544
rect 202389 298482 202699 298516
rect 202389 298454 202437 298482
rect 202465 298454 202499 298482
rect 202527 298454 202561 298482
rect 202589 298454 202623 298482
rect 202651 298454 202699 298482
rect 202389 298420 202699 298454
rect 202389 298392 202437 298420
rect 202465 298392 202499 298420
rect 202527 298392 202561 298420
rect 202589 298392 202623 298420
rect 202651 298392 202699 298420
rect 202389 290175 202699 298392
rect 202389 290147 202437 290175
rect 202465 290147 202499 290175
rect 202527 290147 202561 290175
rect 202589 290147 202623 290175
rect 202651 290147 202699 290175
rect 202389 290113 202699 290147
rect 202389 290085 202437 290113
rect 202465 290085 202499 290113
rect 202527 290085 202561 290113
rect 202589 290085 202623 290113
rect 202651 290085 202699 290113
rect 202389 290051 202699 290085
rect 202389 290023 202437 290051
rect 202465 290023 202499 290051
rect 202527 290023 202561 290051
rect 202589 290023 202623 290051
rect 202651 290023 202699 290051
rect 202389 289989 202699 290023
rect 202389 289961 202437 289989
rect 202465 289961 202499 289989
rect 202527 289961 202561 289989
rect 202589 289961 202623 289989
rect 202651 289961 202699 289989
rect 202389 281175 202699 289961
rect 202389 281147 202437 281175
rect 202465 281147 202499 281175
rect 202527 281147 202561 281175
rect 202589 281147 202623 281175
rect 202651 281147 202699 281175
rect 202389 281113 202699 281147
rect 202389 281085 202437 281113
rect 202465 281085 202499 281113
rect 202527 281085 202561 281113
rect 202589 281085 202623 281113
rect 202651 281085 202699 281113
rect 202389 281051 202699 281085
rect 202389 281023 202437 281051
rect 202465 281023 202499 281051
rect 202527 281023 202561 281051
rect 202589 281023 202623 281051
rect 202651 281023 202699 281051
rect 202389 280989 202699 281023
rect 202389 280961 202437 280989
rect 202465 280961 202499 280989
rect 202527 280961 202561 280989
rect 202589 280961 202623 280989
rect 202651 280961 202699 280989
rect 202389 272175 202699 280961
rect 202389 272147 202437 272175
rect 202465 272147 202499 272175
rect 202527 272147 202561 272175
rect 202589 272147 202623 272175
rect 202651 272147 202699 272175
rect 202389 272113 202699 272147
rect 202389 272085 202437 272113
rect 202465 272085 202499 272113
rect 202527 272085 202561 272113
rect 202589 272085 202623 272113
rect 202651 272085 202699 272113
rect 202389 272051 202699 272085
rect 202389 272023 202437 272051
rect 202465 272023 202499 272051
rect 202527 272023 202561 272051
rect 202589 272023 202623 272051
rect 202651 272023 202699 272051
rect 202389 271989 202699 272023
rect 202389 271961 202437 271989
rect 202465 271961 202499 271989
rect 202527 271961 202561 271989
rect 202589 271961 202623 271989
rect 202651 271961 202699 271989
rect 202389 263175 202699 271961
rect 202389 263147 202437 263175
rect 202465 263147 202499 263175
rect 202527 263147 202561 263175
rect 202589 263147 202623 263175
rect 202651 263147 202699 263175
rect 202389 263113 202699 263147
rect 202389 263085 202437 263113
rect 202465 263085 202499 263113
rect 202527 263085 202561 263113
rect 202589 263085 202623 263113
rect 202651 263085 202699 263113
rect 202389 263051 202699 263085
rect 202389 263023 202437 263051
rect 202465 263023 202499 263051
rect 202527 263023 202561 263051
rect 202589 263023 202623 263051
rect 202651 263023 202699 263051
rect 202389 262989 202699 263023
rect 202389 262961 202437 262989
rect 202465 262961 202499 262989
rect 202527 262961 202561 262989
rect 202589 262961 202623 262989
rect 202651 262961 202699 262989
rect 202389 254175 202699 262961
rect 202389 254147 202437 254175
rect 202465 254147 202499 254175
rect 202527 254147 202561 254175
rect 202589 254147 202623 254175
rect 202651 254147 202699 254175
rect 202389 254113 202699 254147
rect 202389 254085 202437 254113
rect 202465 254085 202499 254113
rect 202527 254085 202561 254113
rect 202589 254085 202623 254113
rect 202651 254085 202699 254113
rect 202389 254051 202699 254085
rect 202389 254023 202437 254051
rect 202465 254023 202499 254051
rect 202527 254023 202561 254051
rect 202589 254023 202623 254051
rect 202651 254023 202699 254051
rect 202389 253989 202699 254023
rect 202389 253961 202437 253989
rect 202465 253961 202499 253989
rect 202527 253961 202561 253989
rect 202589 253961 202623 253989
rect 202651 253961 202699 253989
rect 202389 245175 202699 253961
rect 202389 245147 202437 245175
rect 202465 245147 202499 245175
rect 202527 245147 202561 245175
rect 202589 245147 202623 245175
rect 202651 245147 202699 245175
rect 202389 245113 202699 245147
rect 202389 245085 202437 245113
rect 202465 245085 202499 245113
rect 202527 245085 202561 245113
rect 202589 245085 202623 245113
rect 202651 245085 202699 245113
rect 202389 245051 202699 245085
rect 202389 245023 202437 245051
rect 202465 245023 202499 245051
rect 202527 245023 202561 245051
rect 202589 245023 202623 245051
rect 202651 245023 202699 245051
rect 202389 244989 202699 245023
rect 202389 244961 202437 244989
rect 202465 244961 202499 244989
rect 202527 244961 202561 244989
rect 202589 244961 202623 244989
rect 202651 244961 202699 244989
rect 202389 236175 202699 244961
rect 202389 236147 202437 236175
rect 202465 236147 202499 236175
rect 202527 236147 202561 236175
rect 202589 236147 202623 236175
rect 202651 236147 202699 236175
rect 202389 236113 202699 236147
rect 202389 236085 202437 236113
rect 202465 236085 202499 236113
rect 202527 236085 202561 236113
rect 202589 236085 202623 236113
rect 202651 236085 202699 236113
rect 202389 236051 202699 236085
rect 202389 236023 202437 236051
rect 202465 236023 202499 236051
rect 202527 236023 202561 236051
rect 202589 236023 202623 236051
rect 202651 236023 202699 236051
rect 202389 235989 202699 236023
rect 202389 235961 202437 235989
rect 202465 235961 202499 235989
rect 202527 235961 202561 235989
rect 202589 235961 202623 235989
rect 202651 235961 202699 235989
rect 202389 227175 202699 235961
rect 202389 227147 202437 227175
rect 202465 227147 202499 227175
rect 202527 227147 202561 227175
rect 202589 227147 202623 227175
rect 202651 227147 202699 227175
rect 202389 227113 202699 227147
rect 202389 227085 202437 227113
rect 202465 227085 202499 227113
rect 202527 227085 202561 227113
rect 202589 227085 202623 227113
rect 202651 227085 202699 227113
rect 202389 227051 202699 227085
rect 202389 227023 202437 227051
rect 202465 227023 202499 227051
rect 202527 227023 202561 227051
rect 202589 227023 202623 227051
rect 202651 227023 202699 227051
rect 202389 226989 202699 227023
rect 202389 226961 202437 226989
rect 202465 226961 202499 226989
rect 202527 226961 202561 226989
rect 202589 226961 202623 226989
rect 202651 226961 202699 226989
rect 202389 218175 202699 226961
rect 202389 218147 202437 218175
rect 202465 218147 202499 218175
rect 202527 218147 202561 218175
rect 202589 218147 202623 218175
rect 202651 218147 202699 218175
rect 202389 218113 202699 218147
rect 202389 218085 202437 218113
rect 202465 218085 202499 218113
rect 202527 218085 202561 218113
rect 202589 218085 202623 218113
rect 202651 218085 202699 218113
rect 202389 218051 202699 218085
rect 202389 218023 202437 218051
rect 202465 218023 202499 218051
rect 202527 218023 202561 218051
rect 202589 218023 202623 218051
rect 202651 218023 202699 218051
rect 202389 217989 202699 218023
rect 202389 217961 202437 217989
rect 202465 217961 202499 217989
rect 202527 217961 202561 217989
rect 202589 217961 202623 217989
rect 202651 217961 202699 217989
rect 202389 209175 202699 217961
rect 202389 209147 202437 209175
rect 202465 209147 202499 209175
rect 202527 209147 202561 209175
rect 202589 209147 202623 209175
rect 202651 209147 202699 209175
rect 202389 209113 202699 209147
rect 202389 209085 202437 209113
rect 202465 209085 202499 209113
rect 202527 209085 202561 209113
rect 202589 209085 202623 209113
rect 202651 209085 202699 209113
rect 202389 209051 202699 209085
rect 202389 209023 202437 209051
rect 202465 209023 202499 209051
rect 202527 209023 202561 209051
rect 202589 209023 202623 209051
rect 202651 209023 202699 209051
rect 202389 208989 202699 209023
rect 202389 208961 202437 208989
rect 202465 208961 202499 208989
rect 202527 208961 202561 208989
rect 202589 208961 202623 208989
rect 202651 208961 202699 208989
rect 202389 200175 202699 208961
rect 202389 200147 202437 200175
rect 202465 200147 202499 200175
rect 202527 200147 202561 200175
rect 202589 200147 202623 200175
rect 202651 200147 202699 200175
rect 202389 200113 202699 200147
rect 202389 200085 202437 200113
rect 202465 200085 202499 200113
rect 202527 200085 202561 200113
rect 202589 200085 202623 200113
rect 202651 200085 202699 200113
rect 202389 200051 202699 200085
rect 202389 200023 202437 200051
rect 202465 200023 202499 200051
rect 202527 200023 202561 200051
rect 202589 200023 202623 200051
rect 202651 200023 202699 200051
rect 202389 199989 202699 200023
rect 202389 199961 202437 199989
rect 202465 199961 202499 199989
rect 202527 199961 202561 199989
rect 202589 199961 202623 199989
rect 202651 199961 202699 199989
rect 202389 191175 202699 199961
rect 202389 191147 202437 191175
rect 202465 191147 202499 191175
rect 202527 191147 202561 191175
rect 202589 191147 202623 191175
rect 202651 191147 202699 191175
rect 202389 191113 202699 191147
rect 202389 191085 202437 191113
rect 202465 191085 202499 191113
rect 202527 191085 202561 191113
rect 202589 191085 202623 191113
rect 202651 191085 202699 191113
rect 202389 191051 202699 191085
rect 202389 191023 202437 191051
rect 202465 191023 202499 191051
rect 202527 191023 202561 191051
rect 202589 191023 202623 191051
rect 202651 191023 202699 191051
rect 202389 190989 202699 191023
rect 202389 190961 202437 190989
rect 202465 190961 202499 190989
rect 202527 190961 202561 190989
rect 202589 190961 202623 190989
rect 202651 190961 202699 190989
rect 202389 182175 202699 190961
rect 202389 182147 202437 182175
rect 202465 182147 202499 182175
rect 202527 182147 202561 182175
rect 202589 182147 202623 182175
rect 202651 182147 202699 182175
rect 202389 182113 202699 182147
rect 202389 182085 202437 182113
rect 202465 182085 202499 182113
rect 202527 182085 202561 182113
rect 202589 182085 202623 182113
rect 202651 182085 202699 182113
rect 202389 182051 202699 182085
rect 202389 182023 202437 182051
rect 202465 182023 202499 182051
rect 202527 182023 202561 182051
rect 202589 182023 202623 182051
rect 202651 182023 202699 182051
rect 202389 181989 202699 182023
rect 202389 181961 202437 181989
rect 202465 181961 202499 181989
rect 202527 181961 202561 181989
rect 202589 181961 202623 181989
rect 202651 181961 202699 181989
rect 192544 173175 192704 173192
rect 192544 173147 192579 173175
rect 192607 173147 192641 173175
rect 192669 173147 192704 173175
rect 192544 173113 192704 173147
rect 192544 173085 192579 173113
rect 192607 173085 192641 173113
rect 192669 173085 192704 173113
rect 192544 173051 192704 173085
rect 192544 173023 192579 173051
rect 192607 173023 192641 173051
rect 192669 173023 192704 173051
rect 192544 172989 192704 173023
rect 192544 172961 192579 172989
rect 192607 172961 192641 172989
rect 192669 172961 192704 172989
rect 192544 172944 192704 172961
rect 202389 173175 202699 181961
rect 202389 173147 202437 173175
rect 202465 173147 202499 173175
rect 202527 173147 202561 173175
rect 202589 173147 202623 173175
rect 202651 173147 202699 173175
rect 202389 173113 202699 173147
rect 202389 173085 202437 173113
rect 202465 173085 202499 173113
rect 202527 173085 202561 173113
rect 202589 173085 202623 173113
rect 202651 173085 202699 173113
rect 202389 173051 202699 173085
rect 202389 173023 202437 173051
rect 202465 173023 202499 173051
rect 202527 173023 202561 173051
rect 202589 173023 202623 173051
rect 202651 173023 202699 173051
rect 202389 172989 202699 173023
rect 202389 172961 202437 172989
rect 202465 172961 202499 172989
rect 202527 172961 202561 172989
rect 202589 172961 202623 172989
rect 202651 172961 202699 172989
rect 188889 167147 188937 167175
rect 188965 167147 188999 167175
rect 189027 167147 189061 167175
rect 189089 167147 189123 167175
rect 189151 167147 189199 167175
rect 188889 167113 189199 167147
rect 188889 167085 188937 167113
rect 188965 167085 188999 167113
rect 189027 167085 189061 167113
rect 189089 167085 189123 167113
rect 189151 167085 189199 167113
rect 188889 167051 189199 167085
rect 188889 167023 188937 167051
rect 188965 167023 188999 167051
rect 189027 167023 189061 167051
rect 189089 167023 189123 167051
rect 189151 167023 189199 167051
rect 188889 166989 189199 167023
rect 188889 166961 188937 166989
rect 188965 166961 188999 166989
rect 189027 166961 189061 166989
rect 189089 166961 189123 166989
rect 189151 166961 189199 166989
rect 188889 158175 189199 166961
rect 200224 167175 200384 167192
rect 200224 167147 200259 167175
rect 200287 167147 200321 167175
rect 200349 167147 200384 167175
rect 200224 167113 200384 167147
rect 200224 167085 200259 167113
rect 200287 167085 200321 167113
rect 200349 167085 200384 167113
rect 200224 167051 200384 167085
rect 200224 167023 200259 167051
rect 200287 167023 200321 167051
rect 200349 167023 200384 167051
rect 200224 166989 200384 167023
rect 200224 166961 200259 166989
rect 200287 166961 200321 166989
rect 200349 166961 200384 166989
rect 200224 166944 200384 166961
rect 192544 164175 192704 164192
rect 192544 164147 192579 164175
rect 192607 164147 192641 164175
rect 192669 164147 192704 164175
rect 192544 164113 192704 164147
rect 192544 164085 192579 164113
rect 192607 164085 192641 164113
rect 192669 164085 192704 164113
rect 192544 164051 192704 164085
rect 192544 164023 192579 164051
rect 192607 164023 192641 164051
rect 192669 164023 192704 164051
rect 192544 163989 192704 164023
rect 192544 163961 192579 163989
rect 192607 163961 192641 163989
rect 192669 163961 192704 163989
rect 192544 163944 192704 163961
rect 202389 164175 202699 172961
rect 202389 164147 202437 164175
rect 202465 164147 202499 164175
rect 202527 164147 202561 164175
rect 202589 164147 202623 164175
rect 202651 164147 202699 164175
rect 202389 164113 202699 164147
rect 202389 164085 202437 164113
rect 202465 164085 202499 164113
rect 202527 164085 202561 164113
rect 202589 164085 202623 164113
rect 202651 164085 202699 164113
rect 202389 164051 202699 164085
rect 202389 164023 202437 164051
rect 202465 164023 202499 164051
rect 202527 164023 202561 164051
rect 202589 164023 202623 164051
rect 202651 164023 202699 164051
rect 202389 163989 202699 164023
rect 202389 163961 202437 163989
rect 202465 163961 202499 163989
rect 202527 163961 202561 163989
rect 202589 163961 202623 163989
rect 202651 163961 202699 163989
rect 188889 158147 188937 158175
rect 188965 158147 188999 158175
rect 189027 158147 189061 158175
rect 189089 158147 189123 158175
rect 189151 158147 189199 158175
rect 188889 158113 189199 158147
rect 188889 158085 188937 158113
rect 188965 158085 188999 158113
rect 189027 158085 189061 158113
rect 189089 158085 189123 158113
rect 189151 158085 189199 158113
rect 188889 158051 189199 158085
rect 188889 158023 188937 158051
rect 188965 158023 188999 158051
rect 189027 158023 189061 158051
rect 189089 158023 189123 158051
rect 189151 158023 189199 158051
rect 188889 157989 189199 158023
rect 188889 157961 188937 157989
rect 188965 157961 188999 157989
rect 189027 157961 189061 157989
rect 189089 157961 189123 157989
rect 189151 157961 189199 157989
rect 188889 149175 189199 157961
rect 200224 158175 200384 158192
rect 200224 158147 200259 158175
rect 200287 158147 200321 158175
rect 200349 158147 200384 158175
rect 200224 158113 200384 158147
rect 200224 158085 200259 158113
rect 200287 158085 200321 158113
rect 200349 158085 200384 158113
rect 200224 158051 200384 158085
rect 200224 158023 200259 158051
rect 200287 158023 200321 158051
rect 200349 158023 200384 158051
rect 200224 157989 200384 158023
rect 200224 157961 200259 157989
rect 200287 157961 200321 157989
rect 200349 157961 200384 157989
rect 200224 157944 200384 157961
rect 192544 155175 192704 155192
rect 192544 155147 192579 155175
rect 192607 155147 192641 155175
rect 192669 155147 192704 155175
rect 192544 155113 192704 155147
rect 192544 155085 192579 155113
rect 192607 155085 192641 155113
rect 192669 155085 192704 155113
rect 192544 155051 192704 155085
rect 192544 155023 192579 155051
rect 192607 155023 192641 155051
rect 192669 155023 192704 155051
rect 192544 154989 192704 155023
rect 192544 154961 192579 154989
rect 192607 154961 192641 154989
rect 192669 154961 192704 154989
rect 192544 154944 192704 154961
rect 202389 155175 202699 163961
rect 202389 155147 202437 155175
rect 202465 155147 202499 155175
rect 202527 155147 202561 155175
rect 202589 155147 202623 155175
rect 202651 155147 202699 155175
rect 202389 155113 202699 155147
rect 202389 155085 202437 155113
rect 202465 155085 202499 155113
rect 202527 155085 202561 155113
rect 202589 155085 202623 155113
rect 202651 155085 202699 155113
rect 202389 155051 202699 155085
rect 202389 155023 202437 155051
rect 202465 155023 202499 155051
rect 202527 155023 202561 155051
rect 202589 155023 202623 155051
rect 202651 155023 202699 155051
rect 202389 154989 202699 155023
rect 202389 154961 202437 154989
rect 202465 154961 202499 154989
rect 202527 154961 202561 154989
rect 202589 154961 202623 154989
rect 202651 154961 202699 154989
rect 188889 149147 188937 149175
rect 188965 149147 188999 149175
rect 189027 149147 189061 149175
rect 189089 149147 189123 149175
rect 189151 149147 189199 149175
rect 188889 149113 189199 149147
rect 188889 149085 188937 149113
rect 188965 149085 188999 149113
rect 189027 149085 189061 149113
rect 189089 149085 189123 149113
rect 189151 149085 189199 149113
rect 188889 149051 189199 149085
rect 188889 149023 188937 149051
rect 188965 149023 188999 149051
rect 189027 149023 189061 149051
rect 189089 149023 189123 149051
rect 189151 149023 189199 149051
rect 188889 148989 189199 149023
rect 188889 148961 188937 148989
rect 188965 148961 188999 148989
rect 189027 148961 189061 148989
rect 189089 148961 189123 148989
rect 189151 148961 189199 148989
rect 188889 140175 189199 148961
rect 200224 149175 200384 149192
rect 200224 149147 200259 149175
rect 200287 149147 200321 149175
rect 200349 149147 200384 149175
rect 200224 149113 200384 149147
rect 200224 149085 200259 149113
rect 200287 149085 200321 149113
rect 200349 149085 200384 149113
rect 200224 149051 200384 149085
rect 200224 149023 200259 149051
rect 200287 149023 200321 149051
rect 200349 149023 200384 149051
rect 200224 148989 200384 149023
rect 200224 148961 200259 148989
rect 200287 148961 200321 148989
rect 200349 148961 200384 148989
rect 200224 148944 200384 148961
rect 192544 146175 192704 146192
rect 192544 146147 192579 146175
rect 192607 146147 192641 146175
rect 192669 146147 192704 146175
rect 192544 146113 192704 146147
rect 192544 146085 192579 146113
rect 192607 146085 192641 146113
rect 192669 146085 192704 146113
rect 192544 146051 192704 146085
rect 192544 146023 192579 146051
rect 192607 146023 192641 146051
rect 192669 146023 192704 146051
rect 192544 145989 192704 146023
rect 192544 145961 192579 145989
rect 192607 145961 192641 145989
rect 192669 145961 192704 145989
rect 192544 145944 192704 145961
rect 202389 146175 202699 154961
rect 202389 146147 202437 146175
rect 202465 146147 202499 146175
rect 202527 146147 202561 146175
rect 202589 146147 202623 146175
rect 202651 146147 202699 146175
rect 202389 146113 202699 146147
rect 202389 146085 202437 146113
rect 202465 146085 202499 146113
rect 202527 146085 202561 146113
rect 202589 146085 202623 146113
rect 202651 146085 202699 146113
rect 202389 146051 202699 146085
rect 202389 146023 202437 146051
rect 202465 146023 202499 146051
rect 202527 146023 202561 146051
rect 202589 146023 202623 146051
rect 202651 146023 202699 146051
rect 202389 145989 202699 146023
rect 202389 145961 202437 145989
rect 202465 145961 202499 145989
rect 202527 145961 202561 145989
rect 202589 145961 202623 145989
rect 202651 145961 202699 145989
rect 188889 140147 188937 140175
rect 188965 140147 188999 140175
rect 189027 140147 189061 140175
rect 189089 140147 189123 140175
rect 189151 140147 189199 140175
rect 188889 140113 189199 140147
rect 188889 140085 188937 140113
rect 188965 140085 188999 140113
rect 189027 140085 189061 140113
rect 189089 140085 189123 140113
rect 189151 140085 189199 140113
rect 188889 140051 189199 140085
rect 188889 140023 188937 140051
rect 188965 140023 188999 140051
rect 189027 140023 189061 140051
rect 189089 140023 189123 140051
rect 189151 140023 189199 140051
rect 188889 139989 189199 140023
rect 188889 139961 188937 139989
rect 188965 139961 188999 139989
rect 189027 139961 189061 139989
rect 189089 139961 189123 139989
rect 189151 139961 189199 139989
rect 188889 131175 189199 139961
rect 200224 140175 200384 140192
rect 200224 140147 200259 140175
rect 200287 140147 200321 140175
rect 200349 140147 200384 140175
rect 200224 140113 200384 140147
rect 200224 140085 200259 140113
rect 200287 140085 200321 140113
rect 200349 140085 200384 140113
rect 200224 140051 200384 140085
rect 200224 140023 200259 140051
rect 200287 140023 200321 140051
rect 200349 140023 200384 140051
rect 200224 139989 200384 140023
rect 200224 139961 200259 139989
rect 200287 139961 200321 139989
rect 200349 139961 200384 139989
rect 200224 139944 200384 139961
rect 192544 137175 192704 137192
rect 192544 137147 192579 137175
rect 192607 137147 192641 137175
rect 192669 137147 192704 137175
rect 192544 137113 192704 137147
rect 192544 137085 192579 137113
rect 192607 137085 192641 137113
rect 192669 137085 192704 137113
rect 192544 137051 192704 137085
rect 192544 137023 192579 137051
rect 192607 137023 192641 137051
rect 192669 137023 192704 137051
rect 192544 136989 192704 137023
rect 192544 136961 192579 136989
rect 192607 136961 192641 136989
rect 192669 136961 192704 136989
rect 192544 136944 192704 136961
rect 202389 137175 202699 145961
rect 202389 137147 202437 137175
rect 202465 137147 202499 137175
rect 202527 137147 202561 137175
rect 202589 137147 202623 137175
rect 202651 137147 202699 137175
rect 202389 137113 202699 137147
rect 202389 137085 202437 137113
rect 202465 137085 202499 137113
rect 202527 137085 202561 137113
rect 202589 137085 202623 137113
rect 202651 137085 202699 137113
rect 202389 137051 202699 137085
rect 202389 137023 202437 137051
rect 202465 137023 202499 137051
rect 202527 137023 202561 137051
rect 202589 137023 202623 137051
rect 202651 137023 202699 137051
rect 202389 136989 202699 137023
rect 202389 136961 202437 136989
rect 202465 136961 202499 136989
rect 202527 136961 202561 136989
rect 202589 136961 202623 136989
rect 202651 136961 202699 136989
rect 188889 131147 188937 131175
rect 188965 131147 188999 131175
rect 189027 131147 189061 131175
rect 189089 131147 189123 131175
rect 189151 131147 189199 131175
rect 188889 131113 189199 131147
rect 188889 131085 188937 131113
rect 188965 131085 188999 131113
rect 189027 131085 189061 131113
rect 189089 131085 189123 131113
rect 189151 131085 189199 131113
rect 188889 131051 189199 131085
rect 188889 131023 188937 131051
rect 188965 131023 188999 131051
rect 189027 131023 189061 131051
rect 189089 131023 189123 131051
rect 189151 131023 189199 131051
rect 188889 130989 189199 131023
rect 188889 130961 188937 130989
rect 188965 130961 188999 130989
rect 189027 130961 189061 130989
rect 189089 130961 189123 130989
rect 189151 130961 189199 130989
rect 188889 122175 189199 130961
rect 200224 131175 200384 131192
rect 200224 131147 200259 131175
rect 200287 131147 200321 131175
rect 200349 131147 200384 131175
rect 200224 131113 200384 131147
rect 200224 131085 200259 131113
rect 200287 131085 200321 131113
rect 200349 131085 200384 131113
rect 200224 131051 200384 131085
rect 200224 131023 200259 131051
rect 200287 131023 200321 131051
rect 200349 131023 200384 131051
rect 200224 130989 200384 131023
rect 200224 130961 200259 130989
rect 200287 130961 200321 130989
rect 200349 130961 200384 130989
rect 200224 130944 200384 130961
rect 192544 128175 192704 128192
rect 192544 128147 192579 128175
rect 192607 128147 192641 128175
rect 192669 128147 192704 128175
rect 192544 128113 192704 128147
rect 192544 128085 192579 128113
rect 192607 128085 192641 128113
rect 192669 128085 192704 128113
rect 192544 128051 192704 128085
rect 192544 128023 192579 128051
rect 192607 128023 192641 128051
rect 192669 128023 192704 128051
rect 192544 127989 192704 128023
rect 192544 127961 192579 127989
rect 192607 127961 192641 127989
rect 192669 127961 192704 127989
rect 192544 127944 192704 127961
rect 202389 128175 202699 136961
rect 202389 128147 202437 128175
rect 202465 128147 202499 128175
rect 202527 128147 202561 128175
rect 202589 128147 202623 128175
rect 202651 128147 202699 128175
rect 202389 128113 202699 128147
rect 202389 128085 202437 128113
rect 202465 128085 202499 128113
rect 202527 128085 202561 128113
rect 202589 128085 202623 128113
rect 202651 128085 202699 128113
rect 202389 128051 202699 128085
rect 202389 128023 202437 128051
rect 202465 128023 202499 128051
rect 202527 128023 202561 128051
rect 202589 128023 202623 128051
rect 202651 128023 202699 128051
rect 202389 127989 202699 128023
rect 202389 127961 202437 127989
rect 202465 127961 202499 127989
rect 202527 127961 202561 127989
rect 202589 127961 202623 127989
rect 202651 127961 202699 127989
rect 188889 122147 188937 122175
rect 188965 122147 188999 122175
rect 189027 122147 189061 122175
rect 189089 122147 189123 122175
rect 189151 122147 189199 122175
rect 188889 122113 189199 122147
rect 188889 122085 188937 122113
rect 188965 122085 188999 122113
rect 189027 122085 189061 122113
rect 189089 122085 189123 122113
rect 189151 122085 189199 122113
rect 188889 122051 189199 122085
rect 188889 122023 188937 122051
rect 188965 122023 188999 122051
rect 189027 122023 189061 122051
rect 189089 122023 189123 122051
rect 189151 122023 189199 122051
rect 188889 121989 189199 122023
rect 188889 121961 188937 121989
rect 188965 121961 188999 121989
rect 189027 121961 189061 121989
rect 189089 121961 189123 121989
rect 189151 121961 189199 121989
rect 188889 113175 189199 121961
rect 200224 122175 200384 122192
rect 200224 122147 200259 122175
rect 200287 122147 200321 122175
rect 200349 122147 200384 122175
rect 200224 122113 200384 122147
rect 200224 122085 200259 122113
rect 200287 122085 200321 122113
rect 200349 122085 200384 122113
rect 200224 122051 200384 122085
rect 200224 122023 200259 122051
rect 200287 122023 200321 122051
rect 200349 122023 200384 122051
rect 200224 121989 200384 122023
rect 200224 121961 200259 121989
rect 200287 121961 200321 121989
rect 200349 121961 200384 121989
rect 200224 121944 200384 121961
rect 192544 119175 192704 119192
rect 192544 119147 192579 119175
rect 192607 119147 192641 119175
rect 192669 119147 192704 119175
rect 192544 119113 192704 119147
rect 192544 119085 192579 119113
rect 192607 119085 192641 119113
rect 192669 119085 192704 119113
rect 192544 119051 192704 119085
rect 192544 119023 192579 119051
rect 192607 119023 192641 119051
rect 192669 119023 192704 119051
rect 192544 118989 192704 119023
rect 192544 118961 192579 118989
rect 192607 118961 192641 118989
rect 192669 118961 192704 118989
rect 192544 118944 192704 118961
rect 202389 119175 202699 127961
rect 202389 119147 202437 119175
rect 202465 119147 202499 119175
rect 202527 119147 202561 119175
rect 202589 119147 202623 119175
rect 202651 119147 202699 119175
rect 202389 119113 202699 119147
rect 202389 119085 202437 119113
rect 202465 119085 202499 119113
rect 202527 119085 202561 119113
rect 202589 119085 202623 119113
rect 202651 119085 202699 119113
rect 202389 119051 202699 119085
rect 202389 119023 202437 119051
rect 202465 119023 202499 119051
rect 202527 119023 202561 119051
rect 202589 119023 202623 119051
rect 202651 119023 202699 119051
rect 202389 118989 202699 119023
rect 202389 118961 202437 118989
rect 202465 118961 202499 118989
rect 202527 118961 202561 118989
rect 202589 118961 202623 118989
rect 202651 118961 202699 118989
rect 188889 113147 188937 113175
rect 188965 113147 188999 113175
rect 189027 113147 189061 113175
rect 189089 113147 189123 113175
rect 189151 113147 189199 113175
rect 188889 113113 189199 113147
rect 188889 113085 188937 113113
rect 188965 113085 188999 113113
rect 189027 113085 189061 113113
rect 189089 113085 189123 113113
rect 189151 113085 189199 113113
rect 188889 113051 189199 113085
rect 188889 113023 188937 113051
rect 188965 113023 188999 113051
rect 189027 113023 189061 113051
rect 189089 113023 189123 113051
rect 189151 113023 189199 113051
rect 188889 112989 189199 113023
rect 188889 112961 188937 112989
rect 188965 112961 188999 112989
rect 189027 112961 189061 112989
rect 189089 112961 189123 112989
rect 189151 112961 189199 112989
rect 188889 104175 189199 112961
rect 200224 113175 200384 113192
rect 200224 113147 200259 113175
rect 200287 113147 200321 113175
rect 200349 113147 200384 113175
rect 200224 113113 200384 113147
rect 200224 113085 200259 113113
rect 200287 113085 200321 113113
rect 200349 113085 200384 113113
rect 200224 113051 200384 113085
rect 200224 113023 200259 113051
rect 200287 113023 200321 113051
rect 200349 113023 200384 113051
rect 200224 112989 200384 113023
rect 200224 112961 200259 112989
rect 200287 112961 200321 112989
rect 200349 112961 200384 112989
rect 200224 112944 200384 112961
rect 192544 110175 192704 110192
rect 192544 110147 192579 110175
rect 192607 110147 192641 110175
rect 192669 110147 192704 110175
rect 192544 110113 192704 110147
rect 192544 110085 192579 110113
rect 192607 110085 192641 110113
rect 192669 110085 192704 110113
rect 192544 110051 192704 110085
rect 192544 110023 192579 110051
rect 192607 110023 192641 110051
rect 192669 110023 192704 110051
rect 192544 109989 192704 110023
rect 192544 109961 192579 109989
rect 192607 109961 192641 109989
rect 192669 109961 192704 109989
rect 192544 109944 192704 109961
rect 202389 110175 202699 118961
rect 202389 110147 202437 110175
rect 202465 110147 202499 110175
rect 202527 110147 202561 110175
rect 202589 110147 202623 110175
rect 202651 110147 202699 110175
rect 202389 110113 202699 110147
rect 202389 110085 202437 110113
rect 202465 110085 202499 110113
rect 202527 110085 202561 110113
rect 202589 110085 202623 110113
rect 202651 110085 202699 110113
rect 202389 110051 202699 110085
rect 202389 110023 202437 110051
rect 202465 110023 202499 110051
rect 202527 110023 202561 110051
rect 202589 110023 202623 110051
rect 202651 110023 202699 110051
rect 202389 109989 202699 110023
rect 202389 109961 202437 109989
rect 202465 109961 202499 109989
rect 202527 109961 202561 109989
rect 202589 109961 202623 109989
rect 202651 109961 202699 109989
rect 188889 104147 188937 104175
rect 188965 104147 188999 104175
rect 189027 104147 189061 104175
rect 189089 104147 189123 104175
rect 189151 104147 189199 104175
rect 188889 104113 189199 104147
rect 188889 104085 188937 104113
rect 188965 104085 188999 104113
rect 189027 104085 189061 104113
rect 189089 104085 189123 104113
rect 189151 104085 189199 104113
rect 188889 104051 189199 104085
rect 188889 104023 188937 104051
rect 188965 104023 188999 104051
rect 189027 104023 189061 104051
rect 189089 104023 189123 104051
rect 189151 104023 189199 104051
rect 188889 103989 189199 104023
rect 188889 103961 188937 103989
rect 188965 103961 188999 103989
rect 189027 103961 189061 103989
rect 189089 103961 189123 103989
rect 189151 103961 189199 103989
rect 188889 95175 189199 103961
rect 200224 104175 200384 104192
rect 200224 104147 200259 104175
rect 200287 104147 200321 104175
rect 200349 104147 200384 104175
rect 200224 104113 200384 104147
rect 200224 104085 200259 104113
rect 200287 104085 200321 104113
rect 200349 104085 200384 104113
rect 200224 104051 200384 104085
rect 200224 104023 200259 104051
rect 200287 104023 200321 104051
rect 200349 104023 200384 104051
rect 200224 103989 200384 104023
rect 200224 103961 200259 103989
rect 200287 103961 200321 103989
rect 200349 103961 200384 103989
rect 200224 103944 200384 103961
rect 192544 101175 192704 101192
rect 192544 101147 192579 101175
rect 192607 101147 192641 101175
rect 192669 101147 192704 101175
rect 192544 101113 192704 101147
rect 192544 101085 192579 101113
rect 192607 101085 192641 101113
rect 192669 101085 192704 101113
rect 192544 101051 192704 101085
rect 192544 101023 192579 101051
rect 192607 101023 192641 101051
rect 192669 101023 192704 101051
rect 192544 100989 192704 101023
rect 192544 100961 192579 100989
rect 192607 100961 192641 100989
rect 192669 100961 192704 100989
rect 192544 100944 192704 100961
rect 202389 101175 202699 109961
rect 202389 101147 202437 101175
rect 202465 101147 202499 101175
rect 202527 101147 202561 101175
rect 202589 101147 202623 101175
rect 202651 101147 202699 101175
rect 202389 101113 202699 101147
rect 202389 101085 202437 101113
rect 202465 101085 202499 101113
rect 202527 101085 202561 101113
rect 202589 101085 202623 101113
rect 202651 101085 202699 101113
rect 202389 101051 202699 101085
rect 202389 101023 202437 101051
rect 202465 101023 202499 101051
rect 202527 101023 202561 101051
rect 202589 101023 202623 101051
rect 202651 101023 202699 101051
rect 202389 100989 202699 101023
rect 202389 100961 202437 100989
rect 202465 100961 202499 100989
rect 202527 100961 202561 100989
rect 202589 100961 202623 100989
rect 202651 100961 202699 100989
rect 188889 95147 188937 95175
rect 188965 95147 188999 95175
rect 189027 95147 189061 95175
rect 189089 95147 189123 95175
rect 189151 95147 189199 95175
rect 188889 95113 189199 95147
rect 188889 95085 188937 95113
rect 188965 95085 188999 95113
rect 189027 95085 189061 95113
rect 189089 95085 189123 95113
rect 189151 95085 189199 95113
rect 188889 95051 189199 95085
rect 188889 95023 188937 95051
rect 188965 95023 188999 95051
rect 189027 95023 189061 95051
rect 189089 95023 189123 95051
rect 189151 95023 189199 95051
rect 188889 94989 189199 95023
rect 188889 94961 188937 94989
rect 188965 94961 188999 94989
rect 189027 94961 189061 94989
rect 189089 94961 189123 94989
rect 189151 94961 189199 94989
rect 188889 86175 189199 94961
rect 200224 95175 200384 95192
rect 200224 95147 200259 95175
rect 200287 95147 200321 95175
rect 200349 95147 200384 95175
rect 200224 95113 200384 95147
rect 200224 95085 200259 95113
rect 200287 95085 200321 95113
rect 200349 95085 200384 95113
rect 200224 95051 200384 95085
rect 200224 95023 200259 95051
rect 200287 95023 200321 95051
rect 200349 95023 200384 95051
rect 200224 94989 200384 95023
rect 200224 94961 200259 94989
rect 200287 94961 200321 94989
rect 200349 94961 200384 94989
rect 200224 94944 200384 94961
rect 192544 92175 192704 92192
rect 192544 92147 192579 92175
rect 192607 92147 192641 92175
rect 192669 92147 192704 92175
rect 192544 92113 192704 92147
rect 192544 92085 192579 92113
rect 192607 92085 192641 92113
rect 192669 92085 192704 92113
rect 192544 92051 192704 92085
rect 192544 92023 192579 92051
rect 192607 92023 192641 92051
rect 192669 92023 192704 92051
rect 192544 91989 192704 92023
rect 192544 91961 192579 91989
rect 192607 91961 192641 91989
rect 192669 91961 192704 91989
rect 192544 91944 192704 91961
rect 202389 92175 202699 100961
rect 202389 92147 202437 92175
rect 202465 92147 202499 92175
rect 202527 92147 202561 92175
rect 202589 92147 202623 92175
rect 202651 92147 202699 92175
rect 202389 92113 202699 92147
rect 202389 92085 202437 92113
rect 202465 92085 202499 92113
rect 202527 92085 202561 92113
rect 202589 92085 202623 92113
rect 202651 92085 202699 92113
rect 202389 92051 202699 92085
rect 202389 92023 202437 92051
rect 202465 92023 202499 92051
rect 202527 92023 202561 92051
rect 202589 92023 202623 92051
rect 202651 92023 202699 92051
rect 202389 91989 202699 92023
rect 202389 91961 202437 91989
rect 202465 91961 202499 91989
rect 202527 91961 202561 91989
rect 202589 91961 202623 91989
rect 202651 91961 202699 91989
rect 188889 86147 188937 86175
rect 188965 86147 188999 86175
rect 189027 86147 189061 86175
rect 189089 86147 189123 86175
rect 189151 86147 189199 86175
rect 188889 86113 189199 86147
rect 188889 86085 188937 86113
rect 188965 86085 188999 86113
rect 189027 86085 189061 86113
rect 189089 86085 189123 86113
rect 189151 86085 189199 86113
rect 188889 86051 189199 86085
rect 188889 86023 188937 86051
rect 188965 86023 188999 86051
rect 189027 86023 189061 86051
rect 189089 86023 189123 86051
rect 189151 86023 189199 86051
rect 188889 85989 189199 86023
rect 188889 85961 188937 85989
rect 188965 85961 188999 85989
rect 189027 85961 189061 85989
rect 189089 85961 189123 85989
rect 189151 85961 189199 85989
rect 188889 77175 189199 85961
rect 200224 86175 200384 86192
rect 200224 86147 200259 86175
rect 200287 86147 200321 86175
rect 200349 86147 200384 86175
rect 200224 86113 200384 86147
rect 200224 86085 200259 86113
rect 200287 86085 200321 86113
rect 200349 86085 200384 86113
rect 200224 86051 200384 86085
rect 200224 86023 200259 86051
rect 200287 86023 200321 86051
rect 200349 86023 200384 86051
rect 200224 85989 200384 86023
rect 200224 85961 200259 85989
rect 200287 85961 200321 85989
rect 200349 85961 200384 85989
rect 200224 85944 200384 85961
rect 192544 83175 192704 83192
rect 192544 83147 192579 83175
rect 192607 83147 192641 83175
rect 192669 83147 192704 83175
rect 192544 83113 192704 83147
rect 192544 83085 192579 83113
rect 192607 83085 192641 83113
rect 192669 83085 192704 83113
rect 192544 83051 192704 83085
rect 192544 83023 192579 83051
rect 192607 83023 192641 83051
rect 192669 83023 192704 83051
rect 192544 82989 192704 83023
rect 192544 82961 192579 82989
rect 192607 82961 192641 82989
rect 192669 82961 192704 82989
rect 192544 82944 192704 82961
rect 202389 83175 202699 91961
rect 202389 83147 202437 83175
rect 202465 83147 202499 83175
rect 202527 83147 202561 83175
rect 202589 83147 202623 83175
rect 202651 83147 202699 83175
rect 202389 83113 202699 83147
rect 202389 83085 202437 83113
rect 202465 83085 202499 83113
rect 202527 83085 202561 83113
rect 202589 83085 202623 83113
rect 202651 83085 202699 83113
rect 202389 83051 202699 83085
rect 202389 83023 202437 83051
rect 202465 83023 202499 83051
rect 202527 83023 202561 83051
rect 202589 83023 202623 83051
rect 202651 83023 202699 83051
rect 202389 82989 202699 83023
rect 202389 82961 202437 82989
rect 202465 82961 202499 82989
rect 202527 82961 202561 82989
rect 202589 82961 202623 82989
rect 202651 82961 202699 82989
rect 188889 77147 188937 77175
rect 188965 77147 188999 77175
rect 189027 77147 189061 77175
rect 189089 77147 189123 77175
rect 189151 77147 189199 77175
rect 188889 77113 189199 77147
rect 188889 77085 188937 77113
rect 188965 77085 188999 77113
rect 189027 77085 189061 77113
rect 189089 77085 189123 77113
rect 189151 77085 189199 77113
rect 188889 77051 189199 77085
rect 188889 77023 188937 77051
rect 188965 77023 188999 77051
rect 189027 77023 189061 77051
rect 189089 77023 189123 77051
rect 189151 77023 189199 77051
rect 188889 76989 189199 77023
rect 188889 76961 188937 76989
rect 188965 76961 188999 76989
rect 189027 76961 189061 76989
rect 189089 76961 189123 76989
rect 189151 76961 189199 76989
rect 188889 68175 189199 76961
rect 200224 77175 200384 77192
rect 200224 77147 200259 77175
rect 200287 77147 200321 77175
rect 200349 77147 200384 77175
rect 200224 77113 200384 77147
rect 200224 77085 200259 77113
rect 200287 77085 200321 77113
rect 200349 77085 200384 77113
rect 200224 77051 200384 77085
rect 200224 77023 200259 77051
rect 200287 77023 200321 77051
rect 200349 77023 200384 77051
rect 200224 76989 200384 77023
rect 200224 76961 200259 76989
rect 200287 76961 200321 76989
rect 200349 76961 200384 76989
rect 200224 76944 200384 76961
rect 192544 74175 192704 74192
rect 192544 74147 192579 74175
rect 192607 74147 192641 74175
rect 192669 74147 192704 74175
rect 192544 74113 192704 74147
rect 192544 74085 192579 74113
rect 192607 74085 192641 74113
rect 192669 74085 192704 74113
rect 192544 74051 192704 74085
rect 192544 74023 192579 74051
rect 192607 74023 192641 74051
rect 192669 74023 192704 74051
rect 192544 73989 192704 74023
rect 192544 73961 192579 73989
rect 192607 73961 192641 73989
rect 192669 73961 192704 73989
rect 192544 73944 192704 73961
rect 202389 74175 202699 82961
rect 202389 74147 202437 74175
rect 202465 74147 202499 74175
rect 202527 74147 202561 74175
rect 202589 74147 202623 74175
rect 202651 74147 202699 74175
rect 202389 74113 202699 74147
rect 202389 74085 202437 74113
rect 202465 74085 202499 74113
rect 202527 74085 202561 74113
rect 202589 74085 202623 74113
rect 202651 74085 202699 74113
rect 202389 74051 202699 74085
rect 202389 74023 202437 74051
rect 202465 74023 202499 74051
rect 202527 74023 202561 74051
rect 202589 74023 202623 74051
rect 202651 74023 202699 74051
rect 202389 73989 202699 74023
rect 202389 73961 202437 73989
rect 202465 73961 202499 73989
rect 202527 73961 202561 73989
rect 202589 73961 202623 73989
rect 202651 73961 202699 73989
rect 188889 68147 188937 68175
rect 188965 68147 188999 68175
rect 189027 68147 189061 68175
rect 189089 68147 189123 68175
rect 189151 68147 189199 68175
rect 188889 68113 189199 68147
rect 188889 68085 188937 68113
rect 188965 68085 188999 68113
rect 189027 68085 189061 68113
rect 189089 68085 189123 68113
rect 189151 68085 189199 68113
rect 188889 68051 189199 68085
rect 188889 68023 188937 68051
rect 188965 68023 188999 68051
rect 189027 68023 189061 68051
rect 189089 68023 189123 68051
rect 189151 68023 189199 68051
rect 188889 67989 189199 68023
rect 188889 67961 188937 67989
rect 188965 67961 188999 67989
rect 189027 67961 189061 67989
rect 189089 67961 189123 67989
rect 189151 67961 189199 67989
rect 188889 59175 189199 67961
rect 200224 68175 200384 68192
rect 200224 68147 200259 68175
rect 200287 68147 200321 68175
rect 200349 68147 200384 68175
rect 200224 68113 200384 68147
rect 200224 68085 200259 68113
rect 200287 68085 200321 68113
rect 200349 68085 200384 68113
rect 200224 68051 200384 68085
rect 200224 68023 200259 68051
rect 200287 68023 200321 68051
rect 200349 68023 200384 68051
rect 200224 67989 200384 68023
rect 200224 67961 200259 67989
rect 200287 67961 200321 67989
rect 200349 67961 200384 67989
rect 200224 67944 200384 67961
rect 192544 65175 192704 65192
rect 192544 65147 192579 65175
rect 192607 65147 192641 65175
rect 192669 65147 192704 65175
rect 192544 65113 192704 65147
rect 192544 65085 192579 65113
rect 192607 65085 192641 65113
rect 192669 65085 192704 65113
rect 192544 65051 192704 65085
rect 192544 65023 192579 65051
rect 192607 65023 192641 65051
rect 192669 65023 192704 65051
rect 192544 64989 192704 65023
rect 192544 64961 192579 64989
rect 192607 64961 192641 64989
rect 192669 64961 192704 64989
rect 192544 64944 192704 64961
rect 202389 65175 202699 73961
rect 202389 65147 202437 65175
rect 202465 65147 202499 65175
rect 202527 65147 202561 65175
rect 202589 65147 202623 65175
rect 202651 65147 202699 65175
rect 202389 65113 202699 65147
rect 202389 65085 202437 65113
rect 202465 65085 202499 65113
rect 202527 65085 202561 65113
rect 202589 65085 202623 65113
rect 202651 65085 202699 65113
rect 202389 65051 202699 65085
rect 202389 65023 202437 65051
rect 202465 65023 202499 65051
rect 202527 65023 202561 65051
rect 202589 65023 202623 65051
rect 202651 65023 202699 65051
rect 202389 64989 202699 65023
rect 202389 64961 202437 64989
rect 202465 64961 202499 64989
rect 202527 64961 202561 64989
rect 202589 64961 202623 64989
rect 202651 64961 202699 64989
rect 188889 59147 188937 59175
rect 188965 59147 188999 59175
rect 189027 59147 189061 59175
rect 189089 59147 189123 59175
rect 189151 59147 189199 59175
rect 188889 59113 189199 59147
rect 188889 59085 188937 59113
rect 188965 59085 188999 59113
rect 189027 59085 189061 59113
rect 189089 59085 189123 59113
rect 189151 59085 189199 59113
rect 188889 59051 189199 59085
rect 188889 59023 188937 59051
rect 188965 59023 188999 59051
rect 189027 59023 189061 59051
rect 189089 59023 189123 59051
rect 189151 59023 189199 59051
rect 188889 58989 189199 59023
rect 188889 58961 188937 58989
rect 188965 58961 188999 58989
rect 189027 58961 189061 58989
rect 189089 58961 189123 58989
rect 189151 58961 189199 58989
rect 188889 50175 189199 58961
rect 200224 59175 200384 59192
rect 200224 59147 200259 59175
rect 200287 59147 200321 59175
rect 200349 59147 200384 59175
rect 200224 59113 200384 59147
rect 200224 59085 200259 59113
rect 200287 59085 200321 59113
rect 200349 59085 200384 59113
rect 200224 59051 200384 59085
rect 200224 59023 200259 59051
rect 200287 59023 200321 59051
rect 200349 59023 200384 59051
rect 200224 58989 200384 59023
rect 200224 58961 200259 58989
rect 200287 58961 200321 58989
rect 200349 58961 200384 58989
rect 200224 58944 200384 58961
rect 192544 56175 192704 56192
rect 192544 56147 192579 56175
rect 192607 56147 192641 56175
rect 192669 56147 192704 56175
rect 192544 56113 192704 56147
rect 192544 56085 192579 56113
rect 192607 56085 192641 56113
rect 192669 56085 192704 56113
rect 192544 56051 192704 56085
rect 192544 56023 192579 56051
rect 192607 56023 192641 56051
rect 192669 56023 192704 56051
rect 192544 55989 192704 56023
rect 192544 55961 192579 55989
rect 192607 55961 192641 55989
rect 192669 55961 192704 55989
rect 192544 55944 192704 55961
rect 202389 56175 202699 64961
rect 202389 56147 202437 56175
rect 202465 56147 202499 56175
rect 202527 56147 202561 56175
rect 202589 56147 202623 56175
rect 202651 56147 202699 56175
rect 202389 56113 202699 56147
rect 202389 56085 202437 56113
rect 202465 56085 202499 56113
rect 202527 56085 202561 56113
rect 202589 56085 202623 56113
rect 202651 56085 202699 56113
rect 202389 56051 202699 56085
rect 202389 56023 202437 56051
rect 202465 56023 202499 56051
rect 202527 56023 202561 56051
rect 202589 56023 202623 56051
rect 202651 56023 202699 56051
rect 202389 55989 202699 56023
rect 202389 55961 202437 55989
rect 202465 55961 202499 55989
rect 202527 55961 202561 55989
rect 202589 55961 202623 55989
rect 202651 55961 202699 55989
rect 188889 50147 188937 50175
rect 188965 50147 188999 50175
rect 189027 50147 189061 50175
rect 189089 50147 189123 50175
rect 189151 50147 189199 50175
rect 188889 50113 189199 50147
rect 188889 50085 188937 50113
rect 188965 50085 188999 50113
rect 189027 50085 189061 50113
rect 189089 50085 189123 50113
rect 189151 50085 189199 50113
rect 188889 50051 189199 50085
rect 188889 50023 188937 50051
rect 188965 50023 188999 50051
rect 189027 50023 189061 50051
rect 189089 50023 189123 50051
rect 189151 50023 189199 50051
rect 188889 49989 189199 50023
rect 188889 49961 188937 49989
rect 188965 49961 188999 49989
rect 189027 49961 189061 49989
rect 189089 49961 189123 49989
rect 189151 49961 189199 49989
rect 188889 41175 189199 49961
rect 200224 50175 200384 50192
rect 200224 50147 200259 50175
rect 200287 50147 200321 50175
rect 200349 50147 200384 50175
rect 200224 50113 200384 50147
rect 200224 50085 200259 50113
rect 200287 50085 200321 50113
rect 200349 50085 200384 50113
rect 200224 50051 200384 50085
rect 200224 50023 200259 50051
rect 200287 50023 200321 50051
rect 200349 50023 200384 50051
rect 200224 49989 200384 50023
rect 200224 49961 200259 49989
rect 200287 49961 200321 49989
rect 200349 49961 200384 49989
rect 200224 49944 200384 49961
rect 192544 47175 192704 47192
rect 192544 47147 192579 47175
rect 192607 47147 192641 47175
rect 192669 47147 192704 47175
rect 192544 47113 192704 47147
rect 192544 47085 192579 47113
rect 192607 47085 192641 47113
rect 192669 47085 192704 47113
rect 192544 47051 192704 47085
rect 192544 47023 192579 47051
rect 192607 47023 192641 47051
rect 192669 47023 192704 47051
rect 192544 46989 192704 47023
rect 192544 46961 192579 46989
rect 192607 46961 192641 46989
rect 192669 46961 192704 46989
rect 192544 46944 192704 46961
rect 202389 47175 202699 55961
rect 202389 47147 202437 47175
rect 202465 47147 202499 47175
rect 202527 47147 202561 47175
rect 202589 47147 202623 47175
rect 202651 47147 202699 47175
rect 202389 47113 202699 47147
rect 202389 47085 202437 47113
rect 202465 47085 202499 47113
rect 202527 47085 202561 47113
rect 202589 47085 202623 47113
rect 202651 47085 202699 47113
rect 202389 47051 202699 47085
rect 202389 47023 202437 47051
rect 202465 47023 202499 47051
rect 202527 47023 202561 47051
rect 202589 47023 202623 47051
rect 202651 47023 202699 47051
rect 202389 46989 202699 47023
rect 202389 46961 202437 46989
rect 202465 46961 202499 46989
rect 202527 46961 202561 46989
rect 202589 46961 202623 46989
rect 202651 46961 202699 46989
rect 188889 41147 188937 41175
rect 188965 41147 188999 41175
rect 189027 41147 189061 41175
rect 189089 41147 189123 41175
rect 189151 41147 189199 41175
rect 188889 41113 189199 41147
rect 188889 41085 188937 41113
rect 188965 41085 188999 41113
rect 189027 41085 189061 41113
rect 189089 41085 189123 41113
rect 189151 41085 189199 41113
rect 188889 41051 189199 41085
rect 188889 41023 188937 41051
rect 188965 41023 188999 41051
rect 189027 41023 189061 41051
rect 189089 41023 189123 41051
rect 189151 41023 189199 41051
rect 188889 40989 189199 41023
rect 188889 40961 188937 40989
rect 188965 40961 188999 40989
rect 189027 40961 189061 40989
rect 189089 40961 189123 40989
rect 189151 40961 189199 40989
rect 188889 32175 189199 40961
rect 200224 41175 200384 41192
rect 200224 41147 200259 41175
rect 200287 41147 200321 41175
rect 200349 41147 200384 41175
rect 200224 41113 200384 41147
rect 200224 41085 200259 41113
rect 200287 41085 200321 41113
rect 200349 41085 200384 41113
rect 200224 41051 200384 41085
rect 200224 41023 200259 41051
rect 200287 41023 200321 41051
rect 200349 41023 200384 41051
rect 200224 40989 200384 41023
rect 200224 40961 200259 40989
rect 200287 40961 200321 40989
rect 200349 40961 200384 40989
rect 200224 40944 200384 40961
rect 192544 38175 192704 38192
rect 192544 38147 192579 38175
rect 192607 38147 192641 38175
rect 192669 38147 192704 38175
rect 192544 38113 192704 38147
rect 192544 38085 192579 38113
rect 192607 38085 192641 38113
rect 192669 38085 192704 38113
rect 192544 38051 192704 38085
rect 192544 38023 192579 38051
rect 192607 38023 192641 38051
rect 192669 38023 192704 38051
rect 192544 37989 192704 38023
rect 192544 37961 192579 37989
rect 192607 37961 192641 37989
rect 192669 37961 192704 37989
rect 192544 37944 192704 37961
rect 202389 38175 202699 46961
rect 202389 38147 202437 38175
rect 202465 38147 202499 38175
rect 202527 38147 202561 38175
rect 202589 38147 202623 38175
rect 202651 38147 202699 38175
rect 202389 38113 202699 38147
rect 202389 38085 202437 38113
rect 202465 38085 202499 38113
rect 202527 38085 202561 38113
rect 202589 38085 202623 38113
rect 202651 38085 202699 38113
rect 202389 38051 202699 38085
rect 202389 38023 202437 38051
rect 202465 38023 202499 38051
rect 202527 38023 202561 38051
rect 202589 38023 202623 38051
rect 202651 38023 202699 38051
rect 202389 37989 202699 38023
rect 202389 37961 202437 37989
rect 202465 37961 202499 37989
rect 202527 37961 202561 37989
rect 202589 37961 202623 37989
rect 202651 37961 202699 37989
rect 188889 32147 188937 32175
rect 188965 32147 188999 32175
rect 189027 32147 189061 32175
rect 189089 32147 189123 32175
rect 189151 32147 189199 32175
rect 188889 32113 189199 32147
rect 188889 32085 188937 32113
rect 188965 32085 188999 32113
rect 189027 32085 189061 32113
rect 189089 32085 189123 32113
rect 189151 32085 189199 32113
rect 188889 32051 189199 32085
rect 188889 32023 188937 32051
rect 188965 32023 188999 32051
rect 189027 32023 189061 32051
rect 189089 32023 189123 32051
rect 189151 32023 189199 32051
rect 188889 31989 189199 32023
rect 188889 31961 188937 31989
rect 188965 31961 188999 31989
rect 189027 31961 189061 31989
rect 189089 31961 189123 31989
rect 189151 31961 189199 31989
rect 188889 23175 189199 31961
rect 200224 32175 200384 32192
rect 200224 32147 200259 32175
rect 200287 32147 200321 32175
rect 200349 32147 200384 32175
rect 200224 32113 200384 32147
rect 200224 32085 200259 32113
rect 200287 32085 200321 32113
rect 200349 32085 200384 32113
rect 200224 32051 200384 32085
rect 200224 32023 200259 32051
rect 200287 32023 200321 32051
rect 200349 32023 200384 32051
rect 200224 31989 200384 32023
rect 200224 31961 200259 31989
rect 200287 31961 200321 31989
rect 200349 31961 200384 31989
rect 200224 31944 200384 31961
rect 192544 29175 192704 29192
rect 192544 29147 192579 29175
rect 192607 29147 192641 29175
rect 192669 29147 192704 29175
rect 192544 29113 192704 29147
rect 192544 29085 192579 29113
rect 192607 29085 192641 29113
rect 192669 29085 192704 29113
rect 192544 29051 192704 29085
rect 192544 29023 192579 29051
rect 192607 29023 192641 29051
rect 192669 29023 192704 29051
rect 192544 28989 192704 29023
rect 192544 28961 192579 28989
rect 192607 28961 192641 28989
rect 192669 28961 192704 28989
rect 192544 28944 192704 28961
rect 202389 29175 202699 37961
rect 202389 29147 202437 29175
rect 202465 29147 202499 29175
rect 202527 29147 202561 29175
rect 202589 29147 202623 29175
rect 202651 29147 202699 29175
rect 202389 29113 202699 29147
rect 202389 29085 202437 29113
rect 202465 29085 202499 29113
rect 202527 29085 202561 29113
rect 202589 29085 202623 29113
rect 202651 29085 202699 29113
rect 202389 29051 202699 29085
rect 202389 29023 202437 29051
rect 202465 29023 202499 29051
rect 202527 29023 202561 29051
rect 202589 29023 202623 29051
rect 202651 29023 202699 29051
rect 202389 28989 202699 29023
rect 202389 28961 202437 28989
rect 202465 28961 202499 28989
rect 202527 28961 202561 28989
rect 202589 28961 202623 28989
rect 202651 28961 202699 28989
rect 188889 23147 188937 23175
rect 188965 23147 188999 23175
rect 189027 23147 189061 23175
rect 189089 23147 189123 23175
rect 189151 23147 189199 23175
rect 188889 23113 189199 23147
rect 188889 23085 188937 23113
rect 188965 23085 188999 23113
rect 189027 23085 189061 23113
rect 189089 23085 189123 23113
rect 189151 23085 189199 23113
rect 188889 23051 189199 23085
rect 188889 23023 188937 23051
rect 188965 23023 188999 23051
rect 189027 23023 189061 23051
rect 189089 23023 189123 23051
rect 189151 23023 189199 23051
rect 188889 22989 189199 23023
rect 188889 22961 188937 22989
rect 188965 22961 188999 22989
rect 189027 22961 189061 22989
rect 189089 22961 189123 22989
rect 189151 22961 189199 22989
rect 188889 14175 189199 22961
rect 200224 23175 200384 23192
rect 200224 23147 200259 23175
rect 200287 23147 200321 23175
rect 200349 23147 200384 23175
rect 200224 23113 200384 23147
rect 200224 23085 200259 23113
rect 200287 23085 200321 23113
rect 200349 23085 200384 23113
rect 200224 23051 200384 23085
rect 200224 23023 200259 23051
rect 200287 23023 200321 23051
rect 200349 23023 200384 23051
rect 200224 22989 200384 23023
rect 200224 22961 200259 22989
rect 200287 22961 200321 22989
rect 200349 22961 200384 22989
rect 200224 22944 200384 22961
rect 192544 20175 192704 20192
rect 192544 20147 192579 20175
rect 192607 20147 192641 20175
rect 192669 20147 192704 20175
rect 192544 20113 192704 20147
rect 192544 20085 192579 20113
rect 192607 20085 192641 20113
rect 192669 20085 192704 20113
rect 192544 20051 192704 20085
rect 192544 20023 192579 20051
rect 192607 20023 192641 20051
rect 192669 20023 192704 20051
rect 192544 19989 192704 20023
rect 192544 19961 192579 19989
rect 192607 19961 192641 19989
rect 192669 19961 192704 19989
rect 192544 19944 192704 19961
rect 202389 20175 202699 28961
rect 202389 20147 202437 20175
rect 202465 20147 202499 20175
rect 202527 20147 202561 20175
rect 202589 20147 202623 20175
rect 202651 20147 202699 20175
rect 202389 20113 202699 20147
rect 202389 20085 202437 20113
rect 202465 20085 202499 20113
rect 202527 20085 202561 20113
rect 202589 20085 202623 20113
rect 202651 20085 202699 20113
rect 202389 20051 202699 20085
rect 202389 20023 202437 20051
rect 202465 20023 202499 20051
rect 202527 20023 202561 20051
rect 202589 20023 202623 20051
rect 202651 20023 202699 20051
rect 202389 19989 202699 20023
rect 202389 19961 202437 19989
rect 202465 19961 202499 19989
rect 202527 19961 202561 19989
rect 202589 19961 202623 19989
rect 202651 19961 202699 19989
rect 188889 14147 188937 14175
rect 188965 14147 188999 14175
rect 189027 14147 189061 14175
rect 189089 14147 189123 14175
rect 189151 14147 189199 14175
rect 188889 14113 189199 14147
rect 188889 14085 188937 14113
rect 188965 14085 188999 14113
rect 189027 14085 189061 14113
rect 189089 14085 189123 14113
rect 189151 14085 189199 14113
rect 188889 14051 189199 14085
rect 188889 14023 188937 14051
rect 188965 14023 188999 14051
rect 189027 14023 189061 14051
rect 189089 14023 189123 14051
rect 189151 14023 189199 14051
rect 188889 13989 189199 14023
rect 188889 13961 188937 13989
rect 188965 13961 188999 13989
rect 189027 13961 189061 13989
rect 189089 13961 189123 13989
rect 189151 13961 189199 13989
rect 188889 5175 189199 13961
rect 200224 14175 200384 14192
rect 200224 14147 200259 14175
rect 200287 14147 200321 14175
rect 200349 14147 200384 14175
rect 200224 14113 200384 14147
rect 200224 14085 200259 14113
rect 200287 14085 200321 14113
rect 200349 14085 200384 14113
rect 200224 14051 200384 14085
rect 200224 14023 200259 14051
rect 200287 14023 200321 14051
rect 200349 14023 200384 14051
rect 200224 13989 200384 14023
rect 200224 13961 200259 13989
rect 200287 13961 200321 13989
rect 200349 13961 200384 13989
rect 200224 13944 200384 13961
rect 192544 11175 192704 11192
rect 192544 11147 192579 11175
rect 192607 11147 192641 11175
rect 192669 11147 192704 11175
rect 192544 11113 192704 11147
rect 192544 11085 192579 11113
rect 192607 11085 192641 11113
rect 192669 11085 192704 11113
rect 192544 11051 192704 11085
rect 192544 11023 192579 11051
rect 192607 11023 192641 11051
rect 192669 11023 192704 11051
rect 192544 10989 192704 11023
rect 192544 10961 192579 10989
rect 192607 10961 192641 10989
rect 192669 10961 192704 10989
rect 192544 10944 192704 10961
rect 202389 11175 202699 19961
rect 202389 11147 202437 11175
rect 202465 11147 202499 11175
rect 202527 11147 202561 11175
rect 202589 11147 202623 11175
rect 202651 11147 202699 11175
rect 202389 11113 202699 11147
rect 202389 11085 202437 11113
rect 202465 11085 202499 11113
rect 202527 11085 202561 11113
rect 202589 11085 202623 11113
rect 202651 11085 202699 11113
rect 202389 11051 202699 11085
rect 202389 11023 202437 11051
rect 202465 11023 202499 11051
rect 202527 11023 202561 11051
rect 202589 11023 202623 11051
rect 202651 11023 202699 11051
rect 202389 10989 202699 11023
rect 202389 10961 202437 10989
rect 202465 10961 202499 10989
rect 202527 10961 202561 10989
rect 202589 10961 202623 10989
rect 202651 10961 202699 10989
rect 188889 5147 188937 5175
rect 188965 5147 188999 5175
rect 189027 5147 189061 5175
rect 189089 5147 189123 5175
rect 189151 5147 189199 5175
rect 188889 5113 189199 5147
rect 188889 5085 188937 5113
rect 188965 5085 188999 5113
rect 189027 5085 189061 5113
rect 189089 5085 189123 5113
rect 189151 5085 189199 5113
rect 188889 5051 189199 5085
rect 188889 5023 188937 5051
rect 188965 5023 188999 5051
rect 189027 5023 189061 5051
rect 189089 5023 189123 5051
rect 189151 5023 189199 5051
rect 188889 4989 189199 5023
rect 188889 4961 188937 4989
rect 188965 4961 188999 4989
rect 189027 4961 189061 4989
rect 189089 4961 189123 4989
rect 189151 4961 189199 4989
rect 188889 -560 189199 4961
rect 200224 5175 200384 5192
rect 200224 5147 200259 5175
rect 200287 5147 200321 5175
rect 200349 5147 200384 5175
rect 200224 5113 200384 5147
rect 200224 5085 200259 5113
rect 200287 5085 200321 5113
rect 200349 5085 200384 5113
rect 200224 5051 200384 5085
rect 200224 5023 200259 5051
rect 200287 5023 200321 5051
rect 200349 5023 200384 5051
rect 200224 4989 200384 5023
rect 200224 4961 200259 4989
rect 200287 4961 200321 4989
rect 200349 4961 200384 4989
rect 200224 4944 200384 4961
rect 188889 -588 188937 -560
rect 188965 -588 188999 -560
rect 189027 -588 189061 -560
rect 189089 -588 189123 -560
rect 189151 -588 189199 -560
rect 188889 -622 189199 -588
rect 188889 -650 188937 -622
rect 188965 -650 188999 -622
rect 189027 -650 189061 -622
rect 189089 -650 189123 -622
rect 189151 -650 189199 -622
rect 188889 -684 189199 -650
rect 188889 -712 188937 -684
rect 188965 -712 188999 -684
rect 189027 -712 189061 -684
rect 189089 -712 189123 -684
rect 189151 -712 189199 -684
rect 188889 -746 189199 -712
rect 188889 -774 188937 -746
rect 188965 -774 188999 -746
rect 189027 -774 189061 -746
rect 189089 -774 189123 -746
rect 189151 -774 189199 -746
rect 188889 -822 189199 -774
rect 202389 2175 202699 10961
rect 202389 2147 202437 2175
rect 202465 2147 202499 2175
rect 202527 2147 202561 2175
rect 202589 2147 202623 2175
rect 202651 2147 202699 2175
rect 202389 2113 202699 2147
rect 202389 2085 202437 2113
rect 202465 2085 202499 2113
rect 202527 2085 202561 2113
rect 202589 2085 202623 2113
rect 202651 2085 202699 2113
rect 202389 2051 202699 2085
rect 202389 2023 202437 2051
rect 202465 2023 202499 2051
rect 202527 2023 202561 2051
rect 202589 2023 202623 2051
rect 202651 2023 202699 2051
rect 202389 1989 202699 2023
rect 202389 1961 202437 1989
rect 202465 1961 202499 1989
rect 202527 1961 202561 1989
rect 202589 1961 202623 1989
rect 202651 1961 202699 1989
rect 202389 -80 202699 1961
rect 202389 -108 202437 -80
rect 202465 -108 202499 -80
rect 202527 -108 202561 -80
rect 202589 -108 202623 -80
rect 202651 -108 202699 -80
rect 202389 -142 202699 -108
rect 202389 -170 202437 -142
rect 202465 -170 202499 -142
rect 202527 -170 202561 -142
rect 202589 -170 202623 -142
rect 202651 -170 202699 -142
rect 202389 -204 202699 -170
rect 202389 -232 202437 -204
rect 202465 -232 202499 -204
rect 202527 -232 202561 -204
rect 202589 -232 202623 -204
rect 202651 -232 202699 -204
rect 202389 -266 202699 -232
rect 202389 -294 202437 -266
rect 202465 -294 202499 -266
rect 202527 -294 202561 -266
rect 202589 -294 202623 -266
rect 202651 -294 202699 -266
rect 202389 -822 202699 -294
rect 204249 299086 204559 299134
rect 204249 299058 204297 299086
rect 204325 299058 204359 299086
rect 204387 299058 204421 299086
rect 204449 299058 204483 299086
rect 204511 299058 204559 299086
rect 204249 299024 204559 299058
rect 204249 298996 204297 299024
rect 204325 298996 204359 299024
rect 204387 298996 204421 299024
rect 204449 298996 204483 299024
rect 204511 298996 204559 299024
rect 204249 298962 204559 298996
rect 204249 298934 204297 298962
rect 204325 298934 204359 298962
rect 204387 298934 204421 298962
rect 204449 298934 204483 298962
rect 204511 298934 204559 298962
rect 204249 298900 204559 298934
rect 204249 298872 204297 298900
rect 204325 298872 204359 298900
rect 204387 298872 204421 298900
rect 204449 298872 204483 298900
rect 204511 298872 204559 298900
rect 204249 293175 204559 298872
rect 204249 293147 204297 293175
rect 204325 293147 204359 293175
rect 204387 293147 204421 293175
rect 204449 293147 204483 293175
rect 204511 293147 204559 293175
rect 204249 293113 204559 293147
rect 204249 293085 204297 293113
rect 204325 293085 204359 293113
rect 204387 293085 204421 293113
rect 204449 293085 204483 293113
rect 204511 293085 204559 293113
rect 204249 293051 204559 293085
rect 204249 293023 204297 293051
rect 204325 293023 204359 293051
rect 204387 293023 204421 293051
rect 204449 293023 204483 293051
rect 204511 293023 204559 293051
rect 204249 292989 204559 293023
rect 204249 292961 204297 292989
rect 204325 292961 204359 292989
rect 204387 292961 204421 292989
rect 204449 292961 204483 292989
rect 204511 292961 204559 292989
rect 204249 284175 204559 292961
rect 204249 284147 204297 284175
rect 204325 284147 204359 284175
rect 204387 284147 204421 284175
rect 204449 284147 204483 284175
rect 204511 284147 204559 284175
rect 204249 284113 204559 284147
rect 204249 284085 204297 284113
rect 204325 284085 204359 284113
rect 204387 284085 204421 284113
rect 204449 284085 204483 284113
rect 204511 284085 204559 284113
rect 204249 284051 204559 284085
rect 204249 284023 204297 284051
rect 204325 284023 204359 284051
rect 204387 284023 204421 284051
rect 204449 284023 204483 284051
rect 204511 284023 204559 284051
rect 204249 283989 204559 284023
rect 204249 283961 204297 283989
rect 204325 283961 204359 283989
rect 204387 283961 204421 283989
rect 204449 283961 204483 283989
rect 204511 283961 204559 283989
rect 204249 275175 204559 283961
rect 204249 275147 204297 275175
rect 204325 275147 204359 275175
rect 204387 275147 204421 275175
rect 204449 275147 204483 275175
rect 204511 275147 204559 275175
rect 204249 275113 204559 275147
rect 204249 275085 204297 275113
rect 204325 275085 204359 275113
rect 204387 275085 204421 275113
rect 204449 275085 204483 275113
rect 204511 275085 204559 275113
rect 204249 275051 204559 275085
rect 204249 275023 204297 275051
rect 204325 275023 204359 275051
rect 204387 275023 204421 275051
rect 204449 275023 204483 275051
rect 204511 275023 204559 275051
rect 204249 274989 204559 275023
rect 204249 274961 204297 274989
rect 204325 274961 204359 274989
rect 204387 274961 204421 274989
rect 204449 274961 204483 274989
rect 204511 274961 204559 274989
rect 204249 266175 204559 274961
rect 204249 266147 204297 266175
rect 204325 266147 204359 266175
rect 204387 266147 204421 266175
rect 204449 266147 204483 266175
rect 204511 266147 204559 266175
rect 204249 266113 204559 266147
rect 204249 266085 204297 266113
rect 204325 266085 204359 266113
rect 204387 266085 204421 266113
rect 204449 266085 204483 266113
rect 204511 266085 204559 266113
rect 204249 266051 204559 266085
rect 204249 266023 204297 266051
rect 204325 266023 204359 266051
rect 204387 266023 204421 266051
rect 204449 266023 204483 266051
rect 204511 266023 204559 266051
rect 204249 265989 204559 266023
rect 204249 265961 204297 265989
rect 204325 265961 204359 265989
rect 204387 265961 204421 265989
rect 204449 265961 204483 265989
rect 204511 265961 204559 265989
rect 204249 257175 204559 265961
rect 204249 257147 204297 257175
rect 204325 257147 204359 257175
rect 204387 257147 204421 257175
rect 204449 257147 204483 257175
rect 204511 257147 204559 257175
rect 204249 257113 204559 257147
rect 204249 257085 204297 257113
rect 204325 257085 204359 257113
rect 204387 257085 204421 257113
rect 204449 257085 204483 257113
rect 204511 257085 204559 257113
rect 204249 257051 204559 257085
rect 204249 257023 204297 257051
rect 204325 257023 204359 257051
rect 204387 257023 204421 257051
rect 204449 257023 204483 257051
rect 204511 257023 204559 257051
rect 204249 256989 204559 257023
rect 204249 256961 204297 256989
rect 204325 256961 204359 256989
rect 204387 256961 204421 256989
rect 204449 256961 204483 256989
rect 204511 256961 204559 256989
rect 204249 248175 204559 256961
rect 204249 248147 204297 248175
rect 204325 248147 204359 248175
rect 204387 248147 204421 248175
rect 204449 248147 204483 248175
rect 204511 248147 204559 248175
rect 204249 248113 204559 248147
rect 204249 248085 204297 248113
rect 204325 248085 204359 248113
rect 204387 248085 204421 248113
rect 204449 248085 204483 248113
rect 204511 248085 204559 248113
rect 204249 248051 204559 248085
rect 204249 248023 204297 248051
rect 204325 248023 204359 248051
rect 204387 248023 204421 248051
rect 204449 248023 204483 248051
rect 204511 248023 204559 248051
rect 204249 247989 204559 248023
rect 204249 247961 204297 247989
rect 204325 247961 204359 247989
rect 204387 247961 204421 247989
rect 204449 247961 204483 247989
rect 204511 247961 204559 247989
rect 204249 239175 204559 247961
rect 204249 239147 204297 239175
rect 204325 239147 204359 239175
rect 204387 239147 204421 239175
rect 204449 239147 204483 239175
rect 204511 239147 204559 239175
rect 204249 239113 204559 239147
rect 204249 239085 204297 239113
rect 204325 239085 204359 239113
rect 204387 239085 204421 239113
rect 204449 239085 204483 239113
rect 204511 239085 204559 239113
rect 204249 239051 204559 239085
rect 204249 239023 204297 239051
rect 204325 239023 204359 239051
rect 204387 239023 204421 239051
rect 204449 239023 204483 239051
rect 204511 239023 204559 239051
rect 204249 238989 204559 239023
rect 204249 238961 204297 238989
rect 204325 238961 204359 238989
rect 204387 238961 204421 238989
rect 204449 238961 204483 238989
rect 204511 238961 204559 238989
rect 204249 230175 204559 238961
rect 204249 230147 204297 230175
rect 204325 230147 204359 230175
rect 204387 230147 204421 230175
rect 204449 230147 204483 230175
rect 204511 230147 204559 230175
rect 204249 230113 204559 230147
rect 204249 230085 204297 230113
rect 204325 230085 204359 230113
rect 204387 230085 204421 230113
rect 204449 230085 204483 230113
rect 204511 230085 204559 230113
rect 204249 230051 204559 230085
rect 204249 230023 204297 230051
rect 204325 230023 204359 230051
rect 204387 230023 204421 230051
rect 204449 230023 204483 230051
rect 204511 230023 204559 230051
rect 204249 229989 204559 230023
rect 204249 229961 204297 229989
rect 204325 229961 204359 229989
rect 204387 229961 204421 229989
rect 204449 229961 204483 229989
rect 204511 229961 204559 229989
rect 204249 221175 204559 229961
rect 204249 221147 204297 221175
rect 204325 221147 204359 221175
rect 204387 221147 204421 221175
rect 204449 221147 204483 221175
rect 204511 221147 204559 221175
rect 204249 221113 204559 221147
rect 204249 221085 204297 221113
rect 204325 221085 204359 221113
rect 204387 221085 204421 221113
rect 204449 221085 204483 221113
rect 204511 221085 204559 221113
rect 204249 221051 204559 221085
rect 204249 221023 204297 221051
rect 204325 221023 204359 221051
rect 204387 221023 204421 221051
rect 204449 221023 204483 221051
rect 204511 221023 204559 221051
rect 204249 220989 204559 221023
rect 204249 220961 204297 220989
rect 204325 220961 204359 220989
rect 204387 220961 204421 220989
rect 204449 220961 204483 220989
rect 204511 220961 204559 220989
rect 204249 212175 204559 220961
rect 204249 212147 204297 212175
rect 204325 212147 204359 212175
rect 204387 212147 204421 212175
rect 204449 212147 204483 212175
rect 204511 212147 204559 212175
rect 204249 212113 204559 212147
rect 204249 212085 204297 212113
rect 204325 212085 204359 212113
rect 204387 212085 204421 212113
rect 204449 212085 204483 212113
rect 204511 212085 204559 212113
rect 204249 212051 204559 212085
rect 204249 212023 204297 212051
rect 204325 212023 204359 212051
rect 204387 212023 204421 212051
rect 204449 212023 204483 212051
rect 204511 212023 204559 212051
rect 204249 211989 204559 212023
rect 204249 211961 204297 211989
rect 204325 211961 204359 211989
rect 204387 211961 204421 211989
rect 204449 211961 204483 211989
rect 204511 211961 204559 211989
rect 204249 203175 204559 211961
rect 204249 203147 204297 203175
rect 204325 203147 204359 203175
rect 204387 203147 204421 203175
rect 204449 203147 204483 203175
rect 204511 203147 204559 203175
rect 204249 203113 204559 203147
rect 204249 203085 204297 203113
rect 204325 203085 204359 203113
rect 204387 203085 204421 203113
rect 204449 203085 204483 203113
rect 204511 203085 204559 203113
rect 204249 203051 204559 203085
rect 204249 203023 204297 203051
rect 204325 203023 204359 203051
rect 204387 203023 204421 203051
rect 204449 203023 204483 203051
rect 204511 203023 204559 203051
rect 204249 202989 204559 203023
rect 204249 202961 204297 202989
rect 204325 202961 204359 202989
rect 204387 202961 204421 202989
rect 204449 202961 204483 202989
rect 204511 202961 204559 202989
rect 204249 194175 204559 202961
rect 204249 194147 204297 194175
rect 204325 194147 204359 194175
rect 204387 194147 204421 194175
rect 204449 194147 204483 194175
rect 204511 194147 204559 194175
rect 204249 194113 204559 194147
rect 204249 194085 204297 194113
rect 204325 194085 204359 194113
rect 204387 194085 204421 194113
rect 204449 194085 204483 194113
rect 204511 194085 204559 194113
rect 204249 194051 204559 194085
rect 204249 194023 204297 194051
rect 204325 194023 204359 194051
rect 204387 194023 204421 194051
rect 204449 194023 204483 194051
rect 204511 194023 204559 194051
rect 204249 193989 204559 194023
rect 204249 193961 204297 193989
rect 204325 193961 204359 193989
rect 204387 193961 204421 193989
rect 204449 193961 204483 193989
rect 204511 193961 204559 193989
rect 204249 185175 204559 193961
rect 204249 185147 204297 185175
rect 204325 185147 204359 185175
rect 204387 185147 204421 185175
rect 204449 185147 204483 185175
rect 204511 185147 204559 185175
rect 204249 185113 204559 185147
rect 204249 185085 204297 185113
rect 204325 185085 204359 185113
rect 204387 185085 204421 185113
rect 204449 185085 204483 185113
rect 204511 185085 204559 185113
rect 204249 185051 204559 185085
rect 204249 185023 204297 185051
rect 204325 185023 204359 185051
rect 204387 185023 204421 185051
rect 204449 185023 204483 185051
rect 204511 185023 204559 185051
rect 204249 184989 204559 185023
rect 204249 184961 204297 184989
rect 204325 184961 204359 184989
rect 204387 184961 204421 184989
rect 204449 184961 204483 184989
rect 204511 184961 204559 184989
rect 204249 176175 204559 184961
rect 204249 176147 204297 176175
rect 204325 176147 204359 176175
rect 204387 176147 204421 176175
rect 204449 176147 204483 176175
rect 204511 176147 204559 176175
rect 204249 176113 204559 176147
rect 204249 176085 204297 176113
rect 204325 176085 204359 176113
rect 204387 176085 204421 176113
rect 204449 176085 204483 176113
rect 204511 176085 204559 176113
rect 204249 176051 204559 176085
rect 204249 176023 204297 176051
rect 204325 176023 204359 176051
rect 204387 176023 204421 176051
rect 204449 176023 204483 176051
rect 204511 176023 204559 176051
rect 204249 175989 204559 176023
rect 204249 175961 204297 175989
rect 204325 175961 204359 175989
rect 204387 175961 204421 175989
rect 204449 175961 204483 175989
rect 204511 175961 204559 175989
rect 204249 167175 204559 175961
rect 217749 298606 218059 299134
rect 217749 298578 217797 298606
rect 217825 298578 217859 298606
rect 217887 298578 217921 298606
rect 217949 298578 217983 298606
rect 218011 298578 218059 298606
rect 217749 298544 218059 298578
rect 217749 298516 217797 298544
rect 217825 298516 217859 298544
rect 217887 298516 217921 298544
rect 217949 298516 217983 298544
rect 218011 298516 218059 298544
rect 217749 298482 218059 298516
rect 217749 298454 217797 298482
rect 217825 298454 217859 298482
rect 217887 298454 217921 298482
rect 217949 298454 217983 298482
rect 218011 298454 218059 298482
rect 217749 298420 218059 298454
rect 217749 298392 217797 298420
rect 217825 298392 217859 298420
rect 217887 298392 217921 298420
rect 217949 298392 217983 298420
rect 218011 298392 218059 298420
rect 217749 290175 218059 298392
rect 217749 290147 217797 290175
rect 217825 290147 217859 290175
rect 217887 290147 217921 290175
rect 217949 290147 217983 290175
rect 218011 290147 218059 290175
rect 217749 290113 218059 290147
rect 217749 290085 217797 290113
rect 217825 290085 217859 290113
rect 217887 290085 217921 290113
rect 217949 290085 217983 290113
rect 218011 290085 218059 290113
rect 217749 290051 218059 290085
rect 217749 290023 217797 290051
rect 217825 290023 217859 290051
rect 217887 290023 217921 290051
rect 217949 290023 217983 290051
rect 218011 290023 218059 290051
rect 217749 289989 218059 290023
rect 217749 289961 217797 289989
rect 217825 289961 217859 289989
rect 217887 289961 217921 289989
rect 217949 289961 217983 289989
rect 218011 289961 218059 289989
rect 217749 281175 218059 289961
rect 217749 281147 217797 281175
rect 217825 281147 217859 281175
rect 217887 281147 217921 281175
rect 217949 281147 217983 281175
rect 218011 281147 218059 281175
rect 217749 281113 218059 281147
rect 217749 281085 217797 281113
rect 217825 281085 217859 281113
rect 217887 281085 217921 281113
rect 217949 281085 217983 281113
rect 218011 281085 218059 281113
rect 217749 281051 218059 281085
rect 217749 281023 217797 281051
rect 217825 281023 217859 281051
rect 217887 281023 217921 281051
rect 217949 281023 217983 281051
rect 218011 281023 218059 281051
rect 217749 280989 218059 281023
rect 217749 280961 217797 280989
rect 217825 280961 217859 280989
rect 217887 280961 217921 280989
rect 217949 280961 217983 280989
rect 218011 280961 218059 280989
rect 217749 272175 218059 280961
rect 217749 272147 217797 272175
rect 217825 272147 217859 272175
rect 217887 272147 217921 272175
rect 217949 272147 217983 272175
rect 218011 272147 218059 272175
rect 217749 272113 218059 272147
rect 217749 272085 217797 272113
rect 217825 272085 217859 272113
rect 217887 272085 217921 272113
rect 217949 272085 217983 272113
rect 218011 272085 218059 272113
rect 217749 272051 218059 272085
rect 217749 272023 217797 272051
rect 217825 272023 217859 272051
rect 217887 272023 217921 272051
rect 217949 272023 217983 272051
rect 218011 272023 218059 272051
rect 217749 271989 218059 272023
rect 217749 271961 217797 271989
rect 217825 271961 217859 271989
rect 217887 271961 217921 271989
rect 217949 271961 217983 271989
rect 218011 271961 218059 271989
rect 217749 263175 218059 271961
rect 217749 263147 217797 263175
rect 217825 263147 217859 263175
rect 217887 263147 217921 263175
rect 217949 263147 217983 263175
rect 218011 263147 218059 263175
rect 217749 263113 218059 263147
rect 217749 263085 217797 263113
rect 217825 263085 217859 263113
rect 217887 263085 217921 263113
rect 217949 263085 217983 263113
rect 218011 263085 218059 263113
rect 217749 263051 218059 263085
rect 217749 263023 217797 263051
rect 217825 263023 217859 263051
rect 217887 263023 217921 263051
rect 217949 263023 217983 263051
rect 218011 263023 218059 263051
rect 217749 262989 218059 263023
rect 217749 262961 217797 262989
rect 217825 262961 217859 262989
rect 217887 262961 217921 262989
rect 217949 262961 217983 262989
rect 218011 262961 218059 262989
rect 217749 254175 218059 262961
rect 217749 254147 217797 254175
rect 217825 254147 217859 254175
rect 217887 254147 217921 254175
rect 217949 254147 217983 254175
rect 218011 254147 218059 254175
rect 217749 254113 218059 254147
rect 217749 254085 217797 254113
rect 217825 254085 217859 254113
rect 217887 254085 217921 254113
rect 217949 254085 217983 254113
rect 218011 254085 218059 254113
rect 217749 254051 218059 254085
rect 217749 254023 217797 254051
rect 217825 254023 217859 254051
rect 217887 254023 217921 254051
rect 217949 254023 217983 254051
rect 218011 254023 218059 254051
rect 217749 253989 218059 254023
rect 217749 253961 217797 253989
rect 217825 253961 217859 253989
rect 217887 253961 217921 253989
rect 217949 253961 217983 253989
rect 218011 253961 218059 253989
rect 217749 245175 218059 253961
rect 217749 245147 217797 245175
rect 217825 245147 217859 245175
rect 217887 245147 217921 245175
rect 217949 245147 217983 245175
rect 218011 245147 218059 245175
rect 217749 245113 218059 245147
rect 217749 245085 217797 245113
rect 217825 245085 217859 245113
rect 217887 245085 217921 245113
rect 217949 245085 217983 245113
rect 218011 245085 218059 245113
rect 217749 245051 218059 245085
rect 217749 245023 217797 245051
rect 217825 245023 217859 245051
rect 217887 245023 217921 245051
rect 217949 245023 217983 245051
rect 218011 245023 218059 245051
rect 217749 244989 218059 245023
rect 217749 244961 217797 244989
rect 217825 244961 217859 244989
rect 217887 244961 217921 244989
rect 217949 244961 217983 244989
rect 218011 244961 218059 244989
rect 217749 236175 218059 244961
rect 217749 236147 217797 236175
rect 217825 236147 217859 236175
rect 217887 236147 217921 236175
rect 217949 236147 217983 236175
rect 218011 236147 218059 236175
rect 217749 236113 218059 236147
rect 217749 236085 217797 236113
rect 217825 236085 217859 236113
rect 217887 236085 217921 236113
rect 217949 236085 217983 236113
rect 218011 236085 218059 236113
rect 217749 236051 218059 236085
rect 217749 236023 217797 236051
rect 217825 236023 217859 236051
rect 217887 236023 217921 236051
rect 217949 236023 217983 236051
rect 218011 236023 218059 236051
rect 217749 235989 218059 236023
rect 217749 235961 217797 235989
rect 217825 235961 217859 235989
rect 217887 235961 217921 235989
rect 217949 235961 217983 235989
rect 218011 235961 218059 235989
rect 217749 227175 218059 235961
rect 217749 227147 217797 227175
rect 217825 227147 217859 227175
rect 217887 227147 217921 227175
rect 217949 227147 217983 227175
rect 218011 227147 218059 227175
rect 217749 227113 218059 227147
rect 217749 227085 217797 227113
rect 217825 227085 217859 227113
rect 217887 227085 217921 227113
rect 217949 227085 217983 227113
rect 218011 227085 218059 227113
rect 217749 227051 218059 227085
rect 217749 227023 217797 227051
rect 217825 227023 217859 227051
rect 217887 227023 217921 227051
rect 217949 227023 217983 227051
rect 218011 227023 218059 227051
rect 217749 226989 218059 227023
rect 217749 226961 217797 226989
rect 217825 226961 217859 226989
rect 217887 226961 217921 226989
rect 217949 226961 217983 226989
rect 218011 226961 218059 226989
rect 217749 218175 218059 226961
rect 217749 218147 217797 218175
rect 217825 218147 217859 218175
rect 217887 218147 217921 218175
rect 217949 218147 217983 218175
rect 218011 218147 218059 218175
rect 217749 218113 218059 218147
rect 217749 218085 217797 218113
rect 217825 218085 217859 218113
rect 217887 218085 217921 218113
rect 217949 218085 217983 218113
rect 218011 218085 218059 218113
rect 217749 218051 218059 218085
rect 217749 218023 217797 218051
rect 217825 218023 217859 218051
rect 217887 218023 217921 218051
rect 217949 218023 217983 218051
rect 218011 218023 218059 218051
rect 217749 217989 218059 218023
rect 217749 217961 217797 217989
rect 217825 217961 217859 217989
rect 217887 217961 217921 217989
rect 217949 217961 217983 217989
rect 218011 217961 218059 217989
rect 217749 209175 218059 217961
rect 217749 209147 217797 209175
rect 217825 209147 217859 209175
rect 217887 209147 217921 209175
rect 217949 209147 217983 209175
rect 218011 209147 218059 209175
rect 217749 209113 218059 209147
rect 217749 209085 217797 209113
rect 217825 209085 217859 209113
rect 217887 209085 217921 209113
rect 217949 209085 217983 209113
rect 218011 209085 218059 209113
rect 217749 209051 218059 209085
rect 217749 209023 217797 209051
rect 217825 209023 217859 209051
rect 217887 209023 217921 209051
rect 217949 209023 217983 209051
rect 218011 209023 218059 209051
rect 217749 208989 218059 209023
rect 217749 208961 217797 208989
rect 217825 208961 217859 208989
rect 217887 208961 217921 208989
rect 217949 208961 217983 208989
rect 218011 208961 218059 208989
rect 217749 200175 218059 208961
rect 217749 200147 217797 200175
rect 217825 200147 217859 200175
rect 217887 200147 217921 200175
rect 217949 200147 217983 200175
rect 218011 200147 218059 200175
rect 217749 200113 218059 200147
rect 217749 200085 217797 200113
rect 217825 200085 217859 200113
rect 217887 200085 217921 200113
rect 217949 200085 217983 200113
rect 218011 200085 218059 200113
rect 217749 200051 218059 200085
rect 217749 200023 217797 200051
rect 217825 200023 217859 200051
rect 217887 200023 217921 200051
rect 217949 200023 217983 200051
rect 218011 200023 218059 200051
rect 217749 199989 218059 200023
rect 217749 199961 217797 199989
rect 217825 199961 217859 199989
rect 217887 199961 217921 199989
rect 217949 199961 217983 199989
rect 218011 199961 218059 199989
rect 217749 191175 218059 199961
rect 217749 191147 217797 191175
rect 217825 191147 217859 191175
rect 217887 191147 217921 191175
rect 217949 191147 217983 191175
rect 218011 191147 218059 191175
rect 217749 191113 218059 191147
rect 217749 191085 217797 191113
rect 217825 191085 217859 191113
rect 217887 191085 217921 191113
rect 217949 191085 217983 191113
rect 218011 191085 218059 191113
rect 217749 191051 218059 191085
rect 217749 191023 217797 191051
rect 217825 191023 217859 191051
rect 217887 191023 217921 191051
rect 217949 191023 217983 191051
rect 218011 191023 218059 191051
rect 217749 190989 218059 191023
rect 217749 190961 217797 190989
rect 217825 190961 217859 190989
rect 217887 190961 217921 190989
rect 217949 190961 217983 190989
rect 218011 190961 218059 190989
rect 217749 182175 218059 190961
rect 217749 182147 217797 182175
rect 217825 182147 217859 182175
rect 217887 182147 217921 182175
rect 217949 182147 217983 182175
rect 218011 182147 218059 182175
rect 217749 182113 218059 182147
rect 217749 182085 217797 182113
rect 217825 182085 217859 182113
rect 217887 182085 217921 182113
rect 217949 182085 217983 182113
rect 218011 182085 218059 182113
rect 217749 182051 218059 182085
rect 217749 182023 217797 182051
rect 217825 182023 217859 182051
rect 217887 182023 217921 182051
rect 217949 182023 217983 182051
rect 218011 182023 218059 182051
rect 217749 181989 218059 182023
rect 217749 181961 217797 181989
rect 217825 181961 217859 181989
rect 217887 181961 217921 181989
rect 217949 181961 217983 181989
rect 218011 181961 218059 181989
rect 207904 173175 208064 173192
rect 207904 173147 207939 173175
rect 207967 173147 208001 173175
rect 208029 173147 208064 173175
rect 207904 173113 208064 173147
rect 207904 173085 207939 173113
rect 207967 173085 208001 173113
rect 208029 173085 208064 173113
rect 207904 173051 208064 173085
rect 207904 173023 207939 173051
rect 207967 173023 208001 173051
rect 208029 173023 208064 173051
rect 207904 172989 208064 173023
rect 207904 172961 207939 172989
rect 207967 172961 208001 172989
rect 208029 172961 208064 172989
rect 207904 172944 208064 172961
rect 217749 173175 218059 181961
rect 217749 173147 217797 173175
rect 217825 173147 217859 173175
rect 217887 173147 217921 173175
rect 217949 173147 217983 173175
rect 218011 173147 218059 173175
rect 217749 173113 218059 173147
rect 217749 173085 217797 173113
rect 217825 173085 217859 173113
rect 217887 173085 217921 173113
rect 217949 173085 217983 173113
rect 218011 173085 218059 173113
rect 217749 173051 218059 173085
rect 217749 173023 217797 173051
rect 217825 173023 217859 173051
rect 217887 173023 217921 173051
rect 217949 173023 217983 173051
rect 218011 173023 218059 173051
rect 217749 172989 218059 173023
rect 217749 172961 217797 172989
rect 217825 172961 217859 172989
rect 217887 172961 217921 172989
rect 217949 172961 217983 172989
rect 218011 172961 218059 172989
rect 204249 167147 204297 167175
rect 204325 167147 204359 167175
rect 204387 167147 204421 167175
rect 204449 167147 204483 167175
rect 204511 167147 204559 167175
rect 204249 167113 204559 167147
rect 204249 167085 204297 167113
rect 204325 167085 204359 167113
rect 204387 167085 204421 167113
rect 204449 167085 204483 167113
rect 204511 167085 204559 167113
rect 204249 167051 204559 167085
rect 204249 167023 204297 167051
rect 204325 167023 204359 167051
rect 204387 167023 204421 167051
rect 204449 167023 204483 167051
rect 204511 167023 204559 167051
rect 204249 166989 204559 167023
rect 204249 166961 204297 166989
rect 204325 166961 204359 166989
rect 204387 166961 204421 166989
rect 204449 166961 204483 166989
rect 204511 166961 204559 166989
rect 204249 158175 204559 166961
rect 215584 167175 215744 167192
rect 215584 167147 215619 167175
rect 215647 167147 215681 167175
rect 215709 167147 215744 167175
rect 215584 167113 215744 167147
rect 215584 167085 215619 167113
rect 215647 167085 215681 167113
rect 215709 167085 215744 167113
rect 215584 167051 215744 167085
rect 215584 167023 215619 167051
rect 215647 167023 215681 167051
rect 215709 167023 215744 167051
rect 215584 166989 215744 167023
rect 215584 166961 215619 166989
rect 215647 166961 215681 166989
rect 215709 166961 215744 166989
rect 215584 166944 215744 166961
rect 207904 164175 208064 164192
rect 207904 164147 207939 164175
rect 207967 164147 208001 164175
rect 208029 164147 208064 164175
rect 207904 164113 208064 164147
rect 207904 164085 207939 164113
rect 207967 164085 208001 164113
rect 208029 164085 208064 164113
rect 207904 164051 208064 164085
rect 207904 164023 207939 164051
rect 207967 164023 208001 164051
rect 208029 164023 208064 164051
rect 207904 163989 208064 164023
rect 207904 163961 207939 163989
rect 207967 163961 208001 163989
rect 208029 163961 208064 163989
rect 207904 163944 208064 163961
rect 217749 164175 218059 172961
rect 217749 164147 217797 164175
rect 217825 164147 217859 164175
rect 217887 164147 217921 164175
rect 217949 164147 217983 164175
rect 218011 164147 218059 164175
rect 217749 164113 218059 164147
rect 217749 164085 217797 164113
rect 217825 164085 217859 164113
rect 217887 164085 217921 164113
rect 217949 164085 217983 164113
rect 218011 164085 218059 164113
rect 217749 164051 218059 164085
rect 217749 164023 217797 164051
rect 217825 164023 217859 164051
rect 217887 164023 217921 164051
rect 217949 164023 217983 164051
rect 218011 164023 218059 164051
rect 217749 163989 218059 164023
rect 217749 163961 217797 163989
rect 217825 163961 217859 163989
rect 217887 163961 217921 163989
rect 217949 163961 217983 163989
rect 218011 163961 218059 163989
rect 204249 158147 204297 158175
rect 204325 158147 204359 158175
rect 204387 158147 204421 158175
rect 204449 158147 204483 158175
rect 204511 158147 204559 158175
rect 204249 158113 204559 158147
rect 204249 158085 204297 158113
rect 204325 158085 204359 158113
rect 204387 158085 204421 158113
rect 204449 158085 204483 158113
rect 204511 158085 204559 158113
rect 204249 158051 204559 158085
rect 204249 158023 204297 158051
rect 204325 158023 204359 158051
rect 204387 158023 204421 158051
rect 204449 158023 204483 158051
rect 204511 158023 204559 158051
rect 204249 157989 204559 158023
rect 204249 157961 204297 157989
rect 204325 157961 204359 157989
rect 204387 157961 204421 157989
rect 204449 157961 204483 157989
rect 204511 157961 204559 157989
rect 204249 149175 204559 157961
rect 215584 158175 215744 158192
rect 215584 158147 215619 158175
rect 215647 158147 215681 158175
rect 215709 158147 215744 158175
rect 215584 158113 215744 158147
rect 215584 158085 215619 158113
rect 215647 158085 215681 158113
rect 215709 158085 215744 158113
rect 215584 158051 215744 158085
rect 215584 158023 215619 158051
rect 215647 158023 215681 158051
rect 215709 158023 215744 158051
rect 215584 157989 215744 158023
rect 215584 157961 215619 157989
rect 215647 157961 215681 157989
rect 215709 157961 215744 157989
rect 215584 157944 215744 157961
rect 207904 155175 208064 155192
rect 207904 155147 207939 155175
rect 207967 155147 208001 155175
rect 208029 155147 208064 155175
rect 207904 155113 208064 155147
rect 207904 155085 207939 155113
rect 207967 155085 208001 155113
rect 208029 155085 208064 155113
rect 207904 155051 208064 155085
rect 207904 155023 207939 155051
rect 207967 155023 208001 155051
rect 208029 155023 208064 155051
rect 207904 154989 208064 155023
rect 207904 154961 207939 154989
rect 207967 154961 208001 154989
rect 208029 154961 208064 154989
rect 207904 154944 208064 154961
rect 217749 155175 218059 163961
rect 217749 155147 217797 155175
rect 217825 155147 217859 155175
rect 217887 155147 217921 155175
rect 217949 155147 217983 155175
rect 218011 155147 218059 155175
rect 217749 155113 218059 155147
rect 217749 155085 217797 155113
rect 217825 155085 217859 155113
rect 217887 155085 217921 155113
rect 217949 155085 217983 155113
rect 218011 155085 218059 155113
rect 217749 155051 218059 155085
rect 217749 155023 217797 155051
rect 217825 155023 217859 155051
rect 217887 155023 217921 155051
rect 217949 155023 217983 155051
rect 218011 155023 218059 155051
rect 217749 154989 218059 155023
rect 217749 154961 217797 154989
rect 217825 154961 217859 154989
rect 217887 154961 217921 154989
rect 217949 154961 217983 154989
rect 218011 154961 218059 154989
rect 204249 149147 204297 149175
rect 204325 149147 204359 149175
rect 204387 149147 204421 149175
rect 204449 149147 204483 149175
rect 204511 149147 204559 149175
rect 204249 149113 204559 149147
rect 204249 149085 204297 149113
rect 204325 149085 204359 149113
rect 204387 149085 204421 149113
rect 204449 149085 204483 149113
rect 204511 149085 204559 149113
rect 204249 149051 204559 149085
rect 204249 149023 204297 149051
rect 204325 149023 204359 149051
rect 204387 149023 204421 149051
rect 204449 149023 204483 149051
rect 204511 149023 204559 149051
rect 204249 148989 204559 149023
rect 204249 148961 204297 148989
rect 204325 148961 204359 148989
rect 204387 148961 204421 148989
rect 204449 148961 204483 148989
rect 204511 148961 204559 148989
rect 204249 140175 204559 148961
rect 215584 149175 215744 149192
rect 215584 149147 215619 149175
rect 215647 149147 215681 149175
rect 215709 149147 215744 149175
rect 215584 149113 215744 149147
rect 215584 149085 215619 149113
rect 215647 149085 215681 149113
rect 215709 149085 215744 149113
rect 215584 149051 215744 149085
rect 215584 149023 215619 149051
rect 215647 149023 215681 149051
rect 215709 149023 215744 149051
rect 215584 148989 215744 149023
rect 215584 148961 215619 148989
rect 215647 148961 215681 148989
rect 215709 148961 215744 148989
rect 215584 148944 215744 148961
rect 207904 146175 208064 146192
rect 207904 146147 207939 146175
rect 207967 146147 208001 146175
rect 208029 146147 208064 146175
rect 207904 146113 208064 146147
rect 207904 146085 207939 146113
rect 207967 146085 208001 146113
rect 208029 146085 208064 146113
rect 207904 146051 208064 146085
rect 207904 146023 207939 146051
rect 207967 146023 208001 146051
rect 208029 146023 208064 146051
rect 207904 145989 208064 146023
rect 207904 145961 207939 145989
rect 207967 145961 208001 145989
rect 208029 145961 208064 145989
rect 207904 145944 208064 145961
rect 217749 146175 218059 154961
rect 217749 146147 217797 146175
rect 217825 146147 217859 146175
rect 217887 146147 217921 146175
rect 217949 146147 217983 146175
rect 218011 146147 218059 146175
rect 217749 146113 218059 146147
rect 217749 146085 217797 146113
rect 217825 146085 217859 146113
rect 217887 146085 217921 146113
rect 217949 146085 217983 146113
rect 218011 146085 218059 146113
rect 217749 146051 218059 146085
rect 217749 146023 217797 146051
rect 217825 146023 217859 146051
rect 217887 146023 217921 146051
rect 217949 146023 217983 146051
rect 218011 146023 218059 146051
rect 217749 145989 218059 146023
rect 217749 145961 217797 145989
rect 217825 145961 217859 145989
rect 217887 145961 217921 145989
rect 217949 145961 217983 145989
rect 218011 145961 218059 145989
rect 204249 140147 204297 140175
rect 204325 140147 204359 140175
rect 204387 140147 204421 140175
rect 204449 140147 204483 140175
rect 204511 140147 204559 140175
rect 204249 140113 204559 140147
rect 204249 140085 204297 140113
rect 204325 140085 204359 140113
rect 204387 140085 204421 140113
rect 204449 140085 204483 140113
rect 204511 140085 204559 140113
rect 204249 140051 204559 140085
rect 204249 140023 204297 140051
rect 204325 140023 204359 140051
rect 204387 140023 204421 140051
rect 204449 140023 204483 140051
rect 204511 140023 204559 140051
rect 204249 139989 204559 140023
rect 204249 139961 204297 139989
rect 204325 139961 204359 139989
rect 204387 139961 204421 139989
rect 204449 139961 204483 139989
rect 204511 139961 204559 139989
rect 204249 131175 204559 139961
rect 215584 140175 215744 140192
rect 215584 140147 215619 140175
rect 215647 140147 215681 140175
rect 215709 140147 215744 140175
rect 215584 140113 215744 140147
rect 215584 140085 215619 140113
rect 215647 140085 215681 140113
rect 215709 140085 215744 140113
rect 215584 140051 215744 140085
rect 215584 140023 215619 140051
rect 215647 140023 215681 140051
rect 215709 140023 215744 140051
rect 215584 139989 215744 140023
rect 215584 139961 215619 139989
rect 215647 139961 215681 139989
rect 215709 139961 215744 139989
rect 215584 139944 215744 139961
rect 207904 137175 208064 137192
rect 207904 137147 207939 137175
rect 207967 137147 208001 137175
rect 208029 137147 208064 137175
rect 207904 137113 208064 137147
rect 207904 137085 207939 137113
rect 207967 137085 208001 137113
rect 208029 137085 208064 137113
rect 207904 137051 208064 137085
rect 207904 137023 207939 137051
rect 207967 137023 208001 137051
rect 208029 137023 208064 137051
rect 207904 136989 208064 137023
rect 207904 136961 207939 136989
rect 207967 136961 208001 136989
rect 208029 136961 208064 136989
rect 207904 136944 208064 136961
rect 217749 137175 218059 145961
rect 217749 137147 217797 137175
rect 217825 137147 217859 137175
rect 217887 137147 217921 137175
rect 217949 137147 217983 137175
rect 218011 137147 218059 137175
rect 217749 137113 218059 137147
rect 217749 137085 217797 137113
rect 217825 137085 217859 137113
rect 217887 137085 217921 137113
rect 217949 137085 217983 137113
rect 218011 137085 218059 137113
rect 217749 137051 218059 137085
rect 217749 137023 217797 137051
rect 217825 137023 217859 137051
rect 217887 137023 217921 137051
rect 217949 137023 217983 137051
rect 218011 137023 218059 137051
rect 217749 136989 218059 137023
rect 217749 136961 217797 136989
rect 217825 136961 217859 136989
rect 217887 136961 217921 136989
rect 217949 136961 217983 136989
rect 218011 136961 218059 136989
rect 204249 131147 204297 131175
rect 204325 131147 204359 131175
rect 204387 131147 204421 131175
rect 204449 131147 204483 131175
rect 204511 131147 204559 131175
rect 204249 131113 204559 131147
rect 204249 131085 204297 131113
rect 204325 131085 204359 131113
rect 204387 131085 204421 131113
rect 204449 131085 204483 131113
rect 204511 131085 204559 131113
rect 204249 131051 204559 131085
rect 204249 131023 204297 131051
rect 204325 131023 204359 131051
rect 204387 131023 204421 131051
rect 204449 131023 204483 131051
rect 204511 131023 204559 131051
rect 204249 130989 204559 131023
rect 204249 130961 204297 130989
rect 204325 130961 204359 130989
rect 204387 130961 204421 130989
rect 204449 130961 204483 130989
rect 204511 130961 204559 130989
rect 204249 122175 204559 130961
rect 215584 131175 215744 131192
rect 215584 131147 215619 131175
rect 215647 131147 215681 131175
rect 215709 131147 215744 131175
rect 215584 131113 215744 131147
rect 215584 131085 215619 131113
rect 215647 131085 215681 131113
rect 215709 131085 215744 131113
rect 215584 131051 215744 131085
rect 215584 131023 215619 131051
rect 215647 131023 215681 131051
rect 215709 131023 215744 131051
rect 215584 130989 215744 131023
rect 215584 130961 215619 130989
rect 215647 130961 215681 130989
rect 215709 130961 215744 130989
rect 215584 130944 215744 130961
rect 207904 128175 208064 128192
rect 207904 128147 207939 128175
rect 207967 128147 208001 128175
rect 208029 128147 208064 128175
rect 207904 128113 208064 128147
rect 207904 128085 207939 128113
rect 207967 128085 208001 128113
rect 208029 128085 208064 128113
rect 207904 128051 208064 128085
rect 207904 128023 207939 128051
rect 207967 128023 208001 128051
rect 208029 128023 208064 128051
rect 207904 127989 208064 128023
rect 207904 127961 207939 127989
rect 207967 127961 208001 127989
rect 208029 127961 208064 127989
rect 207904 127944 208064 127961
rect 217749 128175 218059 136961
rect 217749 128147 217797 128175
rect 217825 128147 217859 128175
rect 217887 128147 217921 128175
rect 217949 128147 217983 128175
rect 218011 128147 218059 128175
rect 217749 128113 218059 128147
rect 217749 128085 217797 128113
rect 217825 128085 217859 128113
rect 217887 128085 217921 128113
rect 217949 128085 217983 128113
rect 218011 128085 218059 128113
rect 217749 128051 218059 128085
rect 217749 128023 217797 128051
rect 217825 128023 217859 128051
rect 217887 128023 217921 128051
rect 217949 128023 217983 128051
rect 218011 128023 218059 128051
rect 217749 127989 218059 128023
rect 217749 127961 217797 127989
rect 217825 127961 217859 127989
rect 217887 127961 217921 127989
rect 217949 127961 217983 127989
rect 218011 127961 218059 127989
rect 204249 122147 204297 122175
rect 204325 122147 204359 122175
rect 204387 122147 204421 122175
rect 204449 122147 204483 122175
rect 204511 122147 204559 122175
rect 204249 122113 204559 122147
rect 204249 122085 204297 122113
rect 204325 122085 204359 122113
rect 204387 122085 204421 122113
rect 204449 122085 204483 122113
rect 204511 122085 204559 122113
rect 204249 122051 204559 122085
rect 204249 122023 204297 122051
rect 204325 122023 204359 122051
rect 204387 122023 204421 122051
rect 204449 122023 204483 122051
rect 204511 122023 204559 122051
rect 204249 121989 204559 122023
rect 204249 121961 204297 121989
rect 204325 121961 204359 121989
rect 204387 121961 204421 121989
rect 204449 121961 204483 121989
rect 204511 121961 204559 121989
rect 204249 113175 204559 121961
rect 215584 122175 215744 122192
rect 215584 122147 215619 122175
rect 215647 122147 215681 122175
rect 215709 122147 215744 122175
rect 215584 122113 215744 122147
rect 215584 122085 215619 122113
rect 215647 122085 215681 122113
rect 215709 122085 215744 122113
rect 215584 122051 215744 122085
rect 215584 122023 215619 122051
rect 215647 122023 215681 122051
rect 215709 122023 215744 122051
rect 215584 121989 215744 122023
rect 215584 121961 215619 121989
rect 215647 121961 215681 121989
rect 215709 121961 215744 121989
rect 215584 121944 215744 121961
rect 207904 119175 208064 119192
rect 207904 119147 207939 119175
rect 207967 119147 208001 119175
rect 208029 119147 208064 119175
rect 207904 119113 208064 119147
rect 207904 119085 207939 119113
rect 207967 119085 208001 119113
rect 208029 119085 208064 119113
rect 207904 119051 208064 119085
rect 207904 119023 207939 119051
rect 207967 119023 208001 119051
rect 208029 119023 208064 119051
rect 207904 118989 208064 119023
rect 207904 118961 207939 118989
rect 207967 118961 208001 118989
rect 208029 118961 208064 118989
rect 207904 118944 208064 118961
rect 217749 119175 218059 127961
rect 217749 119147 217797 119175
rect 217825 119147 217859 119175
rect 217887 119147 217921 119175
rect 217949 119147 217983 119175
rect 218011 119147 218059 119175
rect 217749 119113 218059 119147
rect 217749 119085 217797 119113
rect 217825 119085 217859 119113
rect 217887 119085 217921 119113
rect 217949 119085 217983 119113
rect 218011 119085 218059 119113
rect 217749 119051 218059 119085
rect 217749 119023 217797 119051
rect 217825 119023 217859 119051
rect 217887 119023 217921 119051
rect 217949 119023 217983 119051
rect 218011 119023 218059 119051
rect 217749 118989 218059 119023
rect 217749 118961 217797 118989
rect 217825 118961 217859 118989
rect 217887 118961 217921 118989
rect 217949 118961 217983 118989
rect 218011 118961 218059 118989
rect 204249 113147 204297 113175
rect 204325 113147 204359 113175
rect 204387 113147 204421 113175
rect 204449 113147 204483 113175
rect 204511 113147 204559 113175
rect 204249 113113 204559 113147
rect 204249 113085 204297 113113
rect 204325 113085 204359 113113
rect 204387 113085 204421 113113
rect 204449 113085 204483 113113
rect 204511 113085 204559 113113
rect 204249 113051 204559 113085
rect 204249 113023 204297 113051
rect 204325 113023 204359 113051
rect 204387 113023 204421 113051
rect 204449 113023 204483 113051
rect 204511 113023 204559 113051
rect 204249 112989 204559 113023
rect 204249 112961 204297 112989
rect 204325 112961 204359 112989
rect 204387 112961 204421 112989
rect 204449 112961 204483 112989
rect 204511 112961 204559 112989
rect 204249 104175 204559 112961
rect 215584 113175 215744 113192
rect 215584 113147 215619 113175
rect 215647 113147 215681 113175
rect 215709 113147 215744 113175
rect 215584 113113 215744 113147
rect 215584 113085 215619 113113
rect 215647 113085 215681 113113
rect 215709 113085 215744 113113
rect 215584 113051 215744 113085
rect 215584 113023 215619 113051
rect 215647 113023 215681 113051
rect 215709 113023 215744 113051
rect 215584 112989 215744 113023
rect 215584 112961 215619 112989
rect 215647 112961 215681 112989
rect 215709 112961 215744 112989
rect 215584 112944 215744 112961
rect 207904 110175 208064 110192
rect 207904 110147 207939 110175
rect 207967 110147 208001 110175
rect 208029 110147 208064 110175
rect 207904 110113 208064 110147
rect 207904 110085 207939 110113
rect 207967 110085 208001 110113
rect 208029 110085 208064 110113
rect 207904 110051 208064 110085
rect 207904 110023 207939 110051
rect 207967 110023 208001 110051
rect 208029 110023 208064 110051
rect 207904 109989 208064 110023
rect 207904 109961 207939 109989
rect 207967 109961 208001 109989
rect 208029 109961 208064 109989
rect 207904 109944 208064 109961
rect 217749 110175 218059 118961
rect 217749 110147 217797 110175
rect 217825 110147 217859 110175
rect 217887 110147 217921 110175
rect 217949 110147 217983 110175
rect 218011 110147 218059 110175
rect 217749 110113 218059 110147
rect 217749 110085 217797 110113
rect 217825 110085 217859 110113
rect 217887 110085 217921 110113
rect 217949 110085 217983 110113
rect 218011 110085 218059 110113
rect 217749 110051 218059 110085
rect 217749 110023 217797 110051
rect 217825 110023 217859 110051
rect 217887 110023 217921 110051
rect 217949 110023 217983 110051
rect 218011 110023 218059 110051
rect 217749 109989 218059 110023
rect 217749 109961 217797 109989
rect 217825 109961 217859 109989
rect 217887 109961 217921 109989
rect 217949 109961 217983 109989
rect 218011 109961 218059 109989
rect 204249 104147 204297 104175
rect 204325 104147 204359 104175
rect 204387 104147 204421 104175
rect 204449 104147 204483 104175
rect 204511 104147 204559 104175
rect 204249 104113 204559 104147
rect 204249 104085 204297 104113
rect 204325 104085 204359 104113
rect 204387 104085 204421 104113
rect 204449 104085 204483 104113
rect 204511 104085 204559 104113
rect 204249 104051 204559 104085
rect 204249 104023 204297 104051
rect 204325 104023 204359 104051
rect 204387 104023 204421 104051
rect 204449 104023 204483 104051
rect 204511 104023 204559 104051
rect 204249 103989 204559 104023
rect 204249 103961 204297 103989
rect 204325 103961 204359 103989
rect 204387 103961 204421 103989
rect 204449 103961 204483 103989
rect 204511 103961 204559 103989
rect 204249 95175 204559 103961
rect 215584 104175 215744 104192
rect 215584 104147 215619 104175
rect 215647 104147 215681 104175
rect 215709 104147 215744 104175
rect 215584 104113 215744 104147
rect 215584 104085 215619 104113
rect 215647 104085 215681 104113
rect 215709 104085 215744 104113
rect 215584 104051 215744 104085
rect 215584 104023 215619 104051
rect 215647 104023 215681 104051
rect 215709 104023 215744 104051
rect 215584 103989 215744 104023
rect 215584 103961 215619 103989
rect 215647 103961 215681 103989
rect 215709 103961 215744 103989
rect 215584 103944 215744 103961
rect 207904 101175 208064 101192
rect 207904 101147 207939 101175
rect 207967 101147 208001 101175
rect 208029 101147 208064 101175
rect 207904 101113 208064 101147
rect 207904 101085 207939 101113
rect 207967 101085 208001 101113
rect 208029 101085 208064 101113
rect 207904 101051 208064 101085
rect 207904 101023 207939 101051
rect 207967 101023 208001 101051
rect 208029 101023 208064 101051
rect 207904 100989 208064 101023
rect 207904 100961 207939 100989
rect 207967 100961 208001 100989
rect 208029 100961 208064 100989
rect 207904 100944 208064 100961
rect 217749 101175 218059 109961
rect 217749 101147 217797 101175
rect 217825 101147 217859 101175
rect 217887 101147 217921 101175
rect 217949 101147 217983 101175
rect 218011 101147 218059 101175
rect 217749 101113 218059 101147
rect 217749 101085 217797 101113
rect 217825 101085 217859 101113
rect 217887 101085 217921 101113
rect 217949 101085 217983 101113
rect 218011 101085 218059 101113
rect 217749 101051 218059 101085
rect 217749 101023 217797 101051
rect 217825 101023 217859 101051
rect 217887 101023 217921 101051
rect 217949 101023 217983 101051
rect 218011 101023 218059 101051
rect 217749 100989 218059 101023
rect 217749 100961 217797 100989
rect 217825 100961 217859 100989
rect 217887 100961 217921 100989
rect 217949 100961 217983 100989
rect 218011 100961 218059 100989
rect 204249 95147 204297 95175
rect 204325 95147 204359 95175
rect 204387 95147 204421 95175
rect 204449 95147 204483 95175
rect 204511 95147 204559 95175
rect 204249 95113 204559 95147
rect 204249 95085 204297 95113
rect 204325 95085 204359 95113
rect 204387 95085 204421 95113
rect 204449 95085 204483 95113
rect 204511 95085 204559 95113
rect 204249 95051 204559 95085
rect 204249 95023 204297 95051
rect 204325 95023 204359 95051
rect 204387 95023 204421 95051
rect 204449 95023 204483 95051
rect 204511 95023 204559 95051
rect 204249 94989 204559 95023
rect 204249 94961 204297 94989
rect 204325 94961 204359 94989
rect 204387 94961 204421 94989
rect 204449 94961 204483 94989
rect 204511 94961 204559 94989
rect 204249 86175 204559 94961
rect 215584 95175 215744 95192
rect 215584 95147 215619 95175
rect 215647 95147 215681 95175
rect 215709 95147 215744 95175
rect 215584 95113 215744 95147
rect 215584 95085 215619 95113
rect 215647 95085 215681 95113
rect 215709 95085 215744 95113
rect 215584 95051 215744 95085
rect 215584 95023 215619 95051
rect 215647 95023 215681 95051
rect 215709 95023 215744 95051
rect 215584 94989 215744 95023
rect 215584 94961 215619 94989
rect 215647 94961 215681 94989
rect 215709 94961 215744 94989
rect 215584 94944 215744 94961
rect 207904 92175 208064 92192
rect 207904 92147 207939 92175
rect 207967 92147 208001 92175
rect 208029 92147 208064 92175
rect 207904 92113 208064 92147
rect 207904 92085 207939 92113
rect 207967 92085 208001 92113
rect 208029 92085 208064 92113
rect 207904 92051 208064 92085
rect 207904 92023 207939 92051
rect 207967 92023 208001 92051
rect 208029 92023 208064 92051
rect 207904 91989 208064 92023
rect 207904 91961 207939 91989
rect 207967 91961 208001 91989
rect 208029 91961 208064 91989
rect 207904 91944 208064 91961
rect 217749 92175 218059 100961
rect 217749 92147 217797 92175
rect 217825 92147 217859 92175
rect 217887 92147 217921 92175
rect 217949 92147 217983 92175
rect 218011 92147 218059 92175
rect 217749 92113 218059 92147
rect 217749 92085 217797 92113
rect 217825 92085 217859 92113
rect 217887 92085 217921 92113
rect 217949 92085 217983 92113
rect 218011 92085 218059 92113
rect 217749 92051 218059 92085
rect 217749 92023 217797 92051
rect 217825 92023 217859 92051
rect 217887 92023 217921 92051
rect 217949 92023 217983 92051
rect 218011 92023 218059 92051
rect 217749 91989 218059 92023
rect 217749 91961 217797 91989
rect 217825 91961 217859 91989
rect 217887 91961 217921 91989
rect 217949 91961 217983 91989
rect 218011 91961 218059 91989
rect 204249 86147 204297 86175
rect 204325 86147 204359 86175
rect 204387 86147 204421 86175
rect 204449 86147 204483 86175
rect 204511 86147 204559 86175
rect 204249 86113 204559 86147
rect 204249 86085 204297 86113
rect 204325 86085 204359 86113
rect 204387 86085 204421 86113
rect 204449 86085 204483 86113
rect 204511 86085 204559 86113
rect 204249 86051 204559 86085
rect 204249 86023 204297 86051
rect 204325 86023 204359 86051
rect 204387 86023 204421 86051
rect 204449 86023 204483 86051
rect 204511 86023 204559 86051
rect 204249 85989 204559 86023
rect 204249 85961 204297 85989
rect 204325 85961 204359 85989
rect 204387 85961 204421 85989
rect 204449 85961 204483 85989
rect 204511 85961 204559 85989
rect 204249 77175 204559 85961
rect 215584 86175 215744 86192
rect 215584 86147 215619 86175
rect 215647 86147 215681 86175
rect 215709 86147 215744 86175
rect 215584 86113 215744 86147
rect 215584 86085 215619 86113
rect 215647 86085 215681 86113
rect 215709 86085 215744 86113
rect 215584 86051 215744 86085
rect 215584 86023 215619 86051
rect 215647 86023 215681 86051
rect 215709 86023 215744 86051
rect 215584 85989 215744 86023
rect 215584 85961 215619 85989
rect 215647 85961 215681 85989
rect 215709 85961 215744 85989
rect 215584 85944 215744 85961
rect 207904 83175 208064 83192
rect 207904 83147 207939 83175
rect 207967 83147 208001 83175
rect 208029 83147 208064 83175
rect 207904 83113 208064 83147
rect 207904 83085 207939 83113
rect 207967 83085 208001 83113
rect 208029 83085 208064 83113
rect 207904 83051 208064 83085
rect 207904 83023 207939 83051
rect 207967 83023 208001 83051
rect 208029 83023 208064 83051
rect 207904 82989 208064 83023
rect 207904 82961 207939 82989
rect 207967 82961 208001 82989
rect 208029 82961 208064 82989
rect 207904 82944 208064 82961
rect 217749 83175 218059 91961
rect 217749 83147 217797 83175
rect 217825 83147 217859 83175
rect 217887 83147 217921 83175
rect 217949 83147 217983 83175
rect 218011 83147 218059 83175
rect 217749 83113 218059 83147
rect 217749 83085 217797 83113
rect 217825 83085 217859 83113
rect 217887 83085 217921 83113
rect 217949 83085 217983 83113
rect 218011 83085 218059 83113
rect 217749 83051 218059 83085
rect 217749 83023 217797 83051
rect 217825 83023 217859 83051
rect 217887 83023 217921 83051
rect 217949 83023 217983 83051
rect 218011 83023 218059 83051
rect 217749 82989 218059 83023
rect 217749 82961 217797 82989
rect 217825 82961 217859 82989
rect 217887 82961 217921 82989
rect 217949 82961 217983 82989
rect 218011 82961 218059 82989
rect 204249 77147 204297 77175
rect 204325 77147 204359 77175
rect 204387 77147 204421 77175
rect 204449 77147 204483 77175
rect 204511 77147 204559 77175
rect 204249 77113 204559 77147
rect 204249 77085 204297 77113
rect 204325 77085 204359 77113
rect 204387 77085 204421 77113
rect 204449 77085 204483 77113
rect 204511 77085 204559 77113
rect 204249 77051 204559 77085
rect 204249 77023 204297 77051
rect 204325 77023 204359 77051
rect 204387 77023 204421 77051
rect 204449 77023 204483 77051
rect 204511 77023 204559 77051
rect 204249 76989 204559 77023
rect 204249 76961 204297 76989
rect 204325 76961 204359 76989
rect 204387 76961 204421 76989
rect 204449 76961 204483 76989
rect 204511 76961 204559 76989
rect 204249 68175 204559 76961
rect 215584 77175 215744 77192
rect 215584 77147 215619 77175
rect 215647 77147 215681 77175
rect 215709 77147 215744 77175
rect 215584 77113 215744 77147
rect 215584 77085 215619 77113
rect 215647 77085 215681 77113
rect 215709 77085 215744 77113
rect 215584 77051 215744 77085
rect 215584 77023 215619 77051
rect 215647 77023 215681 77051
rect 215709 77023 215744 77051
rect 215584 76989 215744 77023
rect 215584 76961 215619 76989
rect 215647 76961 215681 76989
rect 215709 76961 215744 76989
rect 215584 76944 215744 76961
rect 207904 74175 208064 74192
rect 207904 74147 207939 74175
rect 207967 74147 208001 74175
rect 208029 74147 208064 74175
rect 207904 74113 208064 74147
rect 207904 74085 207939 74113
rect 207967 74085 208001 74113
rect 208029 74085 208064 74113
rect 207904 74051 208064 74085
rect 207904 74023 207939 74051
rect 207967 74023 208001 74051
rect 208029 74023 208064 74051
rect 207904 73989 208064 74023
rect 207904 73961 207939 73989
rect 207967 73961 208001 73989
rect 208029 73961 208064 73989
rect 207904 73944 208064 73961
rect 217749 74175 218059 82961
rect 217749 74147 217797 74175
rect 217825 74147 217859 74175
rect 217887 74147 217921 74175
rect 217949 74147 217983 74175
rect 218011 74147 218059 74175
rect 217749 74113 218059 74147
rect 217749 74085 217797 74113
rect 217825 74085 217859 74113
rect 217887 74085 217921 74113
rect 217949 74085 217983 74113
rect 218011 74085 218059 74113
rect 217749 74051 218059 74085
rect 217749 74023 217797 74051
rect 217825 74023 217859 74051
rect 217887 74023 217921 74051
rect 217949 74023 217983 74051
rect 218011 74023 218059 74051
rect 217749 73989 218059 74023
rect 217749 73961 217797 73989
rect 217825 73961 217859 73989
rect 217887 73961 217921 73989
rect 217949 73961 217983 73989
rect 218011 73961 218059 73989
rect 204249 68147 204297 68175
rect 204325 68147 204359 68175
rect 204387 68147 204421 68175
rect 204449 68147 204483 68175
rect 204511 68147 204559 68175
rect 204249 68113 204559 68147
rect 204249 68085 204297 68113
rect 204325 68085 204359 68113
rect 204387 68085 204421 68113
rect 204449 68085 204483 68113
rect 204511 68085 204559 68113
rect 204249 68051 204559 68085
rect 204249 68023 204297 68051
rect 204325 68023 204359 68051
rect 204387 68023 204421 68051
rect 204449 68023 204483 68051
rect 204511 68023 204559 68051
rect 204249 67989 204559 68023
rect 204249 67961 204297 67989
rect 204325 67961 204359 67989
rect 204387 67961 204421 67989
rect 204449 67961 204483 67989
rect 204511 67961 204559 67989
rect 204249 59175 204559 67961
rect 215584 68175 215744 68192
rect 215584 68147 215619 68175
rect 215647 68147 215681 68175
rect 215709 68147 215744 68175
rect 215584 68113 215744 68147
rect 215584 68085 215619 68113
rect 215647 68085 215681 68113
rect 215709 68085 215744 68113
rect 215584 68051 215744 68085
rect 215584 68023 215619 68051
rect 215647 68023 215681 68051
rect 215709 68023 215744 68051
rect 215584 67989 215744 68023
rect 215584 67961 215619 67989
rect 215647 67961 215681 67989
rect 215709 67961 215744 67989
rect 215584 67944 215744 67961
rect 207904 65175 208064 65192
rect 207904 65147 207939 65175
rect 207967 65147 208001 65175
rect 208029 65147 208064 65175
rect 207904 65113 208064 65147
rect 207904 65085 207939 65113
rect 207967 65085 208001 65113
rect 208029 65085 208064 65113
rect 207904 65051 208064 65085
rect 207904 65023 207939 65051
rect 207967 65023 208001 65051
rect 208029 65023 208064 65051
rect 207904 64989 208064 65023
rect 207904 64961 207939 64989
rect 207967 64961 208001 64989
rect 208029 64961 208064 64989
rect 207904 64944 208064 64961
rect 217749 65175 218059 73961
rect 217749 65147 217797 65175
rect 217825 65147 217859 65175
rect 217887 65147 217921 65175
rect 217949 65147 217983 65175
rect 218011 65147 218059 65175
rect 217749 65113 218059 65147
rect 217749 65085 217797 65113
rect 217825 65085 217859 65113
rect 217887 65085 217921 65113
rect 217949 65085 217983 65113
rect 218011 65085 218059 65113
rect 217749 65051 218059 65085
rect 217749 65023 217797 65051
rect 217825 65023 217859 65051
rect 217887 65023 217921 65051
rect 217949 65023 217983 65051
rect 218011 65023 218059 65051
rect 217749 64989 218059 65023
rect 217749 64961 217797 64989
rect 217825 64961 217859 64989
rect 217887 64961 217921 64989
rect 217949 64961 217983 64989
rect 218011 64961 218059 64989
rect 204249 59147 204297 59175
rect 204325 59147 204359 59175
rect 204387 59147 204421 59175
rect 204449 59147 204483 59175
rect 204511 59147 204559 59175
rect 204249 59113 204559 59147
rect 204249 59085 204297 59113
rect 204325 59085 204359 59113
rect 204387 59085 204421 59113
rect 204449 59085 204483 59113
rect 204511 59085 204559 59113
rect 204249 59051 204559 59085
rect 204249 59023 204297 59051
rect 204325 59023 204359 59051
rect 204387 59023 204421 59051
rect 204449 59023 204483 59051
rect 204511 59023 204559 59051
rect 204249 58989 204559 59023
rect 204249 58961 204297 58989
rect 204325 58961 204359 58989
rect 204387 58961 204421 58989
rect 204449 58961 204483 58989
rect 204511 58961 204559 58989
rect 204249 50175 204559 58961
rect 215584 59175 215744 59192
rect 215584 59147 215619 59175
rect 215647 59147 215681 59175
rect 215709 59147 215744 59175
rect 215584 59113 215744 59147
rect 215584 59085 215619 59113
rect 215647 59085 215681 59113
rect 215709 59085 215744 59113
rect 215584 59051 215744 59085
rect 215584 59023 215619 59051
rect 215647 59023 215681 59051
rect 215709 59023 215744 59051
rect 215584 58989 215744 59023
rect 215584 58961 215619 58989
rect 215647 58961 215681 58989
rect 215709 58961 215744 58989
rect 215584 58944 215744 58961
rect 207904 56175 208064 56192
rect 207904 56147 207939 56175
rect 207967 56147 208001 56175
rect 208029 56147 208064 56175
rect 207904 56113 208064 56147
rect 207904 56085 207939 56113
rect 207967 56085 208001 56113
rect 208029 56085 208064 56113
rect 207904 56051 208064 56085
rect 207904 56023 207939 56051
rect 207967 56023 208001 56051
rect 208029 56023 208064 56051
rect 207904 55989 208064 56023
rect 207904 55961 207939 55989
rect 207967 55961 208001 55989
rect 208029 55961 208064 55989
rect 207904 55944 208064 55961
rect 217749 56175 218059 64961
rect 217749 56147 217797 56175
rect 217825 56147 217859 56175
rect 217887 56147 217921 56175
rect 217949 56147 217983 56175
rect 218011 56147 218059 56175
rect 217749 56113 218059 56147
rect 217749 56085 217797 56113
rect 217825 56085 217859 56113
rect 217887 56085 217921 56113
rect 217949 56085 217983 56113
rect 218011 56085 218059 56113
rect 217749 56051 218059 56085
rect 217749 56023 217797 56051
rect 217825 56023 217859 56051
rect 217887 56023 217921 56051
rect 217949 56023 217983 56051
rect 218011 56023 218059 56051
rect 217749 55989 218059 56023
rect 217749 55961 217797 55989
rect 217825 55961 217859 55989
rect 217887 55961 217921 55989
rect 217949 55961 217983 55989
rect 218011 55961 218059 55989
rect 204249 50147 204297 50175
rect 204325 50147 204359 50175
rect 204387 50147 204421 50175
rect 204449 50147 204483 50175
rect 204511 50147 204559 50175
rect 204249 50113 204559 50147
rect 204249 50085 204297 50113
rect 204325 50085 204359 50113
rect 204387 50085 204421 50113
rect 204449 50085 204483 50113
rect 204511 50085 204559 50113
rect 204249 50051 204559 50085
rect 204249 50023 204297 50051
rect 204325 50023 204359 50051
rect 204387 50023 204421 50051
rect 204449 50023 204483 50051
rect 204511 50023 204559 50051
rect 204249 49989 204559 50023
rect 204249 49961 204297 49989
rect 204325 49961 204359 49989
rect 204387 49961 204421 49989
rect 204449 49961 204483 49989
rect 204511 49961 204559 49989
rect 204249 41175 204559 49961
rect 215584 50175 215744 50192
rect 215584 50147 215619 50175
rect 215647 50147 215681 50175
rect 215709 50147 215744 50175
rect 215584 50113 215744 50147
rect 215584 50085 215619 50113
rect 215647 50085 215681 50113
rect 215709 50085 215744 50113
rect 215584 50051 215744 50085
rect 215584 50023 215619 50051
rect 215647 50023 215681 50051
rect 215709 50023 215744 50051
rect 215584 49989 215744 50023
rect 215584 49961 215619 49989
rect 215647 49961 215681 49989
rect 215709 49961 215744 49989
rect 215584 49944 215744 49961
rect 207904 47175 208064 47192
rect 207904 47147 207939 47175
rect 207967 47147 208001 47175
rect 208029 47147 208064 47175
rect 207904 47113 208064 47147
rect 207904 47085 207939 47113
rect 207967 47085 208001 47113
rect 208029 47085 208064 47113
rect 207904 47051 208064 47085
rect 207904 47023 207939 47051
rect 207967 47023 208001 47051
rect 208029 47023 208064 47051
rect 207904 46989 208064 47023
rect 207904 46961 207939 46989
rect 207967 46961 208001 46989
rect 208029 46961 208064 46989
rect 207904 46944 208064 46961
rect 217749 47175 218059 55961
rect 217749 47147 217797 47175
rect 217825 47147 217859 47175
rect 217887 47147 217921 47175
rect 217949 47147 217983 47175
rect 218011 47147 218059 47175
rect 217749 47113 218059 47147
rect 217749 47085 217797 47113
rect 217825 47085 217859 47113
rect 217887 47085 217921 47113
rect 217949 47085 217983 47113
rect 218011 47085 218059 47113
rect 217749 47051 218059 47085
rect 217749 47023 217797 47051
rect 217825 47023 217859 47051
rect 217887 47023 217921 47051
rect 217949 47023 217983 47051
rect 218011 47023 218059 47051
rect 217749 46989 218059 47023
rect 217749 46961 217797 46989
rect 217825 46961 217859 46989
rect 217887 46961 217921 46989
rect 217949 46961 217983 46989
rect 218011 46961 218059 46989
rect 204249 41147 204297 41175
rect 204325 41147 204359 41175
rect 204387 41147 204421 41175
rect 204449 41147 204483 41175
rect 204511 41147 204559 41175
rect 204249 41113 204559 41147
rect 204249 41085 204297 41113
rect 204325 41085 204359 41113
rect 204387 41085 204421 41113
rect 204449 41085 204483 41113
rect 204511 41085 204559 41113
rect 204249 41051 204559 41085
rect 204249 41023 204297 41051
rect 204325 41023 204359 41051
rect 204387 41023 204421 41051
rect 204449 41023 204483 41051
rect 204511 41023 204559 41051
rect 204249 40989 204559 41023
rect 204249 40961 204297 40989
rect 204325 40961 204359 40989
rect 204387 40961 204421 40989
rect 204449 40961 204483 40989
rect 204511 40961 204559 40989
rect 204249 32175 204559 40961
rect 215584 41175 215744 41192
rect 215584 41147 215619 41175
rect 215647 41147 215681 41175
rect 215709 41147 215744 41175
rect 215584 41113 215744 41147
rect 215584 41085 215619 41113
rect 215647 41085 215681 41113
rect 215709 41085 215744 41113
rect 215584 41051 215744 41085
rect 215584 41023 215619 41051
rect 215647 41023 215681 41051
rect 215709 41023 215744 41051
rect 215584 40989 215744 41023
rect 215584 40961 215619 40989
rect 215647 40961 215681 40989
rect 215709 40961 215744 40989
rect 215584 40944 215744 40961
rect 207904 38175 208064 38192
rect 207904 38147 207939 38175
rect 207967 38147 208001 38175
rect 208029 38147 208064 38175
rect 207904 38113 208064 38147
rect 207904 38085 207939 38113
rect 207967 38085 208001 38113
rect 208029 38085 208064 38113
rect 207904 38051 208064 38085
rect 207904 38023 207939 38051
rect 207967 38023 208001 38051
rect 208029 38023 208064 38051
rect 207904 37989 208064 38023
rect 207904 37961 207939 37989
rect 207967 37961 208001 37989
rect 208029 37961 208064 37989
rect 207904 37944 208064 37961
rect 217749 38175 218059 46961
rect 217749 38147 217797 38175
rect 217825 38147 217859 38175
rect 217887 38147 217921 38175
rect 217949 38147 217983 38175
rect 218011 38147 218059 38175
rect 217749 38113 218059 38147
rect 217749 38085 217797 38113
rect 217825 38085 217859 38113
rect 217887 38085 217921 38113
rect 217949 38085 217983 38113
rect 218011 38085 218059 38113
rect 217749 38051 218059 38085
rect 217749 38023 217797 38051
rect 217825 38023 217859 38051
rect 217887 38023 217921 38051
rect 217949 38023 217983 38051
rect 218011 38023 218059 38051
rect 217749 37989 218059 38023
rect 217749 37961 217797 37989
rect 217825 37961 217859 37989
rect 217887 37961 217921 37989
rect 217949 37961 217983 37989
rect 218011 37961 218059 37989
rect 204249 32147 204297 32175
rect 204325 32147 204359 32175
rect 204387 32147 204421 32175
rect 204449 32147 204483 32175
rect 204511 32147 204559 32175
rect 204249 32113 204559 32147
rect 204249 32085 204297 32113
rect 204325 32085 204359 32113
rect 204387 32085 204421 32113
rect 204449 32085 204483 32113
rect 204511 32085 204559 32113
rect 204249 32051 204559 32085
rect 204249 32023 204297 32051
rect 204325 32023 204359 32051
rect 204387 32023 204421 32051
rect 204449 32023 204483 32051
rect 204511 32023 204559 32051
rect 204249 31989 204559 32023
rect 204249 31961 204297 31989
rect 204325 31961 204359 31989
rect 204387 31961 204421 31989
rect 204449 31961 204483 31989
rect 204511 31961 204559 31989
rect 204249 23175 204559 31961
rect 215584 32175 215744 32192
rect 215584 32147 215619 32175
rect 215647 32147 215681 32175
rect 215709 32147 215744 32175
rect 215584 32113 215744 32147
rect 215584 32085 215619 32113
rect 215647 32085 215681 32113
rect 215709 32085 215744 32113
rect 215584 32051 215744 32085
rect 215584 32023 215619 32051
rect 215647 32023 215681 32051
rect 215709 32023 215744 32051
rect 215584 31989 215744 32023
rect 215584 31961 215619 31989
rect 215647 31961 215681 31989
rect 215709 31961 215744 31989
rect 215584 31944 215744 31961
rect 207904 29175 208064 29192
rect 207904 29147 207939 29175
rect 207967 29147 208001 29175
rect 208029 29147 208064 29175
rect 207904 29113 208064 29147
rect 207904 29085 207939 29113
rect 207967 29085 208001 29113
rect 208029 29085 208064 29113
rect 207904 29051 208064 29085
rect 207904 29023 207939 29051
rect 207967 29023 208001 29051
rect 208029 29023 208064 29051
rect 207904 28989 208064 29023
rect 207904 28961 207939 28989
rect 207967 28961 208001 28989
rect 208029 28961 208064 28989
rect 207904 28944 208064 28961
rect 217749 29175 218059 37961
rect 217749 29147 217797 29175
rect 217825 29147 217859 29175
rect 217887 29147 217921 29175
rect 217949 29147 217983 29175
rect 218011 29147 218059 29175
rect 217749 29113 218059 29147
rect 217749 29085 217797 29113
rect 217825 29085 217859 29113
rect 217887 29085 217921 29113
rect 217949 29085 217983 29113
rect 218011 29085 218059 29113
rect 217749 29051 218059 29085
rect 217749 29023 217797 29051
rect 217825 29023 217859 29051
rect 217887 29023 217921 29051
rect 217949 29023 217983 29051
rect 218011 29023 218059 29051
rect 217749 28989 218059 29023
rect 217749 28961 217797 28989
rect 217825 28961 217859 28989
rect 217887 28961 217921 28989
rect 217949 28961 217983 28989
rect 218011 28961 218059 28989
rect 204249 23147 204297 23175
rect 204325 23147 204359 23175
rect 204387 23147 204421 23175
rect 204449 23147 204483 23175
rect 204511 23147 204559 23175
rect 204249 23113 204559 23147
rect 204249 23085 204297 23113
rect 204325 23085 204359 23113
rect 204387 23085 204421 23113
rect 204449 23085 204483 23113
rect 204511 23085 204559 23113
rect 204249 23051 204559 23085
rect 204249 23023 204297 23051
rect 204325 23023 204359 23051
rect 204387 23023 204421 23051
rect 204449 23023 204483 23051
rect 204511 23023 204559 23051
rect 204249 22989 204559 23023
rect 204249 22961 204297 22989
rect 204325 22961 204359 22989
rect 204387 22961 204421 22989
rect 204449 22961 204483 22989
rect 204511 22961 204559 22989
rect 204249 14175 204559 22961
rect 215584 23175 215744 23192
rect 215584 23147 215619 23175
rect 215647 23147 215681 23175
rect 215709 23147 215744 23175
rect 215584 23113 215744 23147
rect 215584 23085 215619 23113
rect 215647 23085 215681 23113
rect 215709 23085 215744 23113
rect 215584 23051 215744 23085
rect 215584 23023 215619 23051
rect 215647 23023 215681 23051
rect 215709 23023 215744 23051
rect 215584 22989 215744 23023
rect 215584 22961 215619 22989
rect 215647 22961 215681 22989
rect 215709 22961 215744 22989
rect 215584 22944 215744 22961
rect 207904 20175 208064 20192
rect 207904 20147 207939 20175
rect 207967 20147 208001 20175
rect 208029 20147 208064 20175
rect 207904 20113 208064 20147
rect 207904 20085 207939 20113
rect 207967 20085 208001 20113
rect 208029 20085 208064 20113
rect 207904 20051 208064 20085
rect 207904 20023 207939 20051
rect 207967 20023 208001 20051
rect 208029 20023 208064 20051
rect 207904 19989 208064 20023
rect 207904 19961 207939 19989
rect 207967 19961 208001 19989
rect 208029 19961 208064 19989
rect 207904 19944 208064 19961
rect 217749 20175 218059 28961
rect 217749 20147 217797 20175
rect 217825 20147 217859 20175
rect 217887 20147 217921 20175
rect 217949 20147 217983 20175
rect 218011 20147 218059 20175
rect 217749 20113 218059 20147
rect 217749 20085 217797 20113
rect 217825 20085 217859 20113
rect 217887 20085 217921 20113
rect 217949 20085 217983 20113
rect 218011 20085 218059 20113
rect 217749 20051 218059 20085
rect 217749 20023 217797 20051
rect 217825 20023 217859 20051
rect 217887 20023 217921 20051
rect 217949 20023 217983 20051
rect 218011 20023 218059 20051
rect 217749 19989 218059 20023
rect 217749 19961 217797 19989
rect 217825 19961 217859 19989
rect 217887 19961 217921 19989
rect 217949 19961 217983 19989
rect 218011 19961 218059 19989
rect 204249 14147 204297 14175
rect 204325 14147 204359 14175
rect 204387 14147 204421 14175
rect 204449 14147 204483 14175
rect 204511 14147 204559 14175
rect 204249 14113 204559 14147
rect 204249 14085 204297 14113
rect 204325 14085 204359 14113
rect 204387 14085 204421 14113
rect 204449 14085 204483 14113
rect 204511 14085 204559 14113
rect 204249 14051 204559 14085
rect 204249 14023 204297 14051
rect 204325 14023 204359 14051
rect 204387 14023 204421 14051
rect 204449 14023 204483 14051
rect 204511 14023 204559 14051
rect 204249 13989 204559 14023
rect 204249 13961 204297 13989
rect 204325 13961 204359 13989
rect 204387 13961 204421 13989
rect 204449 13961 204483 13989
rect 204511 13961 204559 13989
rect 204249 5175 204559 13961
rect 215584 14175 215744 14192
rect 215584 14147 215619 14175
rect 215647 14147 215681 14175
rect 215709 14147 215744 14175
rect 215584 14113 215744 14147
rect 215584 14085 215619 14113
rect 215647 14085 215681 14113
rect 215709 14085 215744 14113
rect 215584 14051 215744 14085
rect 215584 14023 215619 14051
rect 215647 14023 215681 14051
rect 215709 14023 215744 14051
rect 215584 13989 215744 14023
rect 215584 13961 215619 13989
rect 215647 13961 215681 13989
rect 215709 13961 215744 13989
rect 215584 13944 215744 13961
rect 207904 11175 208064 11192
rect 207904 11147 207939 11175
rect 207967 11147 208001 11175
rect 208029 11147 208064 11175
rect 207904 11113 208064 11147
rect 207904 11085 207939 11113
rect 207967 11085 208001 11113
rect 208029 11085 208064 11113
rect 207904 11051 208064 11085
rect 207904 11023 207939 11051
rect 207967 11023 208001 11051
rect 208029 11023 208064 11051
rect 207904 10989 208064 11023
rect 207904 10961 207939 10989
rect 207967 10961 208001 10989
rect 208029 10961 208064 10989
rect 207904 10944 208064 10961
rect 217749 11175 218059 19961
rect 217749 11147 217797 11175
rect 217825 11147 217859 11175
rect 217887 11147 217921 11175
rect 217949 11147 217983 11175
rect 218011 11147 218059 11175
rect 217749 11113 218059 11147
rect 217749 11085 217797 11113
rect 217825 11085 217859 11113
rect 217887 11085 217921 11113
rect 217949 11085 217983 11113
rect 218011 11085 218059 11113
rect 217749 11051 218059 11085
rect 217749 11023 217797 11051
rect 217825 11023 217859 11051
rect 217887 11023 217921 11051
rect 217949 11023 217983 11051
rect 218011 11023 218059 11051
rect 217749 10989 218059 11023
rect 217749 10961 217797 10989
rect 217825 10961 217859 10989
rect 217887 10961 217921 10989
rect 217949 10961 217983 10989
rect 218011 10961 218059 10989
rect 204249 5147 204297 5175
rect 204325 5147 204359 5175
rect 204387 5147 204421 5175
rect 204449 5147 204483 5175
rect 204511 5147 204559 5175
rect 204249 5113 204559 5147
rect 204249 5085 204297 5113
rect 204325 5085 204359 5113
rect 204387 5085 204421 5113
rect 204449 5085 204483 5113
rect 204511 5085 204559 5113
rect 204249 5051 204559 5085
rect 204249 5023 204297 5051
rect 204325 5023 204359 5051
rect 204387 5023 204421 5051
rect 204449 5023 204483 5051
rect 204511 5023 204559 5051
rect 204249 4989 204559 5023
rect 204249 4961 204297 4989
rect 204325 4961 204359 4989
rect 204387 4961 204421 4989
rect 204449 4961 204483 4989
rect 204511 4961 204559 4989
rect 204249 -560 204559 4961
rect 215584 5175 215744 5192
rect 215584 5147 215619 5175
rect 215647 5147 215681 5175
rect 215709 5147 215744 5175
rect 215584 5113 215744 5147
rect 215584 5085 215619 5113
rect 215647 5085 215681 5113
rect 215709 5085 215744 5113
rect 215584 5051 215744 5085
rect 215584 5023 215619 5051
rect 215647 5023 215681 5051
rect 215709 5023 215744 5051
rect 215584 4989 215744 5023
rect 215584 4961 215619 4989
rect 215647 4961 215681 4989
rect 215709 4961 215744 4989
rect 215584 4944 215744 4961
rect 204249 -588 204297 -560
rect 204325 -588 204359 -560
rect 204387 -588 204421 -560
rect 204449 -588 204483 -560
rect 204511 -588 204559 -560
rect 204249 -622 204559 -588
rect 204249 -650 204297 -622
rect 204325 -650 204359 -622
rect 204387 -650 204421 -622
rect 204449 -650 204483 -622
rect 204511 -650 204559 -622
rect 204249 -684 204559 -650
rect 204249 -712 204297 -684
rect 204325 -712 204359 -684
rect 204387 -712 204421 -684
rect 204449 -712 204483 -684
rect 204511 -712 204559 -684
rect 204249 -746 204559 -712
rect 204249 -774 204297 -746
rect 204325 -774 204359 -746
rect 204387 -774 204421 -746
rect 204449 -774 204483 -746
rect 204511 -774 204559 -746
rect 204249 -822 204559 -774
rect 217749 2175 218059 10961
rect 217749 2147 217797 2175
rect 217825 2147 217859 2175
rect 217887 2147 217921 2175
rect 217949 2147 217983 2175
rect 218011 2147 218059 2175
rect 217749 2113 218059 2147
rect 217749 2085 217797 2113
rect 217825 2085 217859 2113
rect 217887 2085 217921 2113
rect 217949 2085 217983 2113
rect 218011 2085 218059 2113
rect 217749 2051 218059 2085
rect 217749 2023 217797 2051
rect 217825 2023 217859 2051
rect 217887 2023 217921 2051
rect 217949 2023 217983 2051
rect 218011 2023 218059 2051
rect 217749 1989 218059 2023
rect 217749 1961 217797 1989
rect 217825 1961 217859 1989
rect 217887 1961 217921 1989
rect 217949 1961 217983 1989
rect 218011 1961 218059 1989
rect 217749 -80 218059 1961
rect 217749 -108 217797 -80
rect 217825 -108 217859 -80
rect 217887 -108 217921 -80
rect 217949 -108 217983 -80
rect 218011 -108 218059 -80
rect 217749 -142 218059 -108
rect 217749 -170 217797 -142
rect 217825 -170 217859 -142
rect 217887 -170 217921 -142
rect 217949 -170 217983 -142
rect 218011 -170 218059 -142
rect 217749 -204 218059 -170
rect 217749 -232 217797 -204
rect 217825 -232 217859 -204
rect 217887 -232 217921 -204
rect 217949 -232 217983 -204
rect 218011 -232 218059 -204
rect 217749 -266 218059 -232
rect 217749 -294 217797 -266
rect 217825 -294 217859 -266
rect 217887 -294 217921 -266
rect 217949 -294 217983 -266
rect 218011 -294 218059 -266
rect 217749 -822 218059 -294
rect 219609 299086 219919 299134
rect 219609 299058 219657 299086
rect 219685 299058 219719 299086
rect 219747 299058 219781 299086
rect 219809 299058 219843 299086
rect 219871 299058 219919 299086
rect 219609 299024 219919 299058
rect 219609 298996 219657 299024
rect 219685 298996 219719 299024
rect 219747 298996 219781 299024
rect 219809 298996 219843 299024
rect 219871 298996 219919 299024
rect 219609 298962 219919 298996
rect 219609 298934 219657 298962
rect 219685 298934 219719 298962
rect 219747 298934 219781 298962
rect 219809 298934 219843 298962
rect 219871 298934 219919 298962
rect 219609 298900 219919 298934
rect 219609 298872 219657 298900
rect 219685 298872 219719 298900
rect 219747 298872 219781 298900
rect 219809 298872 219843 298900
rect 219871 298872 219919 298900
rect 219609 293175 219919 298872
rect 219609 293147 219657 293175
rect 219685 293147 219719 293175
rect 219747 293147 219781 293175
rect 219809 293147 219843 293175
rect 219871 293147 219919 293175
rect 219609 293113 219919 293147
rect 219609 293085 219657 293113
rect 219685 293085 219719 293113
rect 219747 293085 219781 293113
rect 219809 293085 219843 293113
rect 219871 293085 219919 293113
rect 219609 293051 219919 293085
rect 219609 293023 219657 293051
rect 219685 293023 219719 293051
rect 219747 293023 219781 293051
rect 219809 293023 219843 293051
rect 219871 293023 219919 293051
rect 219609 292989 219919 293023
rect 219609 292961 219657 292989
rect 219685 292961 219719 292989
rect 219747 292961 219781 292989
rect 219809 292961 219843 292989
rect 219871 292961 219919 292989
rect 219609 284175 219919 292961
rect 219609 284147 219657 284175
rect 219685 284147 219719 284175
rect 219747 284147 219781 284175
rect 219809 284147 219843 284175
rect 219871 284147 219919 284175
rect 219609 284113 219919 284147
rect 219609 284085 219657 284113
rect 219685 284085 219719 284113
rect 219747 284085 219781 284113
rect 219809 284085 219843 284113
rect 219871 284085 219919 284113
rect 219609 284051 219919 284085
rect 219609 284023 219657 284051
rect 219685 284023 219719 284051
rect 219747 284023 219781 284051
rect 219809 284023 219843 284051
rect 219871 284023 219919 284051
rect 219609 283989 219919 284023
rect 219609 283961 219657 283989
rect 219685 283961 219719 283989
rect 219747 283961 219781 283989
rect 219809 283961 219843 283989
rect 219871 283961 219919 283989
rect 219609 275175 219919 283961
rect 219609 275147 219657 275175
rect 219685 275147 219719 275175
rect 219747 275147 219781 275175
rect 219809 275147 219843 275175
rect 219871 275147 219919 275175
rect 219609 275113 219919 275147
rect 219609 275085 219657 275113
rect 219685 275085 219719 275113
rect 219747 275085 219781 275113
rect 219809 275085 219843 275113
rect 219871 275085 219919 275113
rect 219609 275051 219919 275085
rect 219609 275023 219657 275051
rect 219685 275023 219719 275051
rect 219747 275023 219781 275051
rect 219809 275023 219843 275051
rect 219871 275023 219919 275051
rect 219609 274989 219919 275023
rect 219609 274961 219657 274989
rect 219685 274961 219719 274989
rect 219747 274961 219781 274989
rect 219809 274961 219843 274989
rect 219871 274961 219919 274989
rect 219609 266175 219919 274961
rect 219609 266147 219657 266175
rect 219685 266147 219719 266175
rect 219747 266147 219781 266175
rect 219809 266147 219843 266175
rect 219871 266147 219919 266175
rect 219609 266113 219919 266147
rect 219609 266085 219657 266113
rect 219685 266085 219719 266113
rect 219747 266085 219781 266113
rect 219809 266085 219843 266113
rect 219871 266085 219919 266113
rect 219609 266051 219919 266085
rect 219609 266023 219657 266051
rect 219685 266023 219719 266051
rect 219747 266023 219781 266051
rect 219809 266023 219843 266051
rect 219871 266023 219919 266051
rect 219609 265989 219919 266023
rect 219609 265961 219657 265989
rect 219685 265961 219719 265989
rect 219747 265961 219781 265989
rect 219809 265961 219843 265989
rect 219871 265961 219919 265989
rect 219609 257175 219919 265961
rect 219609 257147 219657 257175
rect 219685 257147 219719 257175
rect 219747 257147 219781 257175
rect 219809 257147 219843 257175
rect 219871 257147 219919 257175
rect 219609 257113 219919 257147
rect 219609 257085 219657 257113
rect 219685 257085 219719 257113
rect 219747 257085 219781 257113
rect 219809 257085 219843 257113
rect 219871 257085 219919 257113
rect 219609 257051 219919 257085
rect 219609 257023 219657 257051
rect 219685 257023 219719 257051
rect 219747 257023 219781 257051
rect 219809 257023 219843 257051
rect 219871 257023 219919 257051
rect 219609 256989 219919 257023
rect 219609 256961 219657 256989
rect 219685 256961 219719 256989
rect 219747 256961 219781 256989
rect 219809 256961 219843 256989
rect 219871 256961 219919 256989
rect 219609 248175 219919 256961
rect 219609 248147 219657 248175
rect 219685 248147 219719 248175
rect 219747 248147 219781 248175
rect 219809 248147 219843 248175
rect 219871 248147 219919 248175
rect 219609 248113 219919 248147
rect 219609 248085 219657 248113
rect 219685 248085 219719 248113
rect 219747 248085 219781 248113
rect 219809 248085 219843 248113
rect 219871 248085 219919 248113
rect 219609 248051 219919 248085
rect 219609 248023 219657 248051
rect 219685 248023 219719 248051
rect 219747 248023 219781 248051
rect 219809 248023 219843 248051
rect 219871 248023 219919 248051
rect 219609 247989 219919 248023
rect 219609 247961 219657 247989
rect 219685 247961 219719 247989
rect 219747 247961 219781 247989
rect 219809 247961 219843 247989
rect 219871 247961 219919 247989
rect 219609 239175 219919 247961
rect 219609 239147 219657 239175
rect 219685 239147 219719 239175
rect 219747 239147 219781 239175
rect 219809 239147 219843 239175
rect 219871 239147 219919 239175
rect 219609 239113 219919 239147
rect 219609 239085 219657 239113
rect 219685 239085 219719 239113
rect 219747 239085 219781 239113
rect 219809 239085 219843 239113
rect 219871 239085 219919 239113
rect 219609 239051 219919 239085
rect 219609 239023 219657 239051
rect 219685 239023 219719 239051
rect 219747 239023 219781 239051
rect 219809 239023 219843 239051
rect 219871 239023 219919 239051
rect 219609 238989 219919 239023
rect 219609 238961 219657 238989
rect 219685 238961 219719 238989
rect 219747 238961 219781 238989
rect 219809 238961 219843 238989
rect 219871 238961 219919 238989
rect 219609 230175 219919 238961
rect 219609 230147 219657 230175
rect 219685 230147 219719 230175
rect 219747 230147 219781 230175
rect 219809 230147 219843 230175
rect 219871 230147 219919 230175
rect 219609 230113 219919 230147
rect 219609 230085 219657 230113
rect 219685 230085 219719 230113
rect 219747 230085 219781 230113
rect 219809 230085 219843 230113
rect 219871 230085 219919 230113
rect 219609 230051 219919 230085
rect 219609 230023 219657 230051
rect 219685 230023 219719 230051
rect 219747 230023 219781 230051
rect 219809 230023 219843 230051
rect 219871 230023 219919 230051
rect 219609 229989 219919 230023
rect 219609 229961 219657 229989
rect 219685 229961 219719 229989
rect 219747 229961 219781 229989
rect 219809 229961 219843 229989
rect 219871 229961 219919 229989
rect 219609 221175 219919 229961
rect 219609 221147 219657 221175
rect 219685 221147 219719 221175
rect 219747 221147 219781 221175
rect 219809 221147 219843 221175
rect 219871 221147 219919 221175
rect 219609 221113 219919 221147
rect 219609 221085 219657 221113
rect 219685 221085 219719 221113
rect 219747 221085 219781 221113
rect 219809 221085 219843 221113
rect 219871 221085 219919 221113
rect 219609 221051 219919 221085
rect 219609 221023 219657 221051
rect 219685 221023 219719 221051
rect 219747 221023 219781 221051
rect 219809 221023 219843 221051
rect 219871 221023 219919 221051
rect 219609 220989 219919 221023
rect 219609 220961 219657 220989
rect 219685 220961 219719 220989
rect 219747 220961 219781 220989
rect 219809 220961 219843 220989
rect 219871 220961 219919 220989
rect 219609 212175 219919 220961
rect 219609 212147 219657 212175
rect 219685 212147 219719 212175
rect 219747 212147 219781 212175
rect 219809 212147 219843 212175
rect 219871 212147 219919 212175
rect 219609 212113 219919 212147
rect 219609 212085 219657 212113
rect 219685 212085 219719 212113
rect 219747 212085 219781 212113
rect 219809 212085 219843 212113
rect 219871 212085 219919 212113
rect 219609 212051 219919 212085
rect 219609 212023 219657 212051
rect 219685 212023 219719 212051
rect 219747 212023 219781 212051
rect 219809 212023 219843 212051
rect 219871 212023 219919 212051
rect 219609 211989 219919 212023
rect 219609 211961 219657 211989
rect 219685 211961 219719 211989
rect 219747 211961 219781 211989
rect 219809 211961 219843 211989
rect 219871 211961 219919 211989
rect 219609 203175 219919 211961
rect 219609 203147 219657 203175
rect 219685 203147 219719 203175
rect 219747 203147 219781 203175
rect 219809 203147 219843 203175
rect 219871 203147 219919 203175
rect 219609 203113 219919 203147
rect 219609 203085 219657 203113
rect 219685 203085 219719 203113
rect 219747 203085 219781 203113
rect 219809 203085 219843 203113
rect 219871 203085 219919 203113
rect 219609 203051 219919 203085
rect 219609 203023 219657 203051
rect 219685 203023 219719 203051
rect 219747 203023 219781 203051
rect 219809 203023 219843 203051
rect 219871 203023 219919 203051
rect 219609 202989 219919 203023
rect 219609 202961 219657 202989
rect 219685 202961 219719 202989
rect 219747 202961 219781 202989
rect 219809 202961 219843 202989
rect 219871 202961 219919 202989
rect 219609 194175 219919 202961
rect 219609 194147 219657 194175
rect 219685 194147 219719 194175
rect 219747 194147 219781 194175
rect 219809 194147 219843 194175
rect 219871 194147 219919 194175
rect 219609 194113 219919 194147
rect 219609 194085 219657 194113
rect 219685 194085 219719 194113
rect 219747 194085 219781 194113
rect 219809 194085 219843 194113
rect 219871 194085 219919 194113
rect 219609 194051 219919 194085
rect 219609 194023 219657 194051
rect 219685 194023 219719 194051
rect 219747 194023 219781 194051
rect 219809 194023 219843 194051
rect 219871 194023 219919 194051
rect 219609 193989 219919 194023
rect 219609 193961 219657 193989
rect 219685 193961 219719 193989
rect 219747 193961 219781 193989
rect 219809 193961 219843 193989
rect 219871 193961 219919 193989
rect 219609 185175 219919 193961
rect 219609 185147 219657 185175
rect 219685 185147 219719 185175
rect 219747 185147 219781 185175
rect 219809 185147 219843 185175
rect 219871 185147 219919 185175
rect 219609 185113 219919 185147
rect 219609 185085 219657 185113
rect 219685 185085 219719 185113
rect 219747 185085 219781 185113
rect 219809 185085 219843 185113
rect 219871 185085 219919 185113
rect 219609 185051 219919 185085
rect 219609 185023 219657 185051
rect 219685 185023 219719 185051
rect 219747 185023 219781 185051
rect 219809 185023 219843 185051
rect 219871 185023 219919 185051
rect 219609 184989 219919 185023
rect 219609 184961 219657 184989
rect 219685 184961 219719 184989
rect 219747 184961 219781 184989
rect 219809 184961 219843 184989
rect 219871 184961 219919 184989
rect 219609 176175 219919 184961
rect 219609 176147 219657 176175
rect 219685 176147 219719 176175
rect 219747 176147 219781 176175
rect 219809 176147 219843 176175
rect 219871 176147 219919 176175
rect 219609 176113 219919 176147
rect 219609 176085 219657 176113
rect 219685 176085 219719 176113
rect 219747 176085 219781 176113
rect 219809 176085 219843 176113
rect 219871 176085 219919 176113
rect 219609 176051 219919 176085
rect 219609 176023 219657 176051
rect 219685 176023 219719 176051
rect 219747 176023 219781 176051
rect 219809 176023 219843 176051
rect 219871 176023 219919 176051
rect 219609 175989 219919 176023
rect 219609 175961 219657 175989
rect 219685 175961 219719 175989
rect 219747 175961 219781 175989
rect 219809 175961 219843 175989
rect 219871 175961 219919 175989
rect 219609 167175 219919 175961
rect 233109 298606 233419 299134
rect 233109 298578 233157 298606
rect 233185 298578 233219 298606
rect 233247 298578 233281 298606
rect 233309 298578 233343 298606
rect 233371 298578 233419 298606
rect 233109 298544 233419 298578
rect 233109 298516 233157 298544
rect 233185 298516 233219 298544
rect 233247 298516 233281 298544
rect 233309 298516 233343 298544
rect 233371 298516 233419 298544
rect 233109 298482 233419 298516
rect 233109 298454 233157 298482
rect 233185 298454 233219 298482
rect 233247 298454 233281 298482
rect 233309 298454 233343 298482
rect 233371 298454 233419 298482
rect 233109 298420 233419 298454
rect 233109 298392 233157 298420
rect 233185 298392 233219 298420
rect 233247 298392 233281 298420
rect 233309 298392 233343 298420
rect 233371 298392 233419 298420
rect 233109 290175 233419 298392
rect 233109 290147 233157 290175
rect 233185 290147 233219 290175
rect 233247 290147 233281 290175
rect 233309 290147 233343 290175
rect 233371 290147 233419 290175
rect 233109 290113 233419 290147
rect 233109 290085 233157 290113
rect 233185 290085 233219 290113
rect 233247 290085 233281 290113
rect 233309 290085 233343 290113
rect 233371 290085 233419 290113
rect 233109 290051 233419 290085
rect 233109 290023 233157 290051
rect 233185 290023 233219 290051
rect 233247 290023 233281 290051
rect 233309 290023 233343 290051
rect 233371 290023 233419 290051
rect 233109 289989 233419 290023
rect 233109 289961 233157 289989
rect 233185 289961 233219 289989
rect 233247 289961 233281 289989
rect 233309 289961 233343 289989
rect 233371 289961 233419 289989
rect 233109 281175 233419 289961
rect 233109 281147 233157 281175
rect 233185 281147 233219 281175
rect 233247 281147 233281 281175
rect 233309 281147 233343 281175
rect 233371 281147 233419 281175
rect 233109 281113 233419 281147
rect 233109 281085 233157 281113
rect 233185 281085 233219 281113
rect 233247 281085 233281 281113
rect 233309 281085 233343 281113
rect 233371 281085 233419 281113
rect 233109 281051 233419 281085
rect 233109 281023 233157 281051
rect 233185 281023 233219 281051
rect 233247 281023 233281 281051
rect 233309 281023 233343 281051
rect 233371 281023 233419 281051
rect 233109 280989 233419 281023
rect 233109 280961 233157 280989
rect 233185 280961 233219 280989
rect 233247 280961 233281 280989
rect 233309 280961 233343 280989
rect 233371 280961 233419 280989
rect 233109 272175 233419 280961
rect 233109 272147 233157 272175
rect 233185 272147 233219 272175
rect 233247 272147 233281 272175
rect 233309 272147 233343 272175
rect 233371 272147 233419 272175
rect 233109 272113 233419 272147
rect 233109 272085 233157 272113
rect 233185 272085 233219 272113
rect 233247 272085 233281 272113
rect 233309 272085 233343 272113
rect 233371 272085 233419 272113
rect 233109 272051 233419 272085
rect 233109 272023 233157 272051
rect 233185 272023 233219 272051
rect 233247 272023 233281 272051
rect 233309 272023 233343 272051
rect 233371 272023 233419 272051
rect 233109 271989 233419 272023
rect 233109 271961 233157 271989
rect 233185 271961 233219 271989
rect 233247 271961 233281 271989
rect 233309 271961 233343 271989
rect 233371 271961 233419 271989
rect 233109 263175 233419 271961
rect 233109 263147 233157 263175
rect 233185 263147 233219 263175
rect 233247 263147 233281 263175
rect 233309 263147 233343 263175
rect 233371 263147 233419 263175
rect 233109 263113 233419 263147
rect 233109 263085 233157 263113
rect 233185 263085 233219 263113
rect 233247 263085 233281 263113
rect 233309 263085 233343 263113
rect 233371 263085 233419 263113
rect 233109 263051 233419 263085
rect 233109 263023 233157 263051
rect 233185 263023 233219 263051
rect 233247 263023 233281 263051
rect 233309 263023 233343 263051
rect 233371 263023 233419 263051
rect 233109 262989 233419 263023
rect 233109 262961 233157 262989
rect 233185 262961 233219 262989
rect 233247 262961 233281 262989
rect 233309 262961 233343 262989
rect 233371 262961 233419 262989
rect 233109 254175 233419 262961
rect 233109 254147 233157 254175
rect 233185 254147 233219 254175
rect 233247 254147 233281 254175
rect 233309 254147 233343 254175
rect 233371 254147 233419 254175
rect 233109 254113 233419 254147
rect 233109 254085 233157 254113
rect 233185 254085 233219 254113
rect 233247 254085 233281 254113
rect 233309 254085 233343 254113
rect 233371 254085 233419 254113
rect 233109 254051 233419 254085
rect 233109 254023 233157 254051
rect 233185 254023 233219 254051
rect 233247 254023 233281 254051
rect 233309 254023 233343 254051
rect 233371 254023 233419 254051
rect 233109 253989 233419 254023
rect 233109 253961 233157 253989
rect 233185 253961 233219 253989
rect 233247 253961 233281 253989
rect 233309 253961 233343 253989
rect 233371 253961 233419 253989
rect 233109 245175 233419 253961
rect 233109 245147 233157 245175
rect 233185 245147 233219 245175
rect 233247 245147 233281 245175
rect 233309 245147 233343 245175
rect 233371 245147 233419 245175
rect 233109 245113 233419 245147
rect 233109 245085 233157 245113
rect 233185 245085 233219 245113
rect 233247 245085 233281 245113
rect 233309 245085 233343 245113
rect 233371 245085 233419 245113
rect 233109 245051 233419 245085
rect 233109 245023 233157 245051
rect 233185 245023 233219 245051
rect 233247 245023 233281 245051
rect 233309 245023 233343 245051
rect 233371 245023 233419 245051
rect 233109 244989 233419 245023
rect 233109 244961 233157 244989
rect 233185 244961 233219 244989
rect 233247 244961 233281 244989
rect 233309 244961 233343 244989
rect 233371 244961 233419 244989
rect 233109 236175 233419 244961
rect 233109 236147 233157 236175
rect 233185 236147 233219 236175
rect 233247 236147 233281 236175
rect 233309 236147 233343 236175
rect 233371 236147 233419 236175
rect 233109 236113 233419 236147
rect 233109 236085 233157 236113
rect 233185 236085 233219 236113
rect 233247 236085 233281 236113
rect 233309 236085 233343 236113
rect 233371 236085 233419 236113
rect 233109 236051 233419 236085
rect 233109 236023 233157 236051
rect 233185 236023 233219 236051
rect 233247 236023 233281 236051
rect 233309 236023 233343 236051
rect 233371 236023 233419 236051
rect 233109 235989 233419 236023
rect 233109 235961 233157 235989
rect 233185 235961 233219 235989
rect 233247 235961 233281 235989
rect 233309 235961 233343 235989
rect 233371 235961 233419 235989
rect 233109 227175 233419 235961
rect 233109 227147 233157 227175
rect 233185 227147 233219 227175
rect 233247 227147 233281 227175
rect 233309 227147 233343 227175
rect 233371 227147 233419 227175
rect 233109 227113 233419 227147
rect 233109 227085 233157 227113
rect 233185 227085 233219 227113
rect 233247 227085 233281 227113
rect 233309 227085 233343 227113
rect 233371 227085 233419 227113
rect 233109 227051 233419 227085
rect 233109 227023 233157 227051
rect 233185 227023 233219 227051
rect 233247 227023 233281 227051
rect 233309 227023 233343 227051
rect 233371 227023 233419 227051
rect 233109 226989 233419 227023
rect 233109 226961 233157 226989
rect 233185 226961 233219 226989
rect 233247 226961 233281 226989
rect 233309 226961 233343 226989
rect 233371 226961 233419 226989
rect 233109 218175 233419 226961
rect 233109 218147 233157 218175
rect 233185 218147 233219 218175
rect 233247 218147 233281 218175
rect 233309 218147 233343 218175
rect 233371 218147 233419 218175
rect 233109 218113 233419 218147
rect 233109 218085 233157 218113
rect 233185 218085 233219 218113
rect 233247 218085 233281 218113
rect 233309 218085 233343 218113
rect 233371 218085 233419 218113
rect 233109 218051 233419 218085
rect 233109 218023 233157 218051
rect 233185 218023 233219 218051
rect 233247 218023 233281 218051
rect 233309 218023 233343 218051
rect 233371 218023 233419 218051
rect 233109 217989 233419 218023
rect 233109 217961 233157 217989
rect 233185 217961 233219 217989
rect 233247 217961 233281 217989
rect 233309 217961 233343 217989
rect 233371 217961 233419 217989
rect 233109 209175 233419 217961
rect 233109 209147 233157 209175
rect 233185 209147 233219 209175
rect 233247 209147 233281 209175
rect 233309 209147 233343 209175
rect 233371 209147 233419 209175
rect 233109 209113 233419 209147
rect 233109 209085 233157 209113
rect 233185 209085 233219 209113
rect 233247 209085 233281 209113
rect 233309 209085 233343 209113
rect 233371 209085 233419 209113
rect 233109 209051 233419 209085
rect 233109 209023 233157 209051
rect 233185 209023 233219 209051
rect 233247 209023 233281 209051
rect 233309 209023 233343 209051
rect 233371 209023 233419 209051
rect 233109 208989 233419 209023
rect 233109 208961 233157 208989
rect 233185 208961 233219 208989
rect 233247 208961 233281 208989
rect 233309 208961 233343 208989
rect 233371 208961 233419 208989
rect 233109 200175 233419 208961
rect 233109 200147 233157 200175
rect 233185 200147 233219 200175
rect 233247 200147 233281 200175
rect 233309 200147 233343 200175
rect 233371 200147 233419 200175
rect 233109 200113 233419 200147
rect 233109 200085 233157 200113
rect 233185 200085 233219 200113
rect 233247 200085 233281 200113
rect 233309 200085 233343 200113
rect 233371 200085 233419 200113
rect 233109 200051 233419 200085
rect 233109 200023 233157 200051
rect 233185 200023 233219 200051
rect 233247 200023 233281 200051
rect 233309 200023 233343 200051
rect 233371 200023 233419 200051
rect 233109 199989 233419 200023
rect 233109 199961 233157 199989
rect 233185 199961 233219 199989
rect 233247 199961 233281 199989
rect 233309 199961 233343 199989
rect 233371 199961 233419 199989
rect 233109 191175 233419 199961
rect 233109 191147 233157 191175
rect 233185 191147 233219 191175
rect 233247 191147 233281 191175
rect 233309 191147 233343 191175
rect 233371 191147 233419 191175
rect 233109 191113 233419 191147
rect 233109 191085 233157 191113
rect 233185 191085 233219 191113
rect 233247 191085 233281 191113
rect 233309 191085 233343 191113
rect 233371 191085 233419 191113
rect 233109 191051 233419 191085
rect 233109 191023 233157 191051
rect 233185 191023 233219 191051
rect 233247 191023 233281 191051
rect 233309 191023 233343 191051
rect 233371 191023 233419 191051
rect 233109 190989 233419 191023
rect 233109 190961 233157 190989
rect 233185 190961 233219 190989
rect 233247 190961 233281 190989
rect 233309 190961 233343 190989
rect 233371 190961 233419 190989
rect 233109 182175 233419 190961
rect 233109 182147 233157 182175
rect 233185 182147 233219 182175
rect 233247 182147 233281 182175
rect 233309 182147 233343 182175
rect 233371 182147 233419 182175
rect 233109 182113 233419 182147
rect 233109 182085 233157 182113
rect 233185 182085 233219 182113
rect 233247 182085 233281 182113
rect 233309 182085 233343 182113
rect 233371 182085 233419 182113
rect 233109 182051 233419 182085
rect 233109 182023 233157 182051
rect 233185 182023 233219 182051
rect 233247 182023 233281 182051
rect 233309 182023 233343 182051
rect 233371 182023 233419 182051
rect 233109 181989 233419 182023
rect 233109 181961 233157 181989
rect 233185 181961 233219 181989
rect 233247 181961 233281 181989
rect 233309 181961 233343 181989
rect 233371 181961 233419 181989
rect 223264 173175 223424 173192
rect 223264 173147 223299 173175
rect 223327 173147 223361 173175
rect 223389 173147 223424 173175
rect 223264 173113 223424 173147
rect 223264 173085 223299 173113
rect 223327 173085 223361 173113
rect 223389 173085 223424 173113
rect 223264 173051 223424 173085
rect 223264 173023 223299 173051
rect 223327 173023 223361 173051
rect 223389 173023 223424 173051
rect 223264 172989 223424 173023
rect 223264 172961 223299 172989
rect 223327 172961 223361 172989
rect 223389 172961 223424 172989
rect 223264 172944 223424 172961
rect 233109 173175 233419 181961
rect 233109 173147 233157 173175
rect 233185 173147 233219 173175
rect 233247 173147 233281 173175
rect 233309 173147 233343 173175
rect 233371 173147 233419 173175
rect 233109 173113 233419 173147
rect 233109 173085 233157 173113
rect 233185 173085 233219 173113
rect 233247 173085 233281 173113
rect 233309 173085 233343 173113
rect 233371 173085 233419 173113
rect 233109 173051 233419 173085
rect 233109 173023 233157 173051
rect 233185 173023 233219 173051
rect 233247 173023 233281 173051
rect 233309 173023 233343 173051
rect 233371 173023 233419 173051
rect 233109 172989 233419 173023
rect 233109 172961 233157 172989
rect 233185 172961 233219 172989
rect 233247 172961 233281 172989
rect 233309 172961 233343 172989
rect 233371 172961 233419 172989
rect 219609 167147 219657 167175
rect 219685 167147 219719 167175
rect 219747 167147 219781 167175
rect 219809 167147 219843 167175
rect 219871 167147 219919 167175
rect 219609 167113 219919 167147
rect 219609 167085 219657 167113
rect 219685 167085 219719 167113
rect 219747 167085 219781 167113
rect 219809 167085 219843 167113
rect 219871 167085 219919 167113
rect 219609 167051 219919 167085
rect 219609 167023 219657 167051
rect 219685 167023 219719 167051
rect 219747 167023 219781 167051
rect 219809 167023 219843 167051
rect 219871 167023 219919 167051
rect 219609 166989 219919 167023
rect 219609 166961 219657 166989
rect 219685 166961 219719 166989
rect 219747 166961 219781 166989
rect 219809 166961 219843 166989
rect 219871 166961 219919 166989
rect 219609 158175 219919 166961
rect 230944 167175 231104 167192
rect 230944 167147 230979 167175
rect 231007 167147 231041 167175
rect 231069 167147 231104 167175
rect 230944 167113 231104 167147
rect 230944 167085 230979 167113
rect 231007 167085 231041 167113
rect 231069 167085 231104 167113
rect 230944 167051 231104 167085
rect 230944 167023 230979 167051
rect 231007 167023 231041 167051
rect 231069 167023 231104 167051
rect 230944 166989 231104 167023
rect 230944 166961 230979 166989
rect 231007 166961 231041 166989
rect 231069 166961 231104 166989
rect 230944 166944 231104 166961
rect 223264 164175 223424 164192
rect 223264 164147 223299 164175
rect 223327 164147 223361 164175
rect 223389 164147 223424 164175
rect 223264 164113 223424 164147
rect 223264 164085 223299 164113
rect 223327 164085 223361 164113
rect 223389 164085 223424 164113
rect 223264 164051 223424 164085
rect 223264 164023 223299 164051
rect 223327 164023 223361 164051
rect 223389 164023 223424 164051
rect 223264 163989 223424 164023
rect 223264 163961 223299 163989
rect 223327 163961 223361 163989
rect 223389 163961 223424 163989
rect 223264 163944 223424 163961
rect 233109 164175 233419 172961
rect 233109 164147 233157 164175
rect 233185 164147 233219 164175
rect 233247 164147 233281 164175
rect 233309 164147 233343 164175
rect 233371 164147 233419 164175
rect 233109 164113 233419 164147
rect 233109 164085 233157 164113
rect 233185 164085 233219 164113
rect 233247 164085 233281 164113
rect 233309 164085 233343 164113
rect 233371 164085 233419 164113
rect 233109 164051 233419 164085
rect 233109 164023 233157 164051
rect 233185 164023 233219 164051
rect 233247 164023 233281 164051
rect 233309 164023 233343 164051
rect 233371 164023 233419 164051
rect 233109 163989 233419 164023
rect 233109 163961 233157 163989
rect 233185 163961 233219 163989
rect 233247 163961 233281 163989
rect 233309 163961 233343 163989
rect 233371 163961 233419 163989
rect 219609 158147 219657 158175
rect 219685 158147 219719 158175
rect 219747 158147 219781 158175
rect 219809 158147 219843 158175
rect 219871 158147 219919 158175
rect 219609 158113 219919 158147
rect 219609 158085 219657 158113
rect 219685 158085 219719 158113
rect 219747 158085 219781 158113
rect 219809 158085 219843 158113
rect 219871 158085 219919 158113
rect 219609 158051 219919 158085
rect 219609 158023 219657 158051
rect 219685 158023 219719 158051
rect 219747 158023 219781 158051
rect 219809 158023 219843 158051
rect 219871 158023 219919 158051
rect 219609 157989 219919 158023
rect 219609 157961 219657 157989
rect 219685 157961 219719 157989
rect 219747 157961 219781 157989
rect 219809 157961 219843 157989
rect 219871 157961 219919 157989
rect 219609 149175 219919 157961
rect 230944 158175 231104 158192
rect 230944 158147 230979 158175
rect 231007 158147 231041 158175
rect 231069 158147 231104 158175
rect 230944 158113 231104 158147
rect 230944 158085 230979 158113
rect 231007 158085 231041 158113
rect 231069 158085 231104 158113
rect 230944 158051 231104 158085
rect 230944 158023 230979 158051
rect 231007 158023 231041 158051
rect 231069 158023 231104 158051
rect 230944 157989 231104 158023
rect 230944 157961 230979 157989
rect 231007 157961 231041 157989
rect 231069 157961 231104 157989
rect 230944 157944 231104 157961
rect 223264 155175 223424 155192
rect 223264 155147 223299 155175
rect 223327 155147 223361 155175
rect 223389 155147 223424 155175
rect 223264 155113 223424 155147
rect 223264 155085 223299 155113
rect 223327 155085 223361 155113
rect 223389 155085 223424 155113
rect 223264 155051 223424 155085
rect 223264 155023 223299 155051
rect 223327 155023 223361 155051
rect 223389 155023 223424 155051
rect 223264 154989 223424 155023
rect 223264 154961 223299 154989
rect 223327 154961 223361 154989
rect 223389 154961 223424 154989
rect 223264 154944 223424 154961
rect 233109 155175 233419 163961
rect 233109 155147 233157 155175
rect 233185 155147 233219 155175
rect 233247 155147 233281 155175
rect 233309 155147 233343 155175
rect 233371 155147 233419 155175
rect 233109 155113 233419 155147
rect 233109 155085 233157 155113
rect 233185 155085 233219 155113
rect 233247 155085 233281 155113
rect 233309 155085 233343 155113
rect 233371 155085 233419 155113
rect 233109 155051 233419 155085
rect 233109 155023 233157 155051
rect 233185 155023 233219 155051
rect 233247 155023 233281 155051
rect 233309 155023 233343 155051
rect 233371 155023 233419 155051
rect 233109 154989 233419 155023
rect 233109 154961 233157 154989
rect 233185 154961 233219 154989
rect 233247 154961 233281 154989
rect 233309 154961 233343 154989
rect 233371 154961 233419 154989
rect 219609 149147 219657 149175
rect 219685 149147 219719 149175
rect 219747 149147 219781 149175
rect 219809 149147 219843 149175
rect 219871 149147 219919 149175
rect 219609 149113 219919 149147
rect 219609 149085 219657 149113
rect 219685 149085 219719 149113
rect 219747 149085 219781 149113
rect 219809 149085 219843 149113
rect 219871 149085 219919 149113
rect 219609 149051 219919 149085
rect 219609 149023 219657 149051
rect 219685 149023 219719 149051
rect 219747 149023 219781 149051
rect 219809 149023 219843 149051
rect 219871 149023 219919 149051
rect 219609 148989 219919 149023
rect 219609 148961 219657 148989
rect 219685 148961 219719 148989
rect 219747 148961 219781 148989
rect 219809 148961 219843 148989
rect 219871 148961 219919 148989
rect 219609 140175 219919 148961
rect 230944 149175 231104 149192
rect 230944 149147 230979 149175
rect 231007 149147 231041 149175
rect 231069 149147 231104 149175
rect 230944 149113 231104 149147
rect 230944 149085 230979 149113
rect 231007 149085 231041 149113
rect 231069 149085 231104 149113
rect 230944 149051 231104 149085
rect 230944 149023 230979 149051
rect 231007 149023 231041 149051
rect 231069 149023 231104 149051
rect 230944 148989 231104 149023
rect 230944 148961 230979 148989
rect 231007 148961 231041 148989
rect 231069 148961 231104 148989
rect 230944 148944 231104 148961
rect 223264 146175 223424 146192
rect 223264 146147 223299 146175
rect 223327 146147 223361 146175
rect 223389 146147 223424 146175
rect 223264 146113 223424 146147
rect 223264 146085 223299 146113
rect 223327 146085 223361 146113
rect 223389 146085 223424 146113
rect 223264 146051 223424 146085
rect 223264 146023 223299 146051
rect 223327 146023 223361 146051
rect 223389 146023 223424 146051
rect 223264 145989 223424 146023
rect 223264 145961 223299 145989
rect 223327 145961 223361 145989
rect 223389 145961 223424 145989
rect 223264 145944 223424 145961
rect 233109 146175 233419 154961
rect 233109 146147 233157 146175
rect 233185 146147 233219 146175
rect 233247 146147 233281 146175
rect 233309 146147 233343 146175
rect 233371 146147 233419 146175
rect 233109 146113 233419 146147
rect 233109 146085 233157 146113
rect 233185 146085 233219 146113
rect 233247 146085 233281 146113
rect 233309 146085 233343 146113
rect 233371 146085 233419 146113
rect 233109 146051 233419 146085
rect 233109 146023 233157 146051
rect 233185 146023 233219 146051
rect 233247 146023 233281 146051
rect 233309 146023 233343 146051
rect 233371 146023 233419 146051
rect 233109 145989 233419 146023
rect 233109 145961 233157 145989
rect 233185 145961 233219 145989
rect 233247 145961 233281 145989
rect 233309 145961 233343 145989
rect 233371 145961 233419 145989
rect 219609 140147 219657 140175
rect 219685 140147 219719 140175
rect 219747 140147 219781 140175
rect 219809 140147 219843 140175
rect 219871 140147 219919 140175
rect 219609 140113 219919 140147
rect 219609 140085 219657 140113
rect 219685 140085 219719 140113
rect 219747 140085 219781 140113
rect 219809 140085 219843 140113
rect 219871 140085 219919 140113
rect 219609 140051 219919 140085
rect 219609 140023 219657 140051
rect 219685 140023 219719 140051
rect 219747 140023 219781 140051
rect 219809 140023 219843 140051
rect 219871 140023 219919 140051
rect 219609 139989 219919 140023
rect 219609 139961 219657 139989
rect 219685 139961 219719 139989
rect 219747 139961 219781 139989
rect 219809 139961 219843 139989
rect 219871 139961 219919 139989
rect 219609 131175 219919 139961
rect 230944 140175 231104 140192
rect 230944 140147 230979 140175
rect 231007 140147 231041 140175
rect 231069 140147 231104 140175
rect 230944 140113 231104 140147
rect 230944 140085 230979 140113
rect 231007 140085 231041 140113
rect 231069 140085 231104 140113
rect 230944 140051 231104 140085
rect 230944 140023 230979 140051
rect 231007 140023 231041 140051
rect 231069 140023 231104 140051
rect 230944 139989 231104 140023
rect 230944 139961 230979 139989
rect 231007 139961 231041 139989
rect 231069 139961 231104 139989
rect 230944 139944 231104 139961
rect 223264 137175 223424 137192
rect 223264 137147 223299 137175
rect 223327 137147 223361 137175
rect 223389 137147 223424 137175
rect 223264 137113 223424 137147
rect 223264 137085 223299 137113
rect 223327 137085 223361 137113
rect 223389 137085 223424 137113
rect 223264 137051 223424 137085
rect 223264 137023 223299 137051
rect 223327 137023 223361 137051
rect 223389 137023 223424 137051
rect 223264 136989 223424 137023
rect 223264 136961 223299 136989
rect 223327 136961 223361 136989
rect 223389 136961 223424 136989
rect 223264 136944 223424 136961
rect 233109 137175 233419 145961
rect 233109 137147 233157 137175
rect 233185 137147 233219 137175
rect 233247 137147 233281 137175
rect 233309 137147 233343 137175
rect 233371 137147 233419 137175
rect 233109 137113 233419 137147
rect 233109 137085 233157 137113
rect 233185 137085 233219 137113
rect 233247 137085 233281 137113
rect 233309 137085 233343 137113
rect 233371 137085 233419 137113
rect 233109 137051 233419 137085
rect 233109 137023 233157 137051
rect 233185 137023 233219 137051
rect 233247 137023 233281 137051
rect 233309 137023 233343 137051
rect 233371 137023 233419 137051
rect 233109 136989 233419 137023
rect 233109 136961 233157 136989
rect 233185 136961 233219 136989
rect 233247 136961 233281 136989
rect 233309 136961 233343 136989
rect 233371 136961 233419 136989
rect 219609 131147 219657 131175
rect 219685 131147 219719 131175
rect 219747 131147 219781 131175
rect 219809 131147 219843 131175
rect 219871 131147 219919 131175
rect 219609 131113 219919 131147
rect 219609 131085 219657 131113
rect 219685 131085 219719 131113
rect 219747 131085 219781 131113
rect 219809 131085 219843 131113
rect 219871 131085 219919 131113
rect 219609 131051 219919 131085
rect 219609 131023 219657 131051
rect 219685 131023 219719 131051
rect 219747 131023 219781 131051
rect 219809 131023 219843 131051
rect 219871 131023 219919 131051
rect 219609 130989 219919 131023
rect 219609 130961 219657 130989
rect 219685 130961 219719 130989
rect 219747 130961 219781 130989
rect 219809 130961 219843 130989
rect 219871 130961 219919 130989
rect 219609 122175 219919 130961
rect 230944 131175 231104 131192
rect 230944 131147 230979 131175
rect 231007 131147 231041 131175
rect 231069 131147 231104 131175
rect 230944 131113 231104 131147
rect 230944 131085 230979 131113
rect 231007 131085 231041 131113
rect 231069 131085 231104 131113
rect 230944 131051 231104 131085
rect 230944 131023 230979 131051
rect 231007 131023 231041 131051
rect 231069 131023 231104 131051
rect 230944 130989 231104 131023
rect 230944 130961 230979 130989
rect 231007 130961 231041 130989
rect 231069 130961 231104 130989
rect 230944 130944 231104 130961
rect 223264 128175 223424 128192
rect 223264 128147 223299 128175
rect 223327 128147 223361 128175
rect 223389 128147 223424 128175
rect 223264 128113 223424 128147
rect 223264 128085 223299 128113
rect 223327 128085 223361 128113
rect 223389 128085 223424 128113
rect 223264 128051 223424 128085
rect 223264 128023 223299 128051
rect 223327 128023 223361 128051
rect 223389 128023 223424 128051
rect 223264 127989 223424 128023
rect 223264 127961 223299 127989
rect 223327 127961 223361 127989
rect 223389 127961 223424 127989
rect 223264 127944 223424 127961
rect 233109 128175 233419 136961
rect 233109 128147 233157 128175
rect 233185 128147 233219 128175
rect 233247 128147 233281 128175
rect 233309 128147 233343 128175
rect 233371 128147 233419 128175
rect 233109 128113 233419 128147
rect 233109 128085 233157 128113
rect 233185 128085 233219 128113
rect 233247 128085 233281 128113
rect 233309 128085 233343 128113
rect 233371 128085 233419 128113
rect 233109 128051 233419 128085
rect 233109 128023 233157 128051
rect 233185 128023 233219 128051
rect 233247 128023 233281 128051
rect 233309 128023 233343 128051
rect 233371 128023 233419 128051
rect 233109 127989 233419 128023
rect 233109 127961 233157 127989
rect 233185 127961 233219 127989
rect 233247 127961 233281 127989
rect 233309 127961 233343 127989
rect 233371 127961 233419 127989
rect 219609 122147 219657 122175
rect 219685 122147 219719 122175
rect 219747 122147 219781 122175
rect 219809 122147 219843 122175
rect 219871 122147 219919 122175
rect 219609 122113 219919 122147
rect 219609 122085 219657 122113
rect 219685 122085 219719 122113
rect 219747 122085 219781 122113
rect 219809 122085 219843 122113
rect 219871 122085 219919 122113
rect 219609 122051 219919 122085
rect 219609 122023 219657 122051
rect 219685 122023 219719 122051
rect 219747 122023 219781 122051
rect 219809 122023 219843 122051
rect 219871 122023 219919 122051
rect 219609 121989 219919 122023
rect 219609 121961 219657 121989
rect 219685 121961 219719 121989
rect 219747 121961 219781 121989
rect 219809 121961 219843 121989
rect 219871 121961 219919 121989
rect 219609 113175 219919 121961
rect 230944 122175 231104 122192
rect 230944 122147 230979 122175
rect 231007 122147 231041 122175
rect 231069 122147 231104 122175
rect 230944 122113 231104 122147
rect 230944 122085 230979 122113
rect 231007 122085 231041 122113
rect 231069 122085 231104 122113
rect 230944 122051 231104 122085
rect 230944 122023 230979 122051
rect 231007 122023 231041 122051
rect 231069 122023 231104 122051
rect 230944 121989 231104 122023
rect 230944 121961 230979 121989
rect 231007 121961 231041 121989
rect 231069 121961 231104 121989
rect 230944 121944 231104 121961
rect 223264 119175 223424 119192
rect 223264 119147 223299 119175
rect 223327 119147 223361 119175
rect 223389 119147 223424 119175
rect 223264 119113 223424 119147
rect 223264 119085 223299 119113
rect 223327 119085 223361 119113
rect 223389 119085 223424 119113
rect 223264 119051 223424 119085
rect 223264 119023 223299 119051
rect 223327 119023 223361 119051
rect 223389 119023 223424 119051
rect 223264 118989 223424 119023
rect 223264 118961 223299 118989
rect 223327 118961 223361 118989
rect 223389 118961 223424 118989
rect 223264 118944 223424 118961
rect 233109 119175 233419 127961
rect 233109 119147 233157 119175
rect 233185 119147 233219 119175
rect 233247 119147 233281 119175
rect 233309 119147 233343 119175
rect 233371 119147 233419 119175
rect 233109 119113 233419 119147
rect 233109 119085 233157 119113
rect 233185 119085 233219 119113
rect 233247 119085 233281 119113
rect 233309 119085 233343 119113
rect 233371 119085 233419 119113
rect 233109 119051 233419 119085
rect 233109 119023 233157 119051
rect 233185 119023 233219 119051
rect 233247 119023 233281 119051
rect 233309 119023 233343 119051
rect 233371 119023 233419 119051
rect 233109 118989 233419 119023
rect 233109 118961 233157 118989
rect 233185 118961 233219 118989
rect 233247 118961 233281 118989
rect 233309 118961 233343 118989
rect 233371 118961 233419 118989
rect 219609 113147 219657 113175
rect 219685 113147 219719 113175
rect 219747 113147 219781 113175
rect 219809 113147 219843 113175
rect 219871 113147 219919 113175
rect 219609 113113 219919 113147
rect 219609 113085 219657 113113
rect 219685 113085 219719 113113
rect 219747 113085 219781 113113
rect 219809 113085 219843 113113
rect 219871 113085 219919 113113
rect 219609 113051 219919 113085
rect 219609 113023 219657 113051
rect 219685 113023 219719 113051
rect 219747 113023 219781 113051
rect 219809 113023 219843 113051
rect 219871 113023 219919 113051
rect 219609 112989 219919 113023
rect 219609 112961 219657 112989
rect 219685 112961 219719 112989
rect 219747 112961 219781 112989
rect 219809 112961 219843 112989
rect 219871 112961 219919 112989
rect 219609 104175 219919 112961
rect 230944 113175 231104 113192
rect 230944 113147 230979 113175
rect 231007 113147 231041 113175
rect 231069 113147 231104 113175
rect 230944 113113 231104 113147
rect 230944 113085 230979 113113
rect 231007 113085 231041 113113
rect 231069 113085 231104 113113
rect 230944 113051 231104 113085
rect 230944 113023 230979 113051
rect 231007 113023 231041 113051
rect 231069 113023 231104 113051
rect 230944 112989 231104 113023
rect 230944 112961 230979 112989
rect 231007 112961 231041 112989
rect 231069 112961 231104 112989
rect 230944 112944 231104 112961
rect 223264 110175 223424 110192
rect 223264 110147 223299 110175
rect 223327 110147 223361 110175
rect 223389 110147 223424 110175
rect 223264 110113 223424 110147
rect 223264 110085 223299 110113
rect 223327 110085 223361 110113
rect 223389 110085 223424 110113
rect 223264 110051 223424 110085
rect 223264 110023 223299 110051
rect 223327 110023 223361 110051
rect 223389 110023 223424 110051
rect 223264 109989 223424 110023
rect 223264 109961 223299 109989
rect 223327 109961 223361 109989
rect 223389 109961 223424 109989
rect 223264 109944 223424 109961
rect 233109 110175 233419 118961
rect 233109 110147 233157 110175
rect 233185 110147 233219 110175
rect 233247 110147 233281 110175
rect 233309 110147 233343 110175
rect 233371 110147 233419 110175
rect 233109 110113 233419 110147
rect 233109 110085 233157 110113
rect 233185 110085 233219 110113
rect 233247 110085 233281 110113
rect 233309 110085 233343 110113
rect 233371 110085 233419 110113
rect 233109 110051 233419 110085
rect 233109 110023 233157 110051
rect 233185 110023 233219 110051
rect 233247 110023 233281 110051
rect 233309 110023 233343 110051
rect 233371 110023 233419 110051
rect 233109 109989 233419 110023
rect 233109 109961 233157 109989
rect 233185 109961 233219 109989
rect 233247 109961 233281 109989
rect 233309 109961 233343 109989
rect 233371 109961 233419 109989
rect 219609 104147 219657 104175
rect 219685 104147 219719 104175
rect 219747 104147 219781 104175
rect 219809 104147 219843 104175
rect 219871 104147 219919 104175
rect 219609 104113 219919 104147
rect 219609 104085 219657 104113
rect 219685 104085 219719 104113
rect 219747 104085 219781 104113
rect 219809 104085 219843 104113
rect 219871 104085 219919 104113
rect 219609 104051 219919 104085
rect 219609 104023 219657 104051
rect 219685 104023 219719 104051
rect 219747 104023 219781 104051
rect 219809 104023 219843 104051
rect 219871 104023 219919 104051
rect 219609 103989 219919 104023
rect 219609 103961 219657 103989
rect 219685 103961 219719 103989
rect 219747 103961 219781 103989
rect 219809 103961 219843 103989
rect 219871 103961 219919 103989
rect 219609 95175 219919 103961
rect 230944 104175 231104 104192
rect 230944 104147 230979 104175
rect 231007 104147 231041 104175
rect 231069 104147 231104 104175
rect 230944 104113 231104 104147
rect 230944 104085 230979 104113
rect 231007 104085 231041 104113
rect 231069 104085 231104 104113
rect 230944 104051 231104 104085
rect 230944 104023 230979 104051
rect 231007 104023 231041 104051
rect 231069 104023 231104 104051
rect 230944 103989 231104 104023
rect 230944 103961 230979 103989
rect 231007 103961 231041 103989
rect 231069 103961 231104 103989
rect 230944 103944 231104 103961
rect 223264 101175 223424 101192
rect 223264 101147 223299 101175
rect 223327 101147 223361 101175
rect 223389 101147 223424 101175
rect 223264 101113 223424 101147
rect 223264 101085 223299 101113
rect 223327 101085 223361 101113
rect 223389 101085 223424 101113
rect 223264 101051 223424 101085
rect 223264 101023 223299 101051
rect 223327 101023 223361 101051
rect 223389 101023 223424 101051
rect 223264 100989 223424 101023
rect 223264 100961 223299 100989
rect 223327 100961 223361 100989
rect 223389 100961 223424 100989
rect 223264 100944 223424 100961
rect 233109 101175 233419 109961
rect 233109 101147 233157 101175
rect 233185 101147 233219 101175
rect 233247 101147 233281 101175
rect 233309 101147 233343 101175
rect 233371 101147 233419 101175
rect 233109 101113 233419 101147
rect 233109 101085 233157 101113
rect 233185 101085 233219 101113
rect 233247 101085 233281 101113
rect 233309 101085 233343 101113
rect 233371 101085 233419 101113
rect 233109 101051 233419 101085
rect 233109 101023 233157 101051
rect 233185 101023 233219 101051
rect 233247 101023 233281 101051
rect 233309 101023 233343 101051
rect 233371 101023 233419 101051
rect 233109 100989 233419 101023
rect 233109 100961 233157 100989
rect 233185 100961 233219 100989
rect 233247 100961 233281 100989
rect 233309 100961 233343 100989
rect 233371 100961 233419 100989
rect 219609 95147 219657 95175
rect 219685 95147 219719 95175
rect 219747 95147 219781 95175
rect 219809 95147 219843 95175
rect 219871 95147 219919 95175
rect 219609 95113 219919 95147
rect 219609 95085 219657 95113
rect 219685 95085 219719 95113
rect 219747 95085 219781 95113
rect 219809 95085 219843 95113
rect 219871 95085 219919 95113
rect 219609 95051 219919 95085
rect 219609 95023 219657 95051
rect 219685 95023 219719 95051
rect 219747 95023 219781 95051
rect 219809 95023 219843 95051
rect 219871 95023 219919 95051
rect 219609 94989 219919 95023
rect 219609 94961 219657 94989
rect 219685 94961 219719 94989
rect 219747 94961 219781 94989
rect 219809 94961 219843 94989
rect 219871 94961 219919 94989
rect 219609 86175 219919 94961
rect 230944 95175 231104 95192
rect 230944 95147 230979 95175
rect 231007 95147 231041 95175
rect 231069 95147 231104 95175
rect 230944 95113 231104 95147
rect 230944 95085 230979 95113
rect 231007 95085 231041 95113
rect 231069 95085 231104 95113
rect 230944 95051 231104 95085
rect 230944 95023 230979 95051
rect 231007 95023 231041 95051
rect 231069 95023 231104 95051
rect 230944 94989 231104 95023
rect 230944 94961 230979 94989
rect 231007 94961 231041 94989
rect 231069 94961 231104 94989
rect 230944 94944 231104 94961
rect 223264 92175 223424 92192
rect 223264 92147 223299 92175
rect 223327 92147 223361 92175
rect 223389 92147 223424 92175
rect 223264 92113 223424 92147
rect 223264 92085 223299 92113
rect 223327 92085 223361 92113
rect 223389 92085 223424 92113
rect 223264 92051 223424 92085
rect 223264 92023 223299 92051
rect 223327 92023 223361 92051
rect 223389 92023 223424 92051
rect 223264 91989 223424 92023
rect 223264 91961 223299 91989
rect 223327 91961 223361 91989
rect 223389 91961 223424 91989
rect 223264 91944 223424 91961
rect 233109 92175 233419 100961
rect 233109 92147 233157 92175
rect 233185 92147 233219 92175
rect 233247 92147 233281 92175
rect 233309 92147 233343 92175
rect 233371 92147 233419 92175
rect 233109 92113 233419 92147
rect 233109 92085 233157 92113
rect 233185 92085 233219 92113
rect 233247 92085 233281 92113
rect 233309 92085 233343 92113
rect 233371 92085 233419 92113
rect 233109 92051 233419 92085
rect 233109 92023 233157 92051
rect 233185 92023 233219 92051
rect 233247 92023 233281 92051
rect 233309 92023 233343 92051
rect 233371 92023 233419 92051
rect 233109 91989 233419 92023
rect 233109 91961 233157 91989
rect 233185 91961 233219 91989
rect 233247 91961 233281 91989
rect 233309 91961 233343 91989
rect 233371 91961 233419 91989
rect 219609 86147 219657 86175
rect 219685 86147 219719 86175
rect 219747 86147 219781 86175
rect 219809 86147 219843 86175
rect 219871 86147 219919 86175
rect 219609 86113 219919 86147
rect 219609 86085 219657 86113
rect 219685 86085 219719 86113
rect 219747 86085 219781 86113
rect 219809 86085 219843 86113
rect 219871 86085 219919 86113
rect 219609 86051 219919 86085
rect 219609 86023 219657 86051
rect 219685 86023 219719 86051
rect 219747 86023 219781 86051
rect 219809 86023 219843 86051
rect 219871 86023 219919 86051
rect 219609 85989 219919 86023
rect 219609 85961 219657 85989
rect 219685 85961 219719 85989
rect 219747 85961 219781 85989
rect 219809 85961 219843 85989
rect 219871 85961 219919 85989
rect 219609 77175 219919 85961
rect 230944 86175 231104 86192
rect 230944 86147 230979 86175
rect 231007 86147 231041 86175
rect 231069 86147 231104 86175
rect 230944 86113 231104 86147
rect 230944 86085 230979 86113
rect 231007 86085 231041 86113
rect 231069 86085 231104 86113
rect 230944 86051 231104 86085
rect 230944 86023 230979 86051
rect 231007 86023 231041 86051
rect 231069 86023 231104 86051
rect 230944 85989 231104 86023
rect 230944 85961 230979 85989
rect 231007 85961 231041 85989
rect 231069 85961 231104 85989
rect 230944 85944 231104 85961
rect 223264 83175 223424 83192
rect 223264 83147 223299 83175
rect 223327 83147 223361 83175
rect 223389 83147 223424 83175
rect 223264 83113 223424 83147
rect 223264 83085 223299 83113
rect 223327 83085 223361 83113
rect 223389 83085 223424 83113
rect 223264 83051 223424 83085
rect 223264 83023 223299 83051
rect 223327 83023 223361 83051
rect 223389 83023 223424 83051
rect 223264 82989 223424 83023
rect 223264 82961 223299 82989
rect 223327 82961 223361 82989
rect 223389 82961 223424 82989
rect 223264 82944 223424 82961
rect 233109 83175 233419 91961
rect 233109 83147 233157 83175
rect 233185 83147 233219 83175
rect 233247 83147 233281 83175
rect 233309 83147 233343 83175
rect 233371 83147 233419 83175
rect 233109 83113 233419 83147
rect 233109 83085 233157 83113
rect 233185 83085 233219 83113
rect 233247 83085 233281 83113
rect 233309 83085 233343 83113
rect 233371 83085 233419 83113
rect 233109 83051 233419 83085
rect 233109 83023 233157 83051
rect 233185 83023 233219 83051
rect 233247 83023 233281 83051
rect 233309 83023 233343 83051
rect 233371 83023 233419 83051
rect 233109 82989 233419 83023
rect 233109 82961 233157 82989
rect 233185 82961 233219 82989
rect 233247 82961 233281 82989
rect 233309 82961 233343 82989
rect 233371 82961 233419 82989
rect 219609 77147 219657 77175
rect 219685 77147 219719 77175
rect 219747 77147 219781 77175
rect 219809 77147 219843 77175
rect 219871 77147 219919 77175
rect 219609 77113 219919 77147
rect 219609 77085 219657 77113
rect 219685 77085 219719 77113
rect 219747 77085 219781 77113
rect 219809 77085 219843 77113
rect 219871 77085 219919 77113
rect 219609 77051 219919 77085
rect 219609 77023 219657 77051
rect 219685 77023 219719 77051
rect 219747 77023 219781 77051
rect 219809 77023 219843 77051
rect 219871 77023 219919 77051
rect 219609 76989 219919 77023
rect 219609 76961 219657 76989
rect 219685 76961 219719 76989
rect 219747 76961 219781 76989
rect 219809 76961 219843 76989
rect 219871 76961 219919 76989
rect 219609 68175 219919 76961
rect 230944 77175 231104 77192
rect 230944 77147 230979 77175
rect 231007 77147 231041 77175
rect 231069 77147 231104 77175
rect 230944 77113 231104 77147
rect 230944 77085 230979 77113
rect 231007 77085 231041 77113
rect 231069 77085 231104 77113
rect 230944 77051 231104 77085
rect 230944 77023 230979 77051
rect 231007 77023 231041 77051
rect 231069 77023 231104 77051
rect 230944 76989 231104 77023
rect 230944 76961 230979 76989
rect 231007 76961 231041 76989
rect 231069 76961 231104 76989
rect 230944 76944 231104 76961
rect 223264 74175 223424 74192
rect 223264 74147 223299 74175
rect 223327 74147 223361 74175
rect 223389 74147 223424 74175
rect 223264 74113 223424 74147
rect 223264 74085 223299 74113
rect 223327 74085 223361 74113
rect 223389 74085 223424 74113
rect 223264 74051 223424 74085
rect 223264 74023 223299 74051
rect 223327 74023 223361 74051
rect 223389 74023 223424 74051
rect 223264 73989 223424 74023
rect 223264 73961 223299 73989
rect 223327 73961 223361 73989
rect 223389 73961 223424 73989
rect 223264 73944 223424 73961
rect 233109 74175 233419 82961
rect 233109 74147 233157 74175
rect 233185 74147 233219 74175
rect 233247 74147 233281 74175
rect 233309 74147 233343 74175
rect 233371 74147 233419 74175
rect 233109 74113 233419 74147
rect 233109 74085 233157 74113
rect 233185 74085 233219 74113
rect 233247 74085 233281 74113
rect 233309 74085 233343 74113
rect 233371 74085 233419 74113
rect 233109 74051 233419 74085
rect 233109 74023 233157 74051
rect 233185 74023 233219 74051
rect 233247 74023 233281 74051
rect 233309 74023 233343 74051
rect 233371 74023 233419 74051
rect 233109 73989 233419 74023
rect 233109 73961 233157 73989
rect 233185 73961 233219 73989
rect 233247 73961 233281 73989
rect 233309 73961 233343 73989
rect 233371 73961 233419 73989
rect 219609 68147 219657 68175
rect 219685 68147 219719 68175
rect 219747 68147 219781 68175
rect 219809 68147 219843 68175
rect 219871 68147 219919 68175
rect 219609 68113 219919 68147
rect 219609 68085 219657 68113
rect 219685 68085 219719 68113
rect 219747 68085 219781 68113
rect 219809 68085 219843 68113
rect 219871 68085 219919 68113
rect 219609 68051 219919 68085
rect 219609 68023 219657 68051
rect 219685 68023 219719 68051
rect 219747 68023 219781 68051
rect 219809 68023 219843 68051
rect 219871 68023 219919 68051
rect 219609 67989 219919 68023
rect 219609 67961 219657 67989
rect 219685 67961 219719 67989
rect 219747 67961 219781 67989
rect 219809 67961 219843 67989
rect 219871 67961 219919 67989
rect 219609 59175 219919 67961
rect 230944 68175 231104 68192
rect 230944 68147 230979 68175
rect 231007 68147 231041 68175
rect 231069 68147 231104 68175
rect 230944 68113 231104 68147
rect 230944 68085 230979 68113
rect 231007 68085 231041 68113
rect 231069 68085 231104 68113
rect 230944 68051 231104 68085
rect 230944 68023 230979 68051
rect 231007 68023 231041 68051
rect 231069 68023 231104 68051
rect 230944 67989 231104 68023
rect 230944 67961 230979 67989
rect 231007 67961 231041 67989
rect 231069 67961 231104 67989
rect 230944 67944 231104 67961
rect 223264 65175 223424 65192
rect 223264 65147 223299 65175
rect 223327 65147 223361 65175
rect 223389 65147 223424 65175
rect 223264 65113 223424 65147
rect 223264 65085 223299 65113
rect 223327 65085 223361 65113
rect 223389 65085 223424 65113
rect 223264 65051 223424 65085
rect 223264 65023 223299 65051
rect 223327 65023 223361 65051
rect 223389 65023 223424 65051
rect 223264 64989 223424 65023
rect 223264 64961 223299 64989
rect 223327 64961 223361 64989
rect 223389 64961 223424 64989
rect 223264 64944 223424 64961
rect 233109 65175 233419 73961
rect 233109 65147 233157 65175
rect 233185 65147 233219 65175
rect 233247 65147 233281 65175
rect 233309 65147 233343 65175
rect 233371 65147 233419 65175
rect 233109 65113 233419 65147
rect 233109 65085 233157 65113
rect 233185 65085 233219 65113
rect 233247 65085 233281 65113
rect 233309 65085 233343 65113
rect 233371 65085 233419 65113
rect 233109 65051 233419 65085
rect 233109 65023 233157 65051
rect 233185 65023 233219 65051
rect 233247 65023 233281 65051
rect 233309 65023 233343 65051
rect 233371 65023 233419 65051
rect 233109 64989 233419 65023
rect 233109 64961 233157 64989
rect 233185 64961 233219 64989
rect 233247 64961 233281 64989
rect 233309 64961 233343 64989
rect 233371 64961 233419 64989
rect 219609 59147 219657 59175
rect 219685 59147 219719 59175
rect 219747 59147 219781 59175
rect 219809 59147 219843 59175
rect 219871 59147 219919 59175
rect 219609 59113 219919 59147
rect 219609 59085 219657 59113
rect 219685 59085 219719 59113
rect 219747 59085 219781 59113
rect 219809 59085 219843 59113
rect 219871 59085 219919 59113
rect 219609 59051 219919 59085
rect 219609 59023 219657 59051
rect 219685 59023 219719 59051
rect 219747 59023 219781 59051
rect 219809 59023 219843 59051
rect 219871 59023 219919 59051
rect 219609 58989 219919 59023
rect 219609 58961 219657 58989
rect 219685 58961 219719 58989
rect 219747 58961 219781 58989
rect 219809 58961 219843 58989
rect 219871 58961 219919 58989
rect 219609 50175 219919 58961
rect 230944 59175 231104 59192
rect 230944 59147 230979 59175
rect 231007 59147 231041 59175
rect 231069 59147 231104 59175
rect 230944 59113 231104 59147
rect 230944 59085 230979 59113
rect 231007 59085 231041 59113
rect 231069 59085 231104 59113
rect 230944 59051 231104 59085
rect 230944 59023 230979 59051
rect 231007 59023 231041 59051
rect 231069 59023 231104 59051
rect 230944 58989 231104 59023
rect 230944 58961 230979 58989
rect 231007 58961 231041 58989
rect 231069 58961 231104 58989
rect 230944 58944 231104 58961
rect 223264 56175 223424 56192
rect 223264 56147 223299 56175
rect 223327 56147 223361 56175
rect 223389 56147 223424 56175
rect 223264 56113 223424 56147
rect 223264 56085 223299 56113
rect 223327 56085 223361 56113
rect 223389 56085 223424 56113
rect 223264 56051 223424 56085
rect 223264 56023 223299 56051
rect 223327 56023 223361 56051
rect 223389 56023 223424 56051
rect 223264 55989 223424 56023
rect 223264 55961 223299 55989
rect 223327 55961 223361 55989
rect 223389 55961 223424 55989
rect 223264 55944 223424 55961
rect 233109 56175 233419 64961
rect 233109 56147 233157 56175
rect 233185 56147 233219 56175
rect 233247 56147 233281 56175
rect 233309 56147 233343 56175
rect 233371 56147 233419 56175
rect 233109 56113 233419 56147
rect 233109 56085 233157 56113
rect 233185 56085 233219 56113
rect 233247 56085 233281 56113
rect 233309 56085 233343 56113
rect 233371 56085 233419 56113
rect 233109 56051 233419 56085
rect 233109 56023 233157 56051
rect 233185 56023 233219 56051
rect 233247 56023 233281 56051
rect 233309 56023 233343 56051
rect 233371 56023 233419 56051
rect 233109 55989 233419 56023
rect 233109 55961 233157 55989
rect 233185 55961 233219 55989
rect 233247 55961 233281 55989
rect 233309 55961 233343 55989
rect 233371 55961 233419 55989
rect 219609 50147 219657 50175
rect 219685 50147 219719 50175
rect 219747 50147 219781 50175
rect 219809 50147 219843 50175
rect 219871 50147 219919 50175
rect 219609 50113 219919 50147
rect 219609 50085 219657 50113
rect 219685 50085 219719 50113
rect 219747 50085 219781 50113
rect 219809 50085 219843 50113
rect 219871 50085 219919 50113
rect 219609 50051 219919 50085
rect 219609 50023 219657 50051
rect 219685 50023 219719 50051
rect 219747 50023 219781 50051
rect 219809 50023 219843 50051
rect 219871 50023 219919 50051
rect 219609 49989 219919 50023
rect 219609 49961 219657 49989
rect 219685 49961 219719 49989
rect 219747 49961 219781 49989
rect 219809 49961 219843 49989
rect 219871 49961 219919 49989
rect 219609 41175 219919 49961
rect 230944 50175 231104 50192
rect 230944 50147 230979 50175
rect 231007 50147 231041 50175
rect 231069 50147 231104 50175
rect 230944 50113 231104 50147
rect 230944 50085 230979 50113
rect 231007 50085 231041 50113
rect 231069 50085 231104 50113
rect 230944 50051 231104 50085
rect 230944 50023 230979 50051
rect 231007 50023 231041 50051
rect 231069 50023 231104 50051
rect 230944 49989 231104 50023
rect 230944 49961 230979 49989
rect 231007 49961 231041 49989
rect 231069 49961 231104 49989
rect 230944 49944 231104 49961
rect 223264 47175 223424 47192
rect 223264 47147 223299 47175
rect 223327 47147 223361 47175
rect 223389 47147 223424 47175
rect 223264 47113 223424 47147
rect 223264 47085 223299 47113
rect 223327 47085 223361 47113
rect 223389 47085 223424 47113
rect 223264 47051 223424 47085
rect 223264 47023 223299 47051
rect 223327 47023 223361 47051
rect 223389 47023 223424 47051
rect 223264 46989 223424 47023
rect 223264 46961 223299 46989
rect 223327 46961 223361 46989
rect 223389 46961 223424 46989
rect 223264 46944 223424 46961
rect 233109 47175 233419 55961
rect 233109 47147 233157 47175
rect 233185 47147 233219 47175
rect 233247 47147 233281 47175
rect 233309 47147 233343 47175
rect 233371 47147 233419 47175
rect 233109 47113 233419 47147
rect 233109 47085 233157 47113
rect 233185 47085 233219 47113
rect 233247 47085 233281 47113
rect 233309 47085 233343 47113
rect 233371 47085 233419 47113
rect 233109 47051 233419 47085
rect 233109 47023 233157 47051
rect 233185 47023 233219 47051
rect 233247 47023 233281 47051
rect 233309 47023 233343 47051
rect 233371 47023 233419 47051
rect 233109 46989 233419 47023
rect 233109 46961 233157 46989
rect 233185 46961 233219 46989
rect 233247 46961 233281 46989
rect 233309 46961 233343 46989
rect 233371 46961 233419 46989
rect 219609 41147 219657 41175
rect 219685 41147 219719 41175
rect 219747 41147 219781 41175
rect 219809 41147 219843 41175
rect 219871 41147 219919 41175
rect 219609 41113 219919 41147
rect 219609 41085 219657 41113
rect 219685 41085 219719 41113
rect 219747 41085 219781 41113
rect 219809 41085 219843 41113
rect 219871 41085 219919 41113
rect 219609 41051 219919 41085
rect 219609 41023 219657 41051
rect 219685 41023 219719 41051
rect 219747 41023 219781 41051
rect 219809 41023 219843 41051
rect 219871 41023 219919 41051
rect 219609 40989 219919 41023
rect 219609 40961 219657 40989
rect 219685 40961 219719 40989
rect 219747 40961 219781 40989
rect 219809 40961 219843 40989
rect 219871 40961 219919 40989
rect 219609 32175 219919 40961
rect 230944 41175 231104 41192
rect 230944 41147 230979 41175
rect 231007 41147 231041 41175
rect 231069 41147 231104 41175
rect 230944 41113 231104 41147
rect 230944 41085 230979 41113
rect 231007 41085 231041 41113
rect 231069 41085 231104 41113
rect 230944 41051 231104 41085
rect 230944 41023 230979 41051
rect 231007 41023 231041 41051
rect 231069 41023 231104 41051
rect 230944 40989 231104 41023
rect 230944 40961 230979 40989
rect 231007 40961 231041 40989
rect 231069 40961 231104 40989
rect 230944 40944 231104 40961
rect 223264 38175 223424 38192
rect 223264 38147 223299 38175
rect 223327 38147 223361 38175
rect 223389 38147 223424 38175
rect 223264 38113 223424 38147
rect 223264 38085 223299 38113
rect 223327 38085 223361 38113
rect 223389 38085 223424 38113
rect 223264 38051 223424 38085
rect 223264 38023 223299 38051
rect 223327 38023 223361 38051
rect 223389 38023 223424 38051
rect 223264 37989 223424 38023
rect 223264 37961 223299 37989
rect 223327 37961 223361 37989
rect 223389 37961 223424 37989
rect 223264 37944 223424 37961
rect 233109 38175 233419 46961
rect 233109 38147 233157 38175
rect 233185 38147 233219 38175
rect 233247 38147 233281 38175
rect 233309 38147 233343 38175
rect 233371 38147 233419 38175
rect 233109 38113 233419 38147
rect 233109 38085 233157 38113
rect 233185 38085 233219 38113
rect 233247 38085 233281 38113
rect 233309 38085 233343 38113
rect 233371 38085 233419 38113
rect 233109 38051 233419 38085
rect 233109 38023 233157 38051
rect 233185 38023 233219 38051
rect 233247 38023 233281 38051
rect 233309 38023 233343 38051
rect 233371 38023 233419 38051
rect 233109 37989 233419 38023
rect 233109 37961 233157 37989
rect 233185 37961 233219 37989
rect 233247 37961 233281 37989
rect 233309 37961 233343 37989
rect 233371 37961 233419 37989
rect 219609 32147 219657 32175
rect 219685 32147 219719 32175
rect 219747 32147 219781 32175
rect 219809 32147 219843 32175
rect 219871 32147 219919 32175
rect 219609 32113 219919 32147
rect 219609 32085 219657 32113
rect 219685 32085 219719 32113
rect 219747 32085 219781 32113
rect 219809 32085 219843 32113
rect 219871 32085 219919 32113
rect 219609 32051 219919 32085
rect 219609 32023 219657 32051
rect 219685 32023 219719 32051
rect 219747 32023 219781 32051
rect 219809 32023 219843 32051
rect 219871 32023 219919 32051
rect 219609 31989 219919 32023
rect 219609 31961 219657 31989
rect 219685 31961 219719 31989
rect 219747 31961 219781 31989
rect 219809 31961 219843 31989
rect 219871 31961 219919 31989
rect 219609 23175 219919 31961
rect 230944 32175 231104 32192
rect 230944 32147 230979 32175
rect 231007 32147 231041 32175
rect 231069 32147 231104 32175
rect 230944 32113 231104 32147
rect 230944 32085 230979 32113
rect 231007 32085 231041 32113
rect 231069 32085 231104 32113
rect 230944 32051 231104 32085
rect 230944 32023 230979 32051
rect 231007 32023 231041 32051
rect 231069 32023 231104 32051
rect 230944 31989 231104 32023
rect 230944 31961 230979 31989
rect 231007 31961 231041 31989
rect 231069 31961 231104 31989
rect 230944 31944 231104 31961
rect 223264 29175 223424 29192
rect 223264 29147 223299 29175
rect 223327 29147 223361 29175
rect 223389 29147 223424 29175
rect 223264 29113 223424 29147
rect 223264 29085 223299 29113
rect 223327 29085 223361 29113
rect 223389 29085 223424 29113
rect 223264 29051 223424 29085
rect 223264 29023 223299 29051
rect 223327 29023 223361 29051
rect 223389 29023 223424 29051
rect 223264 28989 223424 29023
rect 223264 28961 223299 28989
rect 223327 28961 223361 28989
rect 223389 28961 223424 28989
rect 223264 28944 223424 28961
rect 233109 29175 233419 37961
rect 233109 29147 233157 29175
rect 233185 29147 233219 29175
rect 233247 29147 233281 29175
rect 233309 29147 233343 29175
rect 233371 29147 233419 29175
rect 233109 29113 233419 29147
rect 233109 29085 233157 29113
rect 233185 29085 233219 29113
rect 233247 29085 233281 29113
rect 233309 29085 233343 29113
rect 233371 29085 233419 29113
rect 233109 29051 233419 29085
rect 233109 29023 233157 29051
rect 233185 29023 233219 29051
rect 233247 29023 233281 29051
rect 233309 29023 233343 29051
rect 233371 29023 233419 29051
rect 233109 28989 233419 29023
rect 233109 28961 233157 28989
rect 233185 28961 233219 28989
rect 233247 28961 233281 28989
rect 233309 28961 233343 28989
rect 233371 28961 233419 28989
rect 219609 23147 219657 23175
rect 219685 23147 219719 23175
rect 219747 23147 219781 23175
rect 219809 23147 219843 23175
rect 219871 23147 219919 23175
rect 219609 23113 219919 23147
rect 219609 23085 219657 23113
rect 219685 23085 219719 23113
rect 219747 23085 219781 23113
rect 219809 23085 219843 23113
rect 219871 23085 219919 23113
rect 219609 23051 219919 23085
rect 219609 23023 219657 23051
rect 219685 23023 219719 23051
rect 219747 23023 219781 23051
rect 219809 23023 219843 23051
rect 219871 23023 219919 23051
rect 219609 22989 219919 23023
rect 219609 22961 219657 22989
rect 219685 22961 219719 22989
rect 219747 22961 219781 22989
rect 219809 22961 219843 22989
rect 219871 22961 219919 22989
rect 219609 14175 219919 22961
rect 230944 23175 231104 23192
rect 230944 23147 230979 23175
rect 231007 23147 231041 23175
rect 231069 23147 231104 23175
rect 230944 23113 231104 23147
rect 230944 23085 230979 23113
rect 231007 23085 231041 23113
rect 231069 23085 231104 23113
rect 230944 23051 231104 23085
rect 230944 23023 230979 23051
rect 231007 23023 231041 23051
rect 231069 23023 231104 23051
rect 230944 22989 231104 23023
rect 230944 22961 230979 22989
rect 231007 22961 231041 22989
rect 231069 22961 231104 22989
rect 230944 22944 231104 22961
rect 223264 20175 223424 20192
rect 223264 20147 223299 20175
rect 223327 20147 223361 20175
rect 223389 20147 223424 20175
rect 223264 20113 223424 20147
rect 223264 20085 223299 20113
rect 223327 20085 223361 20113
rect 223389 20085 223424 20113
rect 223264 20051 223424 20085
rect 223264 20023 223299 20051
rect 223327 20023 223361 20051
rect 223389 20023 223424 20051
rect 223264 19989 223424 20023
rect 223264 19961 223299 19989
rect 223327 19961 223361 19989
rect 223389 19961 223424 19989
rect 223264 19944 223424 19961
rect 233109 20175 233419 28961
rect 233109 20147 233157 20175
rect 233185 20147 233219 20175
rect 233247 20147 233281 20175
rect 233309 20147 233343 20175
rect 233371 20147 233419 20175
rect 233109 20113 233419 20147
rect 233109 20085 233157 20113
rect 233185 20085 233219 20113
rect 233247 20085 233281 20113
rect 233309 20085 233343 20113
rect 233371 20085 233419 20113
rect 233109 20051 233419 20085
rect 233109 20023 233157 20051
rect 233185 20023 233219 20051
rect 233247 20023 233281 20051
rect 233309 20023 233343 20051
rect 233371 20023 233419 20051
rect 233109 19989 233419 20023
rect 233109 19961 233157 19989
rect 233185 19961 233219 19989
rect 233247 19961 233281 19989
rect 233309 19961 233343 19989
rect 233371 19961 233419 19989
rect 219609 14147 219657 14175
rect 219685 14147 219719 14175
rect 219747 14147 219781 14175
rect 219809 14147 219843 14175
rect 219871 14147 219919 14175
rect 219609 14113 219919 14147
rect 219609 14085 219657 14113
rect 219685 14085 219719 14113
rect 219747 14085 219781 14113
rect 219809 14085 219843 14113
rect 219871 14085 219919 14113
rect 219609 14051 219919 14085
rect 219609 14023 219657 14051
rect 219685 14023 219719 14051
rect 219747 14023 219781 14051
rect 219809 14023 219843 14051
rect 219871 14023 219919 14051
rect 219609 13989 219919 14023
rect 219609 13961 219657 13989
rect 219685 13961 219719 13989
rect 219747 13961 219781 13989
rect 219809 13961 219843 13989
rect 219871 13961 219919 13989
rect 219609 5175 219919 13961
rect 230944 14175 231104 14192
rect 230944 14147 230979 14175
rect 231007 14147 231041 14175
rect 231069 14147 231104 14175
rect 230944 14113 231104 14147
rect 230944 14085 230979 14113
rect 231007 14085 231041 14113
rect 231069 14085 231104 14113
rect 230944 14051 231104 14085
rect 230944 14023 230979 14051
rect 231007 14023 231041 14051
rect 231069 14023 231104 14051
rect 230944 13989 231104 14023
rect 230944 13961 230979 13989
rect 231007 13961 231041 13989
rect 231069 13961 231104 13989
rect 230944 13944 231104 13961
rect 223264 11175 223424 11192
rect 223264 11147 223299 11175
rect 223327 11147 223361 11175
rect 223389 11147 223424 11175
rect 223264 11113 223424 11147
rect 223264 11085 223299 11113
rect 223327 11085 223361 11113
rect 223389 11085 223424 11113
rect 223264 11051 223424 11085
rect 223264 11023 223299 11051
rect 223327 11023 223361 11051
rect 223389 11023 223424 11051
rect 223264 10989 223424 11023
rect 223264 10961 223299 10989
rect 223327 10961 223361 10989
rect 223389 10961 223424 10989
rect 223264 10944 223424 10961
rect 233109 11175 233419 19961
rect 233109 11147 233157 11175
rect 233185 11147 233219 11175
rect 233247 11147 233281 11175
rect 233309 11147 233343 11175
rect 233371 11147 233419 11175
rect 233109 11113 233419 11147
rect 233109 11085 233157 11113
rect 233185 11085 233219 11113
rect 233247 11085 233281 11113
rect 233309 11085 233343 11113
rect 233371 11085 233419 11113
rect 233109 11051 233419 11085
rect 233109 11023 233157 11051
rect 233185 11023 233219 11051
rect 233247 11023 233281 11051
rect 233309 11023 233343 11051
rect 233371 11023 233419 11051
rect 233109 10989 233419 11023
rect 233109 10961 233157 10989
rect 233185 10961 233219 10989
rect 233247 10961 233281 10989
rect 233309 10961 233343 10989
rect 233371 10961 233419 10989
rect 219609 5147 219657 5175
rect 219685 5147 219719 5175
rect 219747 5147 219781 5175
rect 219809 5147 219843 5175
rect 219871 5147 219919 5175
rect 219609 5113 219919 5147
rect 219609 5085 219657 5113
rect 219685 5085 219719 5113
rect 219747 5085 219781 5113
rect 219809 5085 219843 5113
rect 219871 5085 219919 5113
rect 219609 5051 219919 5085
rect 219609 5023 219657 5051
rect 219685 5023 219719 5051
rect 219747 5023 219781 5051
rect 219809 5023 219843 5051
rect 219871 5023 219919 5051
rect 219609 4989 219919 5023
rect 219609 4961 219657 4989
rect 219685 4961 219719 4989
rect 219747 4961 219781 4989
rect 219809 4961 219843 4989
rect 219871 4961 219919 4989
rect 219609 -560 219919 4961
rect 230944 5175 231104 5192
rect 230944 5147 230979 5175
rect 231007 5147 231041 5175
rect 231069 5147 231104 5175
rect 230944 5113 231104 5147
rect 230944 5085 230979 5113
rect 231007 5085 231041 5113
rect 231069 5085 231104 5113
rect 230944 5051 231104 5085
rect 230944 5023 230979 5051
rect 231007 5023 231041 5051
rect 231069 5023 231104 5051
rect 230944 4989 231104 5023
rect 230944 4961 230979 4989
rect 231007 4961 231041 4989
rect 231069 4961 231104 4989
rect 230944 4944 231104 4961
rect 219609 -588 219657 -560
rect 219685 -588 219719 -560
rect 219747 -588 219781 -560
rect 219809 -588 219843 -560
rect 219871 -588 219919 -560
rect 219609 -622 219919 -588
rect 219609 -650 219657 -622
rect 219685 -650 219719 -622
rect 219747 -650 219781 -622
rect 219809 -650 219843 -622
rect 219871 -650 219919 -622
rect 219609 -684 219919 -650
rect 219609 -712 219657 -684
rect 219685 -712 219719 -684
rect 219747 -712 219781 -684
rect 219809 -712 219843 -684
rect 219871 -712 219919 -684
rect 219609 -746 219919 -712
rect 219609 -774 219657 -746
rect 219685 -774 219719 -746
rect 219747 -774 219781 -746
rect 219809 -774 219843 -746
rect 219871 -774 219919 -746
rect 219609 -822 219919 -774
rect 233109 2175 233419 10961
rect 233109 2147 233157 2175
rect 233185 2147 233219 2175
rect 233247 2147 233281 2175
rect 233309 2147 233343 2175
rect 233371 2147 233419 2175
rect 233109 2113 233419 2147
rect 233109 2085 233157 2113
rect 233185 2085 233219 2113
rect 233247 2085 233281 2113
rect 233309 2085 233343 2113
rect 233371 2085 233419 2113
rect 233109 2051 233419 2085
rect 233109 2023 233157 2051
rect 233185 2023 233219 2051
rect 233247 2023 233281 2051
rect 233309 2023 233343 2051
rect 233371 2023 233419 2051
rect 233109 1989 233419 2023
rect 233109 1961 233157 1989
rect 233185 1961 233219 1989
rect 233247 1961 233281 1989
rect 233309 1961 233343 1989
rect 233371 1961 233419 1989
rect 233109 -80 233419 1961
rect 233109 -108 233157 -80
rect 233185 -108 233219 -80
rect 233247 -108 233281 -80
rect 233309 -108 233343 -80
rect 233371 -108 233419 -80
rect 233109 -142 233419 -108
rect 233109 -170 233157 -142
rect 233185 -170 233219 -142
rect 233247 -170 233281 -142
rect 233309 -170 233343 -142
rect 233371 -170 233419 -142
rect 233109 -204 233419 -170
rect 233109 -232 233157 -204
rect 233185 -232 233219 -204
rect 233247 -232 233281 -204
rect 233309 -232 233343 -204
rect 233371 -232 233419 -204
rect 233109 -266 233419 -232
rect 233109 -294 233157 -266
rect 233185 -294 233219 -266
rect 233247 -294 233281 -266
rect 233309 -294 233343 -266
rect 233371 -294 233419 -266
rect 233109 -822 233419 -294
rect 234969 299086 235279 299134
rect 234969 299058 235017 299086
rect 235045 299058 235079 299086
rect 235107 299058 235141 299086
rect 235169 299058 235203 299086
rect 235231 299058 235279 299086
rect 234969 299024 235279 299058
rect 234969 298996 235017 299024
rect 235045 298996 235079 299024
rect 235107 298996 235141 299024
rect 235169 298996 235203 299024
rect 235231 298996 235279 299024
rect 234969 298962 235279 298996
rect 234969 298934 235017 298962
rect 235045 298934 235079 298962
rect 235107 298934 235141 298962
rect 235169 298934 235203 298962
rect 235231 298934 235279 298962
rect 234969 298900 235279 298934
rect 234969 298872 235017 298900
rect 235045 298872 235079 298900
rect 235107 298872 235141 298900
rect 235169 298872 235203 298900
rect 235231 298872 235279 298900
rect 234969 293175 235279 298872
rect 234969 293147 235017 293175
rect 235045 293147 235079 293175
rect 235107 293147 235141 293175
rect 235169 293147 235203 293175
rect 235231 293147 235279 293175
rect 234969 293113 235279 293147
rect 234969 293085 235017 293113
rect 235045 293085 235079 293113
rect 235107 293085 235141 293113
rect 235169 293085 235203 293113
rect 235231 293085 235279 293113
rect 234969 293051 235279 293085
rect 234969 293023 235017 293051
rect 235045 293023 235079 293051
rect 235107 293023 235141 293051
rect 235169 293023 235203 293051
rect 235231 293023 235279 293051
rect 234969 292989 235279 293023
rect 234969 292961 235017 292989
rect 235045 292961 235079 292989
rect 235107 292961 235141 292989
rect 235169 292961 235203 292989
rect 235231 292961 235279 292989
rect 234969 284175 235279 292961
rect 234969 284147 235017 284175
rect 235045 284147 235079 284175
rect 235107 284147 235141 284175
rect 235169 284147 235203 284175
rect 235231 284147 235279 284175
rect 234969 284113 235279 284147
rect 234969 284085 235017 284113
rect 235045 284085 235079 284113
rect 235107 284085 235141 284113
rect 235169 284085 235203 284113
rect 235231 284085 235279 284113
rect 234969 284051 235279 284085
rect 234969 284023 235017 284051
rect 235045 284023 235079 284051
rect 235107 284023 235141 284051
rect 235169 284023 235203 284051
rect 235231 284023 235279 284051
rect 234969 283989 235279 284023
rect 234969 283961 235017 283989
rect 235045 283961 235079 283989
rect 235107 283961 235141 283989
rect 235169 283961 235203 283989
rect 235231 283961 235279 283989
rect 234969 275175 235279 283961
rect 234969 275147 235017 275175
rect 235045 275147 235079 275175
rect 235107 275147 235141 275175
rect 235169 275147 235203 275175
rect 235231 275147 235279 275175
rect 234969 275113 235279 275147
rect 234969 275085 235017 275113
rect 235045 275085 235079 275113
rect 235107 275085 235141 275113
rect 235169 275085 235203 275113
rect 235231 275085 235279 275113
rect 234969 275051 235279 275085
rect 234969 275023 235017 275051
rect 235045 275023 235079 275051
rect 235107 275023 235141 275051
rect 235169 275023 235203 275051
rect 235231 275023 235279 275051
rect 234969 274989 235279 275023
rect 234969 274961 235017 274989
rect 235045 274961 235079 274989
rect 235107 274961 235141 274989
rect 235169 274961 235203 274989
rect 235231 274961 235279 274989
rect 234969 266175 235279 274961
rect 234969 266147 235017 266175
rect 235045 266147 235079 266175
rect 235107 266147 235141 266175
rect 235169 266147 235203 266175
rect 235231 266147 235279 266175
rect 234969 266113 235279 266147
rect 234969 266085 235017 266113
rect 235045 266085 235079 266113
rect 235107 266085 235141 266113
rect 235169 266085 235203 266113
rect 235231 266085 235279 266113
rect 234969 266051 235279 266085
rect 234969 266023 235017 266051
rect 235045 266023 235079 266051
rect 235107 266023 235141 266051
rect 235169 266023 235203 266051
rect 235231 266023 235279 266051
rect 234969 265989 235279 266023
rect 234969 265961 235017 265989
rect 235045 265961 235079 265989
rect 235107 265961 235141 265989
rect 235169 265961 235203 265989
rect 235231 265961 235279 265989
rect 234969 257175 235279 265961
rect 234969 257147 235017 257175
rect 235045 257147 235079 257175
rect 235107 257147 235141 257175
rect 235169 257147 235203 257175
rect 235231 257147 235279 257175
rect 234969 257113 235279 257147
rect 234969 257085 235017 257113
rect 235045 257085 235079 257113
rect 235107 257085 235141 257113
rect 235169 257085 235203 257113
rect 235231 257085 235279 257113
rect 234969 257051 235279 257085
rect 234969 257023 235017 257051
rect 235045 257023 235079 257051
rect 235107 257023 235141 257051
rect 235169 257023 235203 257051
rect 235231 257023 235279 257051
rect 234969 256989 235279 257023
rect 234969 256961 235017 256989
rect 235045 256961 235079 256989
rect 235107 256961 235141 256989
rect 235169 256961 235203 256989
rect 235231 256961 235279 256989
rect 234969 248175 235279 256961
rect 234969 248147 235017 248175
rect 235045 248147 235079 248175
rect 235107 248147 235141 248175
rect 235169 248147 235203 248175
rect 235231 248147 235279 248175
rect 234969 248113 235279 248147
rect 234969 248085 235017 248113
rect 235045 248085 235079 248113
rect 235107 248085 235141 248113
rect 235169 248085 235203 248113
rect 235231 248085 235279 248113
rect 234969 248051 235279 248085
rect 234969 248023 235017 248051
rect 235045 248023 235079 248051
rect 235107 248023 235141 248051
rect 235169 248023 235203 248051
rect 235231 248023 235279 248051
rect 234969 247989 235279 248023
rect 234969 247961 235017 247989
rect 235045 247961 235079 247989
rect 235107 247961 235141 247989
rect 235169 247961 235203 247989
rect 235231 247961 235279 247989
rect 234969 239175 235279 247961
rect 234969 239147 235017 239175
rect 235045 239147 235079 239175
rect 235107 239147 235141 239175
rect 235169 239147 235203 239175
rect 235231 239147 235279 239175
rect 234969 239113 235279 239147
rect 234969 239085 235017 239113
rect 235045 239085 235079 239113
rect 235107 239085 235141 239113
rect 235169 239085 235203 239113
rect 235231 239085 235279 239113
rect 234969 239051 235279 239085
rect 234969 239023 235017 239051
rect 235045 239023 235079 239051
rect 235107 239023 235141 239051
rect 235169 239023 235203 239051
rect 235231 239023 235279 239051
rect 234969 238989 235279 239023
rect 234969 238961 235017 238989
rect 235045 238961 235079 238989
rect 235107 238961 235141 238989
rect 235169 238961 235203 238989
rect 235231 238961 235279 238989
rect 234969 230175 235279 238961
rect 234969 230147 235017 230175
rect 235045 230147 235079 230175
rect 235107 230147 235141 230175
rect 235169 230147 235203 230175
rect 235231 230147 235279 230175
rect 234969 230113 235279 230147
rect 234969 230085 235017 230113
rect 235045 230085 235079 230113
rect 235107 230085 235141 230113
rect 235169 230085 235203 230113
rect 235231 230085 235279 230113
rect 234969 230051 235279 230085
rect 234969 230023 235017 230051
rect 235045 230023 235079 230051
rect 235107 230023 235141 230051
rect 235169 230023 235203 230051
rect 235231 230023 235279 230051
rect 234969 229989 235279 230023
rect 234969 229961 235017 229989
rect 235045 229961 235079 229989
rect 235107 229961 235141 229989
rect 235169 229961 235203 229989
rect 235231 229961 235279 229989
rect 234969 221175 235279 229961
rect 234969 221147 235017 221175
rect 235045 221147 235079 221175
rect 235107 221147 235141 221175
rect 235169 221147 235203 221175
rect 235231 221147 235279 221175
rect 234969 221113 235279 221147
rect 234969 221085 235017 221113
rect 235045 221085 235079 221113
rect 235107 221085 235141 221113
rect 235169 221085 235203 221113
rect 235231 221085 235279 221113
rect 234969 221051 235279 221085
rect 234969 221023 235017 221051
rect 235045 221023 235079 221051
rect 235107 221023 235141 221051
rect 235169 221023 235203 221051
rect 235231 221023 235279 221051
rect 234969 220989 235279 221023
rect 234969 220961 235017 220989
rect 235045 220961 235079 220989
rect 235107 220961 235141 220989
rect 235169 220961 235203 220989
rect 235231 220961 235279 220989
rect 234969 212175 235279 220961
rect 234969 212147 235017 212175
rect 235045 212147 235079 212175
rect 235107 212147 235141 212175
rect 235169 212147 235203 212175
rect 235231 212147 235279 212175
rect 234969 212113 235279 212147
rect 234969 212085 235017 212113
rect 235045 212085 235079 212113
rect 235107 212085 235141 212113
rect 235169 212085 235203 212113
rect 235231 212085 235279 212113
rect 234969 212051 235279 212085
rect 234969 212023 235017 212051
rect 235045 212023 235079 212051
rect 235107 212023 235141 212051
rect 235169 212023 235203 212051
rect 235231 212023 235279 212051
rect 234969 211989 235279 212023
rect 234969 211961 235017 211989
rect 235045 211961 235079 211989
rect 235107 211961 235141 211989
rect 235169 211961 235203 211989
rect 235231 211961 235279 211989
rect 234969 203175 235279 211961
rect 234969 203147 235017 203175
rect 235045 203147 235079 203175
rect 235107 203147 235141 203175
rect 235169 203147 235203 203175
rect 235231 203147 235279 203175
rect 234969 203113 235279 203147
rect 234969 203085 235017 203113
rect 235045 203085 235079 203113
rect 235107 203085 235141 203113
rect 235169 203085 235203 203113
rect 235231 203085 235279 203113
rect 234969 203051 235279 203085
rect 234969 203023 235017 203051
rect 235045 203023 235079 203051
rect 235107 203023 235141 203051
rect 235169 203023 235203 203051
rect 235231 203023 235279 203051
rect 234969 202989 235279 203023
rect 234969 202961 235017 202989
rect 235045 202961 235079 202989
rect 235107 202961 235141 202989
rect 235169 202961 235203 202989
rect 235231 202961 235279 202989
rect 234969 194175 235279 202961
rect 234969 194147 235017 194175
rect 235045 194147 235079 194175
rect 235107 194147 235141 194175
rect 235169 194147 235203 194175
rect 235231 194147 235279 194175
rect 234969 194113 235279 194147
rect 234969 194085 235017 194113
rect 235045 194085 235079 194113
rect 235107 194085 235141 194113
rect 235169 194085 235203 194113
rect 235231 194085 235279 194113
rect 234969 194051 235279 194085
rect 234969 194023 235017 194051
rect 235045 194023 235079 194051
rect 235107 194023 235141 194051
rect 235169 194023 235203 194051
rect 235231 194023 235279 194051
rect 234969 193989 235279 194023
rect 234969 193961 235017 193989
rect 235045 193961 235079 193989
rect 235107 193961 235141 193989
rect 235169 193961 235203 193989
rect 235231 193961 235279 193989
rect 234969 185175 235279 193961
rect 234969 185147 235017 185175
rect 235045 185147 235079 185175
rect 235107 185147 235141 185175
rect 235169 185147 235203 185175
rect 235231 185147 235279 185175
rect 234969 185113 235279 185147
rect 234969 185085 235017 185113
rect 235045 185085 235079 185113
rect 235107 185085 235141 185113
rect 235169 185085 235203 185113
rect 235231 185085 235279 185113
rect 234969 185051 235279 185085
rect 234969 185023 235017 185051
rect 235045 185023 235079 185051
rect 235107 185023 235141 185051
rect 235169 185023 235203 185051
rect 235231 185023 235279 185051
rect 234969 184989 235279 185023
rect 234969 184961 235017 184989
rect 235045 184961 235079 184989
rect 235107 184961 235141 184989
rect 235169 184961 235203 184989
rect 235231 184961 235279 184989
rect 234969 176175 235279 184961
rect 234969 176147 235017 176175
rect 235045 176147 235079 176175
rect 235107 176147 235141 176175
rect 235169 176147 235203 176175
rect 235231 176147 235279 176175
rect 234969 176113 235279 176147
rect 234969 176085 235017 176113
rect 235045 176085 235079 176113
rect 235107 176085 235141 176113
rect 235169 176085 235203 176113
rect 235231 176085 235279 176113
rect 234969 176051 235279 176085
rect 234969 176023 235017 176051
rect 235045 176023 235079 176051
rect 235107 176023 235141 176051
rect 235169 176023 235203 176051
rect 235231 176023 235279 176051
rect 234969 175989 235279 176023
rect 234969 175961 235017 175989
rect 235045 175961 235079 175989
rect 235107 175961 235141 175989
rect 235169 175961 235203 175989
rect 235231 175961 235279 175989
rect 234969 167175 235279 175961
rect 248469 298606 248779 299134
rect 248469 298578 248517 298606
rect 248545 298578 248579 298606
rect 248607 298578 248641 298606
rect 248669 298578 248703 298606
rect 248731 298578 248779 298606
rect 248469 298544 248779 298578
rect 248469 298516 248517 298544
rect 248545 298516 248579 298544
rect 248607 298516 248641 298544
rect 248669 298516 248703 298544
rect 248731 298516 248779 298544
rect 248469 298482 248779 298516
rect 248469 298454 248517 298482
rect 248545 298454 248579 298482
rect 248607 298454 248641 298482
rect 248669 298454 248703 298482
rect 248731 298454 248779 298482
rect 248469 298420 248779 298454
rect 248469 298392 248517 298420
rect 248545 298392 248579 298420
rect 248607 298392 248641 298420
rect 248669 298392 248703 298420
rect 248731 298392 248779 298420
rect 248469 290175 248779 298392
rect 248469 290147 248517 290175
rect 248545 290147 248579 290175
rect 248607 290147 248641 290175
rect 248669 290147 248703 290175
rect 248731 290147 248779 290175
rect 248469 290113 248779 290147
rect 248469 290085 248517 290113
rect 248545 290085 248579 290113
rect 248607 290085 248641 290113
rect 248669 290085 248703 290113
rect 248731 290085 248779 290113
rect 248469 290051 248779 290085
rect 248469 290023 248517 290051
rect 248545 290023 248579 290051
rect 248607 290023 248641 290051
rect 248669 290023 248703 290051
rect 248731 290023 248779 290051
rect 248469 289989 248779 290023
rect 248469 289961 248517 289989
rect 248545 289961 248579 289989
rect 248607 289961 248641 289989
rect 248669 289961 248703 289989
rect 248731 289961 248779 289989
rect 248469 281175 248779 289961
rect 248469 281147 248517 281175
rect 248545 281147 248579 281175
rect 248607 281147 248641 281175
rect 248669 281147 248703 281175
rect 248731 281147 248779 281175
rect 248469 281113 248779 281147
rect 248469 281085 248517 281113
rect 248545 281085 248579 281113
rect 248607 281085 248641 281113
rect 248669 281085 248703 281113
rect 248731 281085 248779 281113
rect 248469 281051 248779 281085
rect 248469 281023 248517 281051
rect 248545 281023 248579 281051
rect 248607 281023 248641 281051
rect 248669 281023 248703 281051
rect 248731 281023 248779 281051
rect 248469 280989 248779 281023
rect 248469 280961 248517 280989
rect 248545 280961 248579 280989
rect 248607 280961 248641 280989
rect 248669 280961 248703 280989
rect 248731 280961 248779 280989
rect 248469 272175 248779 280961
rect 248469 272147 248517 272175
rect 248545 272147 248579 272175
rect 248607 272147 248641 272175
rect 248669 272147 248703 272175
rect 248731 272147 248779 272175
rect 248469 272113 248779 272147
rect 248469 272085 248517 272113
rect 248545 272085 248579 272113
rect 248607 272085 248641 272113
rect 248669 272085 248703 272113
rect 248731 272085 248779 272113
rect 248469 272051 248779 272085
rect 248469 272023 248517 272051
rect 248545 272023 248579 272051
rect 248607 272023 248641 272051
rect 248669 272023 248703 272051
rect 248731 272023 248779 272051
rect 248469 271989 248779 272023
rect 248469 271961 248517 271989
rect 248545 271961 248579 271989
rect 248607 271961 248641 271989
rect 248669 271961 248703 271989
rect 248731 271961 248779 271989
rect 248469 263175 248779 271961
rect 248469 263147 248517 263175
rect 248545 263147 248579 263175
rect 248607 263147 248641 263175
rect 248669 263147 248703 263175
rect 248731 263147 248779 263175
rect 248469 263113 248779 263147
rect 248469 263085 248517 263113
rect 248545 263085 248579 263113
rect 248607 263085 248641 263113
rect 248669 263085 248703 263113
rect 248731 263085 248779 263113
rect 248469 263051 248779 263085
rect 248469 263023 248517 263051
rect 248545 263023 248579 263051
rect 248607 263023 248641 263051
rect 248669 263023 248703 263051
rect 248731 263023 248779 263051
rect 248469 262989 248779 263023
rect 248469 262961 248517 262989
rect 248545 262961 248579 262989
rect 248607 262961 248641 262989
rect 248669 262961 248703 262989
rect 248731 262961 248779 262989
rect 248469 254175 248779 262961
rect 248469 254147 248517 254175
rect 248545 254147 248579 254175
rect 248607 254147 248641 254175
rect 248669 254147 248703 254175
rect 248731 254147 248779 254175
rect 248469 254113 248779 254147
rect 248469 254085 248517 254113
rect 248545 254085 248579 254113
rect 248607 254085 248641 254113
rect 248669 254085 248703 254113
rect 248731 254085 248779 254113
rect 248469 254051 248779 254085
rect 248469 254023 248517 254051
rect 248545 254023 248579 254051
rect 248607 254023 248641 254051
rect 248669 254023 248703 254051
rect 248731 254023 248779 254051
rect 248469 253989 248779 254023
rect 248469 253961 248517 253989
rect 248545 253961 248579 253989
rect 248607 253961 248641 253989
rect 248669 253961 248703 253989
rect 248731 253961 248779 253989
rect 248469 245175 248779 253961
rect 248469 245147 248517 245175
rect 248545 245147 248579 245175
rect 248607 245147 248641 245175
rect 248669 245147 248703 245175
rect 248731 245147 248779 245175
rect 248469 245113 248779 245147
rect 248469 245085 248517 245113
rect 248545 245085 248579 245113
rect 248607 245085 248641 245113
rect 248669 245085 248703 245113
rect 248731 245085 248779 245113
rect 248469 245051 248779 245085
rect 248469 245023 248517 245051
rect 248545 245023 248579 245051
rect 248607 245023 248641 245051
rect 248669 245023 248703 245051
rect 248731 245023 248779 245051
rect 248469 244989 248779 245023
rect 248469 244961 248517 244989
rect 248545 244961 248579 244989
rect 248607 244961 248641 244989
rect 248669 244961 248703 244989
rect 248731 244961 248779 244989
rect 248469 236175 248779 244961
rect 248469 236147 248517 236175
rect 248545 236147 248579 236175
rect 248607 236147 248641 236175
rect 248669 236147 248703 236175
rect 248731 236147 248779 236175
rect 248469 236113 248779 236147
rect 248469 236085 248517 236113
rect 248545 236085 248579 236113
rect 248607 236085 248641 236113
rect 248669 236085 248703 236113
rect 248731 236085 248779 236113
rect 248469 236051 248779 236085
rect 248469 236023 248517 236051
rect 248545 236023 248579 236051
rect 248607 236023 248641 236051
rect 248669 236023 248703 236051
rect 248731 236023 248779 236051
rect 248469 235989 248779 236023
rect 248469 235961 248517 235989
rect 248545 235961 248579 235989
rect 248607 235961 248641 235989
rect 248669 235961 248703 235989
rect 248731 235961 248779 235989
rect 248469 227175 248779 235961
rect 248469 227147 248517 227175
rect 248545 227147 248579 227175
rect 248607 227147 248641 227175
rect 248669 227147 248703 227175
rect 248731 227147 248779 227175
rect 248469 227113 248779 227147
rect 248469 227085 248517 227113
rect 248545 227085 248579 227113
rect 248607 227085 248641 227113
rect 248669 227085 248703 227113
rect 248731 227085 248779 227113
rect 248469 227051 248779 227085
rect 248469 227023 248517 227051
rect 248545 227023 248579 227051
rect 248607 227023 248641 227051
rect 248669 227023 248703 227051
rect 248731 227023 248779 227051
rect 248469 226989 248779 227023
rect 248469 226961 248517 226989
rect 248545 226961 248579 226989
rect 248607 226961 248641 226989
rect 248669 226961 248703 226989
rect 248731 226961 248779 226989
rect 248469 218175 248779 226961
rect 248469 218147 248517 218175
rect 248545 218147 248579 218175
rect 248607 218147 248641 218175
rect 248669 218147 248703 218175
rect 248731 218147 248779 218175
rect 248469 218113 248779 218147
rect 248469 218085 248517 218113
rect 248545 218085 248579 218113
rect 248607 218085 248641 218113
rect 248669 218085 248703 218113
rect 248731 218085 248779 218113
rect 248469 218051 248779 218085
rect 248469 218023 248517 218051
rect 248545 218023 248579 218051
rect 248607 218023 248641 218051
rect 248669 218023 248703 218051
rect 248731 218023 248779 218051
rect 248469 217989 248779 218023
rect 248469 217961 248517 217989
rect 248545 217961 248579 217989
rect 248607 217961 248641 217989
rect 248669 217961 248703 217989
rect 248731 217961 248779 217989
rect 248469 209175 248779 217961
rect 248469 209147 248517 209175
rect 248545 209147 248579 209175
rect 248607 209147 248641 209175
rect 248669 209147 248703 209175
rect 248731 209147 248779 209175
rect 248469 209113 248779 209147
rect 248469 209085 248517 209113
rect 248545 209085 248579 209113
rect 248607 209085 248641 209113
rect 248669 209085 248703 209113
rect 248731 209085 248779 209113
rect 248469 209051 248779 209085
rect 248469 209023 248517 209051
rect 248545 209023 248579 209051
rect 248607 209023 248641 209051
rect 248669 209023 248703 209051
rect 248731 209023 248779 209051
rect 248469 208989 248779 209023
rect 248469 208961 248517 208989
rect 248545 208961 248579 208989
rect 248607 208961 248641 208989
rect 248669 208961 248703 208989
rect 248731 208961 248779 208989
rect 248469 200175 248779 208961
rect 248469 200147 248517 200175
rect 248545 200147 248579 200175
rect 248607 200147 248641 200175
rect 248669 200147 248703 200175
rect 248731 200147 248779 200175
rect 248469 200113 248779 200147
rect 248469 200085 248517 200113
rect 248545 200085 248579 200113
rect 248607 200085 248641 200113
rect 248669 200085 248703 200113
rect 248731 200085 248779 200113
rect 248469 200051 248779 200085
rect 248469 200023 248517 200051
rect 248545 200023 248579 200051
rect 248607 200023 248641 200051
rect 248669 200023 248703 200051
rect 248731 200023 248779 200051
rect 248469 199989 248779 200023
rect 248469 199961 248517 199989
rect 248545 199961 248579 199989
rect 248607 199961 248641 199989
rect 248669 199961 248703 199989
rect 248731 199961 248779 199989
rect 248469 191175 248779 199961
rect 248469 191147 248517 191175
rect 248545 191147 248579 191175
rect 248607 191147 248641 191175
rect 248669 191147 248703 191175
rect 248731 191147 248779 191175
rect 248469 191113 248779 191147
rect 248469 191085 248517 191113
rect 248545 191085 248579 191113
rect 248607 191085 248641 191113
rect 248669 191085 248703 191113
rect 248731 191085 248779 191113
rect 248469 191051 248779 191085
rect 248469 191023 248517 191051
rect 248545 191023 248579 191051
rect 248607 191023 248641 191051
rect 248669 191023 248703 191051
rect 248731 191023 248779 191051
rect 248469 190989 248779 191023
rect 248469 190961 248517 190989
rect 248545 190961 248579 190989
rect 248607 190961 248641 190989
rect 248669 190961 248703 190989
rect 248731 190961 248779 190989
rect 248469 182175 248779 190961
rect 248469 182147 248517 182175
rect 248545 182147 248579 182175
rect 248607 182147 248641 182175
rect 248669 182147 248703 182175
rect 248731 182147 248779 182175
rect 248469 182113 248779 182147
rect 248469 182085 248517 182113
rect 248545 182085 248579 182113
rect 248607 182085 248641 182113
rect 248669 182085 248703 182113
rect 248731 182085 248779 182113
rect 248469 182051 248779 182085
rect 248469 182023 248517 182051
rect 248545 182023 248579 182051
rect 248607 182023 248641 182051
rect 248669 182023 248703 182051
rect 248731 182023 248779 182051
rect 248469 181989 248779 182023
rect 248469 181961 248517 181989
rect 248545 181961 248579 181989
rect 248607 181961 248641 181989
rect 248669 181961 248703 181989
rect 248731 181961 248779 181989
rect 238624 173175 238784 173192
rect 238624 173147 238659 173175
rect 238687 173147 238721 173175
rect 238749 173147 238784 173175
rect 238624 173113 238784 173147
rect 238624 173085 238659 173113
rect 238687 173085 238721 173113
rect 238749 173085 238784 173113
rect 238624 173051 238784 173085
rect 238624 173023 238659 173051
rect 238687 173023 238721 173051
rect 238749 173023 238784 173051
rect 238624 172989 238784 173023
rect 238624 172961 238659 172989
rect 238687 172961 238721 172989
rect 238749 172961 238784 172989
rect 238624 172944 238784 172961
rect 248469 173175 248779 181961
rect 248469 173147 248517 173175
rect 248545 173147 248579 173175
rect 248607 173147 248641 173175
rect 248669 173147 248703 173175
rect 248731 173147 248779 173175
rect 248469 173113 248779 173147
rect 248469 173085 248517 173113
rect 248545 173085 248579 173113
rect 248607 173085 248641 173113
rect 248669 173085 248703 173113
rect 248731 173085 248779 173113
rect 248469 173051 248779 173085
rect 248469 173023 248517 173051
rect 248545 173023 248579 173051
rect 248607 173023 248641 173051
rect 248669 173023 248703 173051
rect 248731 173023 248779 173051
rect 248469 172989 248779 173023
rect 248469 172961 248517 172989
rect 248545 172961 248579 172989
rect 248607 172961 248641 172989
rect 248669 172961 248703 172989
rect 248731 172961 248779 172989
rect 234969 167147 235017 167175
rect 235045 167147 235079 167175
rect 235107 167147 235141 167175
rect 235169 167147 235203 167175
rect 235231 167147 235279 167175
rect 234969 167113 235279 167147
rect 234969 167085 235017 167113
rect 235045 167085 235079 167113
rect 235107 167085 235141 167113
rect 235169 167085 235203 167113
rect 235231 167085 235279 167113
rect 234969 167051 235279 167085
rect 234969 167023 235017 167051
rect 235045 167023 235079 167051
rect 235107 167023 235141 167051
rect 235169 167023 235203 167051
rect 235231 167023 235279 167051
rect 234969 166989 235279 167023
rect 234969 166961 235017 166989
rect 235045 166961 235079 166989
rect 235107 166961 235141 166989
rect 235169 166961 235203 166989
rect 235231 166961 235279 166989
rect 234969 158175 235279 166961
rect 246304 167175 246464 167192
rect 246304 167147 246339 167175
rect 246367 167147 246401 167175
rect 246429 167147 246464 167175
rect 246304 167113 246464 167147
rect 246304 167085 246339 167113
rect 246367 167085 246401 167113
rect 246429 167085 246464 167113
rect 246304 167051 246464 167085
rect 246304 167023 246339 167051
rect 246367 167023 246401 167051
rect 246429 167023 246464 167051
rect 246304 166989 246464 167023
rect 246304 166961 246339 166989
rect 246367 166961 246401 166989
rect 246429 166961 246464 166989
rect 246304 166944 246464 166961
rect 238624 164175 238784 164192
rect 238624 164147 238659 164175
rect 238687 164147 238721 164175
rect 238749 164147 238784 164175
rect 238624 164113 238784 164147
rect 238624 164085 238659 164113
rect 238687 164085 238721 164113
rect 238749 164085 238784 164113
rect 238624 164051 238784 164085
rect 238624 164023 238659 164051
rect 238687 164023 238721 164051
rect 238749 164023 238784 164051
rect 238624 163989 238784 164023
rect 238624 163961 238659 163989
rect 238687 163961 238721 163989
rect 238749 163961 238784 163989
rect 238624 163944 238784 163961
rect 248469 164175 248779 172961
rect 248469 164147 248517 164175
rect 248545 164147 248579 164175
rect 248607 164147 248641 164175
rect 248669 164147 248703 164175
rect 248731 164147 248779 164175
rect 248469 164113 248779 164147
rect 248469 164085 248517 164113
rect 248545 164085 248579 164113
rect 248607 164085 248641 164113
rect 248669 164085 248703 164113
rect 248731 164085 248779 164113
rect 248469 164051 248779 164085
rect 248469 164023 248517 164051
rect 248545 164023 248579 164051
rect 248607 164023 248641 164051
rect 248669 164023 248703 164051
rect 248731 164023 248779 164051
rect 248469 163989 248779 164023
rect 248469 163961 248517 163989
rect 248545 163961 248579 163989
rect 248607 163961 248641 163989
rect 248669 163961 248703 163989
rect 248731 163961 248779 163989
rect 234969 158147 235017 158175
rect 235045 158147 235079 158175
rect 235107 158147 235141 158175
rect 235169 158147 235203 158175
rect 235231 158147 235279 158175
rect 234969 158113 235279 158147
rect 234969 158085 235017 158113
rect 235045 158085 235079 158113
rect 235107 158085 235141 158113
rect 235169 158085 235203 158113
rect 235231 158085 235279 158113
rect 234969 158051 235279 158085
rect 234969 158023 235017 158051
rect 235045 158023 235079 158051
rect 235107 158023 235141 158051
rect 235169 158023 235203 158051
rect 235231 158023 235279 158051
rect 234969 157989 235279 158023
rect 234969 157961 235017 157989
rect 235045 157961 235079 157989
rect 235107 157961 235141 157989
rect 235169 157961 235203 157989
rect 235231 157961 235279 157989
rect 234969 149175 235279 157961
rect 246304 158175 246464 158192
rect 246304 158147 246339 158175
rect 246367 158147 246401 158175
rect 246429 158147 246464 158175
rect 246304 158113 246464 158147
rect 246304 158085 246339 158113
rect 246367 158085 246401 158113
rect 246429 158085 246464 158113
rect 246304 158051 246464 158085
rect 246304 158023 246339 158051
rect 246367 158023 246401 158051
rect 246429 158023 246464 158051
rect 246304 157989 246464 158023
rect 246304 157961 246339 157989
rect 246367 157961 246401 157989
rect 246429 157961 246464 157989
rect 246304 157944 246464 157961
rect 238624 155175 238784 155192
rect 238624 155147 238659 155175
rect 238687 155147 238721 155175
rect 238749 155147 238784 155175
rect 238624 155113 238784 155147
rect 238624 155085 238659 155113
rect 238687 155085 238721 155113
rect 238749 155085 238784 155113
rect 238624 155051 238784 155085
rect 238624 155023 238659 155051
rect 238687 155023 238721 155051
rect 238749 155023 238784 155051
rect 238624 154989 238784 155023
rect 238624 154961 238659 154989
rect 238687 154961 238721 154989
rect 238749 154961 238784 154989
rect 238624 154944 238784 154961
rect 248469 155175 248779 163961
rect 248469 155147 248517 155175
rect 248545 155147 248579 155175
rect 248607 155147 248641 155175
rect 248669 155147 248703 155175
rect 248731 155147 248779 155175
rect 248469 155113 248779 155147
rect 248469 155085 248517 155113
rect 248545 155085 248579 155113
rect 248607 155085 248641 155113
rect 248669 155085 248703 155113
rect 248731 155085 248779 155113
rect 248469 155051 248779 155085
rect 248469 155023 248517 155051
rect 248545 155023 248579 155051
rect 248607 155023 248641 155051
rect 248669 155023 248703 155051
rect 248731 155023 248779 155051
rect 248469 154989 248779 155023
rect 248469 154961 248517 154989
rect 248545 154961 248579 154989
rect 248607 154961 248641 154989
rect 248669 154961 248703 154989
rect 248731 154961 248779 154989
rect 234969 149147 235017 149175
rect 235045 149147 235079 149175
rect 235107 149147 235141 149175
rect 235169 149147 235203 149175
rect 235231 149147 235279 149175
rect 234969 149113 235279 149147
rect 234969 149085 235017 149113
rect 235045 149085 235079 149113
rect 235107 149085 235141 149113
rect 235169 149085 235203 149113
rect 235231 149085 235279 149113
rect 234969 149051 235279 149085
rect 234969 149023 235017 149051
rect 235045 149023 235079 149051
rect 235107 149023 235141 149051
rect 235169 149023 235203 149051
rect 235231 149023 235279 149051
rect 234969 148989 235279 149023
rect 234969 148961 235017 148989
rect 235045 148961 235079 148989
rect 235107 148961 235141 148989
rect 235169 148961 235203 148989
rect 235231 148961 235279 148989
rect 234969 140175 235279 148961
rect 246304 149175 246464 149192
rect 246304 149147 246339 149175
rect 246367 149147 246401 149175
rect 246429 149147 246464 149175
rect 246304 149113 246464 149147
rect 246304 149085 246339 149113
rect 246367 149085 246401 149113
rect 246429 149085 246464 149113
rect 246304 149051 246464 149085
rect 246304 149023 246339 149051
rect 246367 149023 246401 149051
rect 246429 149023 246464 149051
rect 246304 148989 246464 149023
rect 246304 148961 246339 148989
rect 246367 148961 246401 148989
rect 246429 148961 246464 148989
rect 246304 148944 246464 148961
rect 238624 146175 238784 146192
rect 238624 146147 238659 146175
rect 238687 146147 238721 146175
rect 238749 146147 238784 146175
rect 238624 146113 238784 146147
rect 238624 146085 238659 146113
rect 238687 146085 238721 146113
rect 238749 146085 238784 146113
rect 238624 146051 238784 146085
rect 238624 146023 238659 146051
rect 238687 146023 238721 146051
rect 238749 146023 238784 146051
rect 238624 145989 238784 146023
rect 238624 145961 238659 145989
rect 238687 145961 238721 145989
rect 238749 145961 238784 145989
rect 238624 145944 238784 145961
rect 248469 146175 248779 154961
rect 248469 146147 248517 146175
rect 248545 146147 248579 146175
rect 248607 146147 248641 146175
rect 248669 146147 248703 146175
rect 248731 146147 248779 146175
rect 248469 146113 248779 146147
rect 248469 146085 248517 146113
rect 248545 146085 248579 146113
rect 248607 146085 248641 146113
rect 248669 146085 248703 146113
rect 248731 146085 248779 146113
rect 248469 146051 248779 146085
rect 248469 146023 248517 146051
rect 248545 146023 248579 146051
rect 248607 146023 248641 146051
rect 248669 146023 248703 146051
rect 248731 146023 248779 146051
rect 248469 145989 248779 146023
rect 248469 145961 248517 145989
rect 248545 145961 248579 145989
rect 248607 145961 248641 145989
rect 248669 145961 248703 145989
rect 248731 145961 248779 145989
rect 234969 140147 235017 140175
rect 235045 140147 235079 140175
rect 235107 140147 235141 140175
rect 235169 140147 235203 140175
rect 235231 140147 235279 140175
rect 234969 140113 235279 140147
rect 234969 140085 235017 140113
rect 235045 140085 235079 140113
rect 235107 140085 235141 140113
rect 235169 140085 235203 140113
rect 235231 140085 235279 140113
rect 234969 140051 235279 140085
rect 234969 140023 235017 140051
rect 235045 140023 235079 140051
rect 235107 140023 235141 140051
rect 235169 140023 235203 140051
rect 235231 140023 235279 140051
rect 234969 139989 235279 140023
rect 234969 139961 235017 139989
rect 235045 139961 235079 139989
rect 235107 139961 235141 139989
rect 235169 139961 235203 139989
rect 235231 139961 235279 139989
rect 234969 131175 235279 139961
rect 246304 140175 246464 140192
rect 246304 140147 246339 140175
rect 246367 140147 246401 140175
rect 246429 140147 246464 140175
rect 246304 140113 246464 140147
rect 246304 140085 246339 140113
rect 246367 140085 246401 140113
rect 246429 140085 246464 140113
rect 246304 140051 246464 140085
rect 246304 140023 246339 140051
rect 246367 140023 246401 140051
rect 246429 140023 246464 140051
rect 246304 139989 246464 140023
rect 246304 139961 246339 139989
rect 246367 139961 246401 139989
rect 246429 139961 246464 139989
rect 246304 139944 246464 139961
rect 238624 137175 238784 137192
rect 238624 137147 238659 137175
rect 238687 137147 238721 137175
rect 238749 137147 238784 137175
rect 238624 137113 238784 137147
rect 238624 137085 238659 137113
rect 238687 137085 238721 137113
rect 238749 137085 238784 137113
rect 238624 137051 238784 137085
rect 238624 137023 238659 137051
rect 238687 137023 238721 137051
rect 238749 137023 238784 137051
rect 238624 136989 238784 137023
rect 238624 136961 238659 136989
rect 238687 136961 238721 136989
rect 238749 136961 238784 136989
rect 238624 136944 238784 136961
rect 248469 137175 248779 145961
rect 248469 137147 248517 137175
rect 248545 137147 248579 137175
rect 248607 137147 248641 137175
rect 248669 137147 248703 137175
rect 248731 137147 248779 137175
rect 248469 137113 248779 137147
rect 248469 137085 248517 137113
rect 248545 137085 248579 137113
rect 248607 137085 248641 137113
rect 248669 137085 248703 137113
rect 248731 137085 248779 137113
rect 248469 137051 248779 137085
rect 248469 137023 248517 137051
rect 248545 137023 248579 137051
rect 248607 137023 248641 137051
rect 248669 137023 248703 137051
rect 248731 137023 248779 137051
rect 248469 136989 248779 137023
rect 248469 136961 248517 136989
rect 248545 136961 248579 136989
rect 248607 136961 248641 136989
rect 248669 136961 248703 136989
rect 248731 136961 248779 136989
rect 234969 131147 235017 131175
rect 235045 131147 235079 131175
rect 235107 131147 235141 131175
rect 235169 131147 235203 131175
rect 235231 131147 235279 131175
rect 234969 131113 235279 131147
rect 234969 131085 235017 131113
rect 235045 131085 235079 131113
rect 235107 131085 235141 131113
rect 235169 131085 235203 131113
rect 235231 131085 235279 131113
rect 234969 131051 235279 131085
rect 234969 131023 235017 131051
rect 235045 131023 235079 131051
rect 235107 131023 235141 131051
rect 235169 131023 235203 131051
rect 235231 131023 235279 131051
rect 234969 130989 235279 131023
rect 234969 130961 235017 130989
rect 235045 130961 235079 130989
rect 235107 130961 235141 130989
rect 235169 130961 235203 130989
rect 235231 130961 235279 130989
rect 234969 122175 235279 130961
rect 246304 131175 246464 131192
rect 246304 131147 246339 131175
rect 246367 131147 246401 131175
rect 246429 131147 246464 131175
rect 246304 131113 246464 131147
rect 246304 131085 246339 131113
rect 246367 131085 246401 131113
rect 246429 131085 246464 131113
rect 246304 131051 246464 131085
rect 246304 131023 246339 131051
rect 246367 131023 246401 131051
rect 246429 131023 246464 131051
rect 246304 130989 246464 131023
rect 246304 130961 246339 130989
rect 246367 130961 246401 130989
rect 246429 130961 246464 130989
rect 246304 130944 246464 130961
rect 238624 128175 238784 128192
rect 238624 128147 238659 128175
rect 238687 128147 238721 128175
rect 238749 128147 238784 128175
rect 238624 128113 238784 128147
rect 238624 128085 238659 128113
rect 238687 128085 238721 128113
rect 238749 128085 238784 128113
rect 238624 128051 238784 128085
rect 238624 128023 238659 128051
rect 238687 128023 238721 128051
rect 238749 128023 238784 128051
rect 238624 127989 238784 128023
rect 238624 127961 238659 127989
rect 238687 127961 238721 127989
rect 238749 127961 238784 127989
rect 238624 127944 238784 127961
rect 248469 128175 248779 136961
rect 248469 128147 248517 128175
rect 248545 128147 248579 128175
rect 248607 128147 248641 128175
rect 248669 128147 248703 128175
rect 248731 128147 248779 128175
rect 248469 128113 248779 128147
rect 248469 128085 248517 128113
rect 248545 128085 248579 128113
rect 248607 128085 248641 128113
rect 248669 128085 248703 128113
rect 248731 128085 248779 128113
rect 248469 128051 248779 128085
rect 248469 128023 248517 128051
rect 248545 128023 248579 128051
rect 248607 128023 248641 128051
rect 248669 128023 248703 128051
rect 248731 128023 248779 128051
rect 248469 127989 248779 128023
rect 248469 127961 248517 127989
rect 248545 127961 248579 127989
rect 248607 127961 248641 127989
rect 248669 127961 248703 127989
rect 248731 127961 248779 127989
rect 234969 122147 235017 122175
rect 235045 122147 235079 122175
rect 235107 122147 235141 122175
rect 235169 122147 235203 122175
rect 235231 122147 235279 122175
rect 234969 122113 235279 122147
rect 234969 122085 235017 122113
rect 235045 122085 235079 122113
rect 235107 122085 235141 122113
rect 235169 122085 235203 122113
rect 235231 122085 235279 122113
rect 234969 122051 235279 122085
rect 234969 122023 235017 122051
rect 235045 122023 235079 122051
rect 235107 122023 235141 122051
rect 235169 122023 235203 122051
rect 235231 122023 235279 122051
rect 234969 121989 235279 122023
rect 234969 121961 235017 121989
rect 235045 121961 235079 121989
rect 235107 121961 235141 121989
rect 235169 121961 235203 121989
rect 235231 121961 235279 121989
rect 234969 113175 235279 121961
rect 246304 122175 246464 122192
rect 246304 122147 246339 122175
rect 246367 122147 246401 122175
rect 246429 122147 246464 122175
rect 246304 122113 246464 122147
rect 246304 122085 246339 122113
rect 246367 122085 246401 122113
rect 246429 122085 246464 122113
rect 246304 122051 246464 122085
rect 246304 122023 246339 122051
rect 246367 122023 246401 122051
rect 246429 122023 246464 122051
rect 246304 121989 246464 122023
rect 246304 121961 246339 121989
rect 246367 121961 246401 121989
rect 246429 121961 246464 121989
rect 246304 121944 246464 121961
rect 238624 119175 238784 119192
rect 238624 119147 238659 119175
rect 238687 119147 238721 119175
rect 238749 119147 238784 119175
rect 238624 119113 238784 119147
rect 238624 119085 238659 119113
rect 238687 119085 238721 119113
rect 238749 119085 238784 119113
rect 238624 119051 238784 119085
rect 238624 119023 238659 119051
rect 238687 119023 238721 119051
rect 238749 119023 238784 119051
rect 238624 118989 238784 119023
rect 238624 118961 238659 118989
rect 238687 118961 238721 118989
rect 238749 118961 238784 118989
rect 238624 118944 238784 118961
rect 248469 119175 248779 127961
rect 248469 119147 248517 119175
rect 248545 119147 248579 119175
rect 248607 119147 248641 119175
rect 248669 119147 248703 119175
rect 248731 119147 248779 119175
rect 248469 119113 248779 119147
rect 248469 119085 248517 119113
rect 248545 119085 248579 119113
rect 248607 119085 248641 119113
rect 248669 119085 248703 119113
rect 248731 119085 248779 119113
rect 248469 119051 248779 119085
rect 248469 119023 248517 119051
rect 248545 119023 248579 119051
rect 248607 119023 248641 119051
rect 248669 119023 248703 119051
rect 248731 119023 248779 119051
rect 248469 118989 248779 119023
rect 248469 118961 248517 118989
rect 248545 118961 248579 118989
rect 248607 118961 248641 118989
rect 248669 118961 248703 118989
rect 248731 118961 248779 118989
rect 234969 113147 235017 113175
rect 235045 113147 235079 113175
rect 235107 113147 235141 113175
rect 235169 113147 235203 113175
rect 235231 113147 235279 113175
rect 234969 113113 235279 113147
rect 234969 113085 235017 113113
rect 235045 113085 235079 113113
rect 235107 113085 235141 113113
rect 235169 113085 235203 113113
rect 235231 113085 235279 113113
rect 234969 113051 235279 113085
rect 234969 113023 235017 113051
rect 235045 113023 235079 113051
rect 235107 113023 235141 113051
rect 235169 113023 235203 113051
rect 235231 113023 235279 113051
rect 234969 112989 235279 113023
rect 234969 112961 235017 112989
rect 235045 112961 235079 112989
rect 235107 112961 235141 112989
rect 235169 112961 235203 112989
rect 235231 112961 235279 112989
rect 234969 104175 235279 112961
rect 246304 113175 246464 113192
rect 246304 113147 246339 113175
rect 246367 113147 246401 113175
rect 246429 113147 246464 113175
rect 246304 113113 246464 113147
rect 246304 113085 246339 113113
rect 246367 113085 246401 113113
rect 246429 113085 246464 113113
rect 246304 113051 246464 113085
rect 246304 113023 246339 113051
rect 246367 113023 246401 113051
rect 246429 113023 246464 113051
rect 246304 112989 246464 113023
rect 246304 112961 246339 112989
rect 246367 112961 246401 112989
rect 246429 112961 246464 112989
rect 246304 112944 246464 112961
rect 238624 110175 238784 110192
rect 238624 110147 238659 110175
rect 238687 110147 238721 110175
rect 238749 110147 238784 110175
rect 238624 110113 238784 110147
rect 238624 110085 238659 110113
rect 238687 110085 238721 110113
rect 238749 110085 238784 110113
rect 238624 110051 238784 110085
rect 238624 110023 238659 110051
rect 238687 110023 238721 110051
rect 238749 110023 238784 110051
rect 238624 109989 238784 110023
rect 238624 109961 238659 109989
rect 238687 109961 238721 109989
rect 238749 109961 238784 109989
rect 238624 109944 238784 109961
rect 248469 110175 248779 118961
rect 248469 110147 248517 110175
rect 248545 110147 248579 110175
rect 248607 110147 248641 110175
rect 248669 110147 248703 110175
rect 248731 110147 248779 110175
rect 248469 110113 248779 110147
rect 248469 110085 248517 110113
rect 248545 110085 248579 110113
rect 248607 110085 248641 110113
rect 248669 110085 248703 110113
rect 248731 110085 248779 110113
rect 248469 110051 248779 110085
rect 248469 110023 248517 110051
rect 248545 110023 248579 110051
rect 248607 110023 248641 110051
rect 248669 110023 248703 110051
rect 248731 110023 248779 110051
rect 248469 109989 248779 110023
rect 248469 109961 248517 109989
rect 248545 109961 248579 109989
rect 248607 109961 248641 109989
rect 248669 109961 248703 109989
rect 248731 109961 248779 109989
rect 234969 104147 235017 104175
rect 235045 104147 235079 104175
rect 235107 104147 235141 104175
rect 235169 104147 235203 104175
rect 235231 104147 235279 104175
rect 234969 104113 235279 104147
rect 234969 104085 235017 104113
rect 235045 104085 235079 104113
rect 235107 104085 235141 104113
rect 235169 104085 235203 104113
rect 235231 104085 235279 104113
rect 234969 104051 235279 104085
rect 234969 104023 235017 104051
rect 235045 104023 235079 104051
rect 235107 104023 235141 104051
rect 235169 104023 235203 104051
rect 235231 104023 235279 104051
rect 234969 103989 235279 104023
rect 234969 103961 235017 103989
rect 235045 103961 235079 103989
rect 235107 103961 235141 103989
rect 235169 103961 235203 103989
rect 235231 103961 235279 103989
rect 234969 95175 235279 103961
rect 246304 104175 246464 104192
rect 246304 104147 246339 104175
rect 246367 104147 246401 104175
rect 246429 104147 246464 104175
rect 246304 104113 246464 104147
rect 246304 104085 246339 104113
rect 246367 104085 246401 104113
rect 246429 104085 246464 104113
rect 246304 104051 246464 104085
rect 246304 104023 246339 104051
rect 246367 104023 246401 104051
rect 246429 104023 246464 104051
rect 246304 103989 246464 104023
rect 246304 103961 246339 103989
rect 246367 103961 246401 103989
rect 246429 103961 246464 103989
rect 246304 103944 246464 103961
rect 238624 101175 238784 101192
rect 238624 101147 238659 101175
rect 238687 101147 238721 101175
rect 238749 101147 238784 101175
rect 238624 101113 238784 101147
rect 238624 101085 238659 101113
rect 238687 101085 238721 101113
rect 238749 101085 238784 101113
rect 238624 101051 238784 101085
rect 238624 101023 238659 101051
rect 238687 101023 238721 101051
rect 238749 101023 238784 101051
rect 238624 100989 238784 101023
rect 238624 100961 238659 100989
rect 238687 100961 238721 100989
rect 238749 100961 238784 100989
rect 238624 100944 238784 100961
rect 248469 101175 248779 109961
rect 248469 101147 248517 101175
rect 248545 101147 248579 101175
rect 248607 101147 248641 101175
rect 248669 101147 248703 101175
rect 248731 101147 248779 101175
rect 248469 101113 248779 101147
rect 248469 101085 248517 101113
rect 248545 101085 248579 101113
rect 248607 101085 248641 101113
rect 248669 101085 248703 101113
rect 248731 101085 248779 101113
rect 248469 101051 248779 101085
rect 248469 101023 248517 101051
rect 248545 101023 248579 101051
rect 248607 101023 248641 101051
rect 248669 101023 248703 101051
rect 248731 101023 248779 101051
rect 248469 100989 248779 101023
rect 248469 100961 248517 100989
rect 248545 100961 248579 100989
rect 248607 100961 248641 100989
rect 248669 100961 248703 100989
rect 248731 100961 248779 100989
rect 234969 95147 235017 95175
rect 235045 95147 235079 95175
rect 235107 95147 235141 95175
rect 235169 95147 235203 95175
rect 235231 95147 235279 95175
rect 234969 95113 235279 95147
rect 234969 95085 235017 95113
rect 235045 95085 235079 95113
rect 235107 95085 235141 95113
rect 235169 95085 235203 95113
rect 235231 95085 235279 95113
rect 234969 95051 235279 95085
rect 234969 95023 235017 95051
rect 235045 95023 235079 95051
rect 235107 95023 235141 95051
rect 235169 95023 235203 95051
rect 235231 95023 235279 95051
rect 234969 94989 235279 95023
rect 234969 94961 235017 94989
rect 235045 94961 235079 94989
rect 235107 94961 235141 94989
rect 235169 94961 235203 94989
rect 235231 94961 235279 94989
rect 234969 86175 235279 94961
rect 246304 95175 246464 95192
rect 246304 95147 246339 95175
rect 246367 95147 246401 95175
rect 246429 95147 246464 95175
rect 246304 95113 246464 95147
rect 246304 95085 246339 95113
rect 246367 95085 246401 95113
rect 246429 95085 246464 95113
rect 246304 95051 246464 95085
rect 246304 95023 246339 95051
rect 246367 95023 246401 95051
rect 246429 95023 246464 95051
rect 246304 94989 246464 95023
rect 246304 94961 246339 94989
rect 246367 94961 246401 94989
rect 246429 94961 246464 94989
rect 246304 94944 246464 94961
rect 238624 92175 238784 92192
rect 238624 92147 238659 92175
rect 238687 92147 238721 92175
rect 238749 92147 238784 92175
rect 238624 92113 238784 92147
rect 238624 92085 238659 92113
rect 238687 92085 238721 92113
rect 238749 92085 238784 92113
rect 238624 92051 238784 92085
rect 238624 92023 238659 92051
rect 238687 92023 238721 92051
rect 238749 92023 238784 92051
rect 238624 91989 238784 92023
rect 238624 91961 238659 91989
rect 238687 91961 238721 91989
rect 238749 91961 238784 91989
rect 238624 91944 238784 91961
rect 248469 92175 248779 100961
rect 248469 92147 248517 92175
rect 248545 92147 248579 92175
rect 248607 92147 248641 92175
rect 248669 92147 248703 92175
rect 248731 92147 248779 92175
rect 248469 92113 248779 92147
rect 248469 92085 248517 92113
rect 248545 92085 248579 92113
rect 248607 92085 248641 92113
rect 248669 92085 248703 92113
rect 248731 92085 248779 92113
rect 248469 92051 248779 92085
rect 248469 92023 248517 92051
rect 248545 92023 248579 92051
rect 248607 92023 248641 92051
rect 248669 92023 248703 92051
rect 248731 92023 248779 92051
rect 248469 91989 248779 92023
rect 248469 91961 248517 91989
rect 248545 91961 248579 91989
rect 248607 91961 248641 91989
rect 248669 91961 248703 91989
rect 248731 91961 248779 91989
rect 234969 86147 235017 86175
rect 235045 86147 235079 86175
rect 235107 86147 235141 86175
rect 235169 86147 235203 86175
rect 235231 86147 235279 86175
rect 234969 86113 235279 86147
rect 234969 86085 235017 86113
rect 235045 86085 235079 86113
rect 235107 86085 235141 86113
rect 235169 86085 235203 86113
rect 235231 86085 235279 86113
rect 234969 86051 235279 86085
rect 234969 86023 235017 86051
rect 235045 86023 235079 86051
rect 235107 86023 235141 86051
rect 235169 86023 235203 86051
rect 235231 86023 235279 86051
rect 234969 85989 235279 86023
rect 234969 85961 235017 85989
rect 235045 85961 235079 85989
rect 235107 85961 235141 85989
rect 235169 85961 235203 85989
rect 235231 85961 235279 85989
rect 234969 77175 235279 85961
rect 246304 86175 246464 86192
rect 246304 86147 246339 86175
rect 246367 86147 246401 86175
rect 246429 86147 246464 86175
rect 246304 86113 246464 86147
rect 246304 86085 246339 86113
rect 246367 86085 246401 86113
rect 246429 86085 246464 86113
rect 246304 86051 246464 86085
rect 246304 86023 246339 86051
rect 246367 86023 246401 86051
rect 246429 86023 246464 86051
rect 246304 85989 246464 86023
rect 246304 85961 246339 85989
rect 246367 85961 246401 85989
rect 246429 85961 246464 85989
rect 246304 85944 246464 85961
rect 238624 83175 238784 83192
rect 238624 83147 238659 83175
rect 238687 83147 238721 83175
rect 238749 83147 238784 83175
rect 238624 83113 238784 83147
rect 238624 83085 238659 83113
rect 238687 83085 238721 83113
rect 238749 83085 238784 83113
rect 238624 83051 238784 83085
rect 238624 83023 238659 83051
rect 238687 83023 238721 83051
rect 238749 83023 238784 83051
rect 238624 82989 238784 83023
rect 238624 82961 238659 82989
rect 238687 82961 238721 82989
rect 238749 82961 238784 82989
rect 238624 82944 238784 82961
rect 248469 83175 248779 91961
rect 248469 83147 248517 83175
rect 248545 83147 248579 83175
rect 248607 83147 248641 83175
rect 248669 83147 248703 83175
rect 248731 83147 248779 83175
rect 248469 83113 248779 83147
rect 248469 83085 248517 83113
rect 248545 83085 248579 83113
rect 248607 83085 248641 83113
rect 248669 83085 248703 83113
rect 248731 83085 248779 83113
rect 248469 83051 248779 83085
rect 248469 83023 248517 83051
rect 248545 83023 248579 83051
rect 248607 83023 248641 83051
rect 248669 83023 248703 83051
rect 248731 83023 248779 83051
rect 248469 82989 248779 83023
rect 248469 82961 248517 82989
rect 248545 82961 248579 82989
rect 248607 82961 248641 82989
rect 248669 82961 248703 82989
rect 248731 82961 248779 82989
rect 234969 77147 235017 77175
rect 235045 77147 235079 77175
rect 235107 77147 235141 77175
rect 235169 77147 235203 77175
rect 235231 77147 235279 77175
rect 234969 77113 235279 77147
rect 234969 77085 235017 77113
rect 235045 77085 235079 77113
rect 235107 77085 235141 77113
rect 235169 77085 235203 77113
rect 235231 77085 235279 77113
rect 234969 77051 235279 77085
rect 234969 77023 235017 77051
rect 235045 77023 235079 77051
rect 235107 77023 235141 77051
rect 235169 77023 235203 77051
rect 235231 77023 235279 77051
rect 234969 76989 235279 77023
rect 234969 76961 235017 76989
rect 235045 76961 235079 76989
rect 235107 76961 235141 76989
rect 235169 76961 235203 76989
rect 235231 76961 235279 76989
rect 234969 68175 235279 76961
rect 246304 77175 246464 77192
rect 246304 77147 246339 77175
rect 246367 77147 246401 77175
rect 246429 77147 246464 77175
rect 246304 77113 246464 77147
rect 246304 77085 246339 77113
rect 246367 77085 246401 77113
rect 246429 77085 246464 77113
rect 246304 77051 246464 77085
rect 246304 77023 246339 77051
rect 246367 77023 246401 77051
rect 246429 77023 246464 77051
rect 246304 76989 246464 77023
rect 246304 76961 246339 76989
rect 246367 76961 246401 76989
rect 246429 76961 246464 76989
rect 246304 76944 246464 76961
rect 238624 74175 238784 74192
rect 238624 74147 238659 74175
rect 238687 74147 238721 74175
rect 238749 74147 238784 74175
rect 238624 74113 238784 74147
rect 238624 74085 238659 74113
rect 238687 74085 238721 74113
rect 238749 74085 238784 74113
rect 238624 74051 238784 74085
rect 238624 74023 238659 74051
rect 238687 74023 238721 74051
rect 238749 74023 238784 74051
rect 238624 73989 238784 74023
rect 238624 73961 238659 73989
rect 238687 73961 238721 73989
rect 238749 73961 238784 73989
rect 238624 73944 238784 73961
rect 248469 74175 248779 82961
rect 248469 74147 248517 74175
rect 248545 74147 248579 74175
rect 248607 74147 248641 74175
rect 248669 74147 248703 74175
rect 248731 74147 248779 74175
rect 248469 74113 248779 74147
rect 248469 74085 248517 74113
rect 248545 74085 248579 74113
rect 248607 74085 248641 74113
rect 248669 74085 248703 74113
rect 248731 74085 248779 74113
rect 248469 74051 248779 74085
rect 248469 74023 248517 74051
rect 248545 74023 248579 74051
rect 248607 74023 248641 74051
rect 248669 74023 248703 74051
rect 248731 74023 248779 74051
rect 248469 73989 248779 74023
rect 248469 73961 248517 73989
rect 248545 73961 248579 73989
rect 248607 73961 248641 73989
rect 248669 73961 248703 73989
rect 248731 73961 248779 73989
rect 234969 68147 235017 68175
rect 235045 68147 235079 68175
rect 235107 68147 235141 68175
rect 235169 68147 235203 68175
rect 235231 68147 235279 68175
rect 234969 68113 235279 68147
rect 234969 68085 235017 68113
rect 235045 68085 235079 68113
rect 235107 68085 235141 68113
rect 235169 68085 235203 68113
rect 235231 68085 235279 68113
rect 234969 68051 235279 68085
rect 234969 68023 235017 68051
rect 235045 68023 235079 68051
rect 235107 68023 235141 68051
rect 235169 68023 235203 68051
rect 235231 68023 235279 68051
rect 234969 67989 235279 68023
rect 234969 67961 235017 67989
rect 235045 67961 235079 67989
rect 235107 67961 235141 67989
rect 235169 67961 235203 67989
rect 235231 67961 235279 67989
rect 234969 59175 235279 67961
rect 246304 68175 246464 68192
rect 246304 68147 246339 68175
rect 246367 68147 246401 68175
rect 246429 68147 246464 68175
rect 246304 68113 246464 68147
rect 246304 68085 246339 68113
rect 246367 68085 246401 68113
rect 246429 68085 246464 68113
rect 246304 68051 246464 68085
rect 246304 68023 246339 68051
rect 246367 68023 246401 68051
rect 246429 68023 246464 68051
rect 246304 67989 246464 68023
rect 246304 67961 246339 67989
rect 246367 67961 246401 67989
rect 246429 67961 246464 67989
rect 246304 67944 246464 67961
rect 238624 65175 238784 65192
rect 238624 65147 238659 65175
rect 238687 65147 238721 65175
rect 238749 65147 238784 65175
rect 238624 65113 238784 65147
rect 238624 65085 238659 65113
rect 238687 65085 238721 65113
rect 238749 65085 238784 65113
rect 238624 65051 238784 65085
rect 238624 65023 238659 65051
rect 238687 65023 238721 65051
rect 238749 65023 238784 65051
rect 238624 64989 238784 65023
rect 238624 64961 238659 64989
rect 238687 64961 238721 64989
rect 238749 64961 238784 64989
rect 238624 64944 238784 64961
rect 248469 65175 248779 73961
rect 248469 65147 248517 65175
rect 248545 65147 248579 65175
rect 248607 65147 248641 65175
rect 248669 65147 248703 65175
rect 248731 65147 248779 65175
rect 248469 65113 248779 65147
rect 248469 65085 248517 65113
rect 248545 65085 248579 65113
rect 248607 65085 248641 65113
rect 248669 65085 248703 65113
rect 248731 65085 248779 65113
rect 248469 65051 248779 65085
rect 248469 65023 248517 65051
rect 248545 65023 248579 65051
rect 248607 65023 248641 65051
rect 248669 65023 248703 65051
rect 248731 65023 248779 65051
rect 248469 64989 248779 65023
rect 248469 64961 248517 64989
rect 248545 64961 248579 64989
rect 248607 64961 248641 64989
rect 248669 64961 248703 64989
rect 248731 64961 248779 64989
rect 234969 59147 235017 59175
rect 235045 59147 235079 59175
rect 235107 59147 235141 59175
rect 235169 59147 235203 59175
rect 235231 59147 235279 59175
rect 234969 59113 235279 59147
rect 234969 59085 235017 59113
rect 235045 59085 235079 59113
rect 235107 59085 235141 59113
rect 235169 59085 235203 59113
rect 235231 59085 235279 59113
rect 234969 59051 235279 59085
rect 234969 59023 235017 59051
rect 235045 59023 235079 59051
rect 235107 59023 235141 59051
rect 235169 59023 235203 59051
rect 235231 59023 235279 59051
rect 234969 58989 235279 59023
rect 234969 58961 235017 58989
rect 235045 58961 235079 58989
rect 235107 58961 235141 58989
rect 235169 58961 235203 58989
rect 235231 58961 235279 58989
rect 234969 50175 235279 58961
rect 246304 59175 246464 59192
rect 246304 59147 246339 59175
rect 246367 59147 246401 59175
rect 246429 59147 246464 59175
rect 246304 59113 246464 59147
rect 246304 59085 246339 59113
rect 246367 59085 246401 59113
rect 246429 59085 246464 59113
rect 246304 59051 246464 59085
rect 246304 59023 246339 59051
rect 246367 59023 246401 59051
rect 246429 59023 246464 59051
rect 246304 58989 246464 59023
rect 246304 58961 246339 58989
rect 246367 58961 246401 58989
rect 246429 58961 246464 58989
rect 246304 58944 246464 58961
rect 238624 56175 238784 56192
rect 238624 56147 238659 56175
rect 238687 56147 238721 56175
rect 238749 56147 238784 56175
rect 238624 56113 238784 56147
rect 238624 56085 238659 56113
rect 238687 56085 238721 56113
rect 238749 56085 238784 56113
rect 238624 56051 238784 56085
rect 238624 56023 238659 56051
rect 238687 56023 238721 56051
rect 238749 56023 238784 56051
rect 238624 55989 238784 56023
rect 238624 55961 238659 55989
rect 238687 55961 238721 55989
rect 238749 55961 238784 55989
rect 238624 55944 238784 55961
rect 248469 56175 248779 64961
rect 248469 56147 248517 56175
rect 248545 56147 248579 56175
rect 248607 56147 248641 56175
rect 248669 56147 248703 56175
rect 248731 56147 248779 56175
rect 248469 56113 248779 56147
rect 248469 56085 248517 56113
rect 248545 56085 248579 56113
rect 248607 56085 248641 56113
rect 248669 56085 248703 56113
rect 248731 56085 248779 56113
rect 248469 56051 248779 56085
rect 248469 56023 248517 56051
rect 248545 56023 248579 56051
rect 248607 56023 248641 56051
rect 248669 56023 248703 56051
rect 248731 56023 248779 56051
rect 248469 55989 248779 56023
rect 248469 55961 248517 55989
rect 248545 55961 248579 55989
rect 248607 55961 248641 55989
rect 248669 55961 248703 55989
rect 248731 55961 248779 55989
rect 234969 50147 235017 50175
rect 235045 50147 235079 50175
rect 235107 50147 235141 50175
rect 235169 50147 235203 50175
rect 235231 50147 235279 50175
rect 234969 50113 235279 50147
rect 234969 50085 235017 50113
rect 235045 50085 235079 50113
rect 235107 50085 235141 50113
rect 235169 50085 235203 50113
rect 235231 50085 235279 50113
rect 234969 50051 235279 50085
rect 234969 50023 235017 50051
rect 235045 50023 235079 50051
rect 235107 50023 235141 50051
rect 235169 50023 235203 50051
rect 235231 50023 235279 50051
rect 234969 49989 235279 50023
rect 234969 49961 235017 49989
rect 235045 49961 235079 49989
rect 235107 49961 235141 49989
rect 235169 49961 235203 49989
rect 235231 49961 235279 49989
rect 234969 41175 235279 49961
rect 246304 50175 246464 50192
rect 246304 50147 246339 50175
rect 246367 50147 246401 50175
rect 246429 50147 246464 50175
rect 246304 50113 246464 50147
rect 246304 50085 246339 50113
rect 246367 50085 246401 50113
rect 246429 50085 246464 50113
rect 246304 50051 246464 50085
rect 246304 50023 246339 50051
rect 246367 50023 246401 50051
rect 246429 50023 246464 50051
rect 246304 49989 246464 50023
rect 246304 49961 246339 49989
rect 246367 49961 246401 49989
rect 246429 49961 246464 49989
rect 246304 49944 246464 49961
rect 238624 47175 238784 47192
rect 238624 47147 238659 47175
rect 238687 47147 238721 47175
rect 238749 47147 238784 47175
rect 238624 47113 238784 47147
rect 238624 47085 238659 47113
rect 238687 47085 238721 47113
rect 238749 47085 238784 47113
rect 238624 47051 238784 47085
rect 238624 47023 238659 47051
rect 238687 47023 238721 47051
rect 238749 47023 238784 47051
rect 238624 46989 238784 47023
rect 238624 46961 238659 46989
rect 238687 46961 238721 46989
rect 238749 46961 238784 46989
rect 238624 46944 238784 46961
rect 248469 47175 248779 55961
rect 248469 47147 248517 47175
rect 248545 47147 248579 47175
rect 248607 47147 248641 47175
rect 248669 47147 248703 47175
rect 248731 47147 248779 47175
rect 248469 47113 248779 47147
rect 248469 47085 248517 47113
rect 248545 47085 248579 47113
rect 248607 47085 248641 47113
rect 248669 47085 248703 47113
rect 248731 47085 248779 47113
rect 248469 47051 248779 47085
rect 248469 47023 248517 47051
rect 248545 47023 248579 47051
rect 248607 47023 248641 47051
rect 248669 47023 248703 47051
rect 248731 47023 248779 47051
rect 248469 46989 248779 47023
rect 248469 46961 248517 46989
rect 248545 46961 248579 46989
rect 248607 46961 248641 46989
rect 248669 46961 248703 46989
rect 248731 46961 248779 46989
rect 234969 41147 235017 41175
rect 235045 41147 235079 41175
rect 235107 41147 235141 41175
rect 235169 41147 235203 41175
rect 235231 41147 235279 41175
rect 234969 41113 235279 41147
rect 234969 41085 235017 41113
rect 235045 41085 235079 41113
rect 235107 41085 235141 41113
rect 235169 41085 235203 41113
rect 235231 41085 235279 41113
rect 234969 41051 235279 41085
rect 234969 41023 235017 41051
rect 235045 41023 235079 41051
rect 235107 41023 235141 41051
rect 235169 41023 235203 41051
rect 235231 41023 235279 41051
rect 234969 40989 235279 41023
rect 234969 40961 235017 40989
rect 235045 40961 235079 40989
rect 235107 40961 235141 40989
rect 235169 40961 235203 40989
rect 235231 40961 235279 40989
rect 234969 32175 235279 40961
rect 246304 41175 246464 41192
rect 246304 41147 246339 41175
rect 246367 41147 246401 41175
rect 246429 41147 246464 41175
rect 246304 41113 246464 41147
rect 246304 41085 246339 41113
rect 246367 41085 246401 41113
rect 246429 41085 246464 41113
rect 246304 41051 246464 41085
rect 246304 41023 246339 41051
rect 246367 41023 246401 41051
rect 246429 41023 246464 41051
rect 246304 40989 246464 41023
rect 246304 40961 246339 40989
rect 246367 40961 246401 40989
rect 246429 40961 246464 40989
rect 246304 40944 246464 40961
rect 238624 38175 238784 38192
rect 238624 38147 238659 38175
rect 238687 38147 238721 38175
rect 238749 38147 238784 38175
rect 238624 38113 238784 38147
rect 238624 38085 238659 38113
rect 238687 38085 238721 38113
rect 238749 38085 238784 38113
rect 238624 38051 238784 38085
rect 238624 38023 238659 38051
rect 238687 38023 238721 38051
rect 238749 38023 238784 38051
rect 238624 37989 238784 38023
rect 238624 37961 238659 37989
rect 238687 37961 238721 37989
rect 238749 37961 238784 37989
rect 238624 37944 238784 37961
rect 248469 38175 248779 46961
rect 248469 38147 248517 38175
rect 248545 38147 248579 38175
rect 248607 38147 248641 38175
rect 248669 38147 248703 38175
rect 248731 38147 248779 38175
rect 248469 38113 248779 38147
rect 248469 38085 248517 38113
rect 248545 38085 248579 38113
rect 248607 38085 248641 38113
rect 248669 38085 248703 38113
rect 248731 38085 248779 38113
rect 248469 38051 248779 38085
rect 248469 38023 248517 38051
rect 248545 38023 248579 38051
rect 248607 38023 248641 38051
rect 248669 38023 248703 38051
rect 248731 38023 248779 38051
rect 248469 37989 248779 38023
rect 248469 37961 248517 37989
rect 248545 37961 248579 37989
rect 248607 37961 248641 37989
rect 248669 37961 248703 37989
rect 248731 37961 248779 37989
rect 234969 32147 235017 32175
rect 235045 32147 235079 32175
rect 235107 32147 235141 32175
rect 235169 32147 235203 32175
rect 235231 32147 235279 32175
rect 234969 32113 235279 32147
rect 234969 32085 235017 32113
rect 235045 32085 235079 32113
rect 235107 32085 235141 32113
rect 235169 32085 235203 32113
rect 235231 32085 235279 32113
rect 234969 32051 235279 32085
rect 234969 32023 235017 32051
rect 235045 32023 235079 32051
rect 235107 32023 235141 32051
rect 235169 32023 235203 32051
rect 235231 32023 235279 32051
rect 234969 31989 235279 32023
rect 234969 31961 235017 31989
rect 235045 31961 235079 31989
rect 235107 31961 235141 31989
rect 235169 31961 235203 31989
rect 235231 31961 235279 31989
rect 234969 23175 235279 31961
rect 246304 32175 246464 32192
rect 246304 32147 246339 32175
rect 246367 32147 246401 32175
rect 246429 32147 246464 32175
rect 246304 32113 246464 32147
rect 246304 32085 246339 32113
rect 246367 32085 246401 32113
rect 246429 32085 246464 32113
rect 246304 32051 246464 32085
rect 246304 32023 246339 32051
rect 246367 32023 246401 32051
rect 246429 32023 246464 32051
rect 246304 31989 246464 32023
rect 246304 31961 246339 31989
rect 246367 31961 246401 31989
rect 246429 31961 246464 31989
rect 246304 31944 246464 31961
rect 238624 29175 238784 29192
rect 238624 29147 238659 29175
rect 238687 29147 238721 29175
rect 238749 29147 238784 29175
rect 238624 29113 238784 29147
rect 238624 29085 238659 29113
rect 238687 29085 238721 29113
rect 238749 29085 238784 29113
rect 238624 29051 238784 29085
rect 238624 29023 238659 29051
rect 238687 29023 238721 29051
rect 238749 29023 238784 29051
rect 238624 28989 238784 29023
rect 238624 28961 238659 28989
rect 238687 28961 238721 28989
rect 238749 28961 238784 28989
rect 238624 28944 238784 28961
rect 248469 29175 248779 37961
rect 248469 29147 248517 29175
rect 248545 29147 248579 29175
rect 248607 29147 248641 29175
rect 248669 29147 248703 29175
rect 248731 29147 248779 29175
rect 248469 29113 248779 29147
rect 248469 29085 248517 29113
rect 248545 29085 248579 29113
rect 248607 29085 248641 29113
rect 248669 29085 248703 29113
rect 248731 29085 248779 29113
rect 248469 29051 248779 29085
rect 248469 29023 248517 29051
rect 248545 29023 248579 29051
rect 248607 29023 248641 29051
rect 248669 29023 248703 29051
rect 248731 29023 248779 29051
rect 248469 28989 248779 29023
rect 248469 28961 248517 28989
rect 248545 28961 248579 28989
rect 248607 28961 248641 28989
rect 248669 28961 248703 28989
rect 248731 28961 248779 28989
rect 234969 23147 235017 23175
rect 235045 23147 235079 23175
rect 235107 23147 235141 23175
rect 235169 23147 235203 23175
rect 235231 23147 235279 23175
rect 234969 23113 235279 23147
rect 234969 23085 235017 23113
rect 235045 23085 235079 23113
rect 235107 23085 235141 23113
rect 235169 23085 235203 23113
rect 235231 23085 235279 23113
rect 234969 23051 235279 23085
rect 234969 23023 235017 23051
rect 235045 23023 235079 23051
rect 235107 23023 235141 23051
rect 235169 23023 235203 23051
rect 235231 23023 235279 23051
rect 234969 22989 235279 23023
rect 234969 22961 235017 22989
rect 235045 22961 235079 22989
rect 235107 22961 235141 22989
rect 235169 22961 235203 22989
rect 235231 22961 235279 22989
rect 234969 14175 235279 22961
rect 246304 23175 246464 23192
rect 246304 23147 246339 23175
rect 246367 23147 246401 23175
rect 246429 23147 246464 23175
rect 246304 23113 246464 23147
rect 246304 23085 246339 23113
rect 246367 23085 246401 23113
rect 246429 23085 246464 23113
rect 246304 23051 246464 23085
rect 246304 23023 246339 23051
rect 246367 23023 246401 23051
rect 246429 23023 246464 23051
rect 246304 22989 246464 23023
rect 246304 22961 246339 22989
rect 246367 22961 246401 22989
rect 246429 22961 246464 22989
rect 246304 22944 246464 22961
rect 238624 20175 238784 20192
rect 238624 20147 238659 20175
rect 238687 20147 238721 20175
rect 238749 20147 238784 20175
rect 238624 20113 238784 20147
rect 238624 20085 238659 20113
rect 238687 20085 238721 20113
rect 238749 20085 238784 20113
rect 238624 20051 238784 20085
rect 238624 20023 238659 20051
rect 238687 20023 238721 20051
rect 238749 20023 238784 20051
rect 238624 19989 238784 20023
rect 238624 19961 238659 19989
rect 238687 19961 238721 19989
rect 238749 19961 238784 19989
rect 238624 19944 238784 19961
rect 248469 20175 248779 28961
rect 248469 20147 248517 20175
rect 248545 20147 248579 20175
rect 248607 20147 248641 20175
rect 248669 20147 248703 20175
rect 248731 20147 248779 20175
rect 248469 20113 248779 20147
rect 248469 20085 248517 20113
rect 248545 20085 248579 20113
rect 248607 20085 248641 20113
rect 248669 20085 248703 20113
rect 248731 20085 248779 20113
rect 248469 20051 248779 20085
rect 248469 20023 248517 20051
rect 248545 20023 248579 20051
rect 248607 20023 248641 20051
rect 248669 20023 248703 20051
rect 248731 20023 248779 20051
rect 248469 19989 248779 20023
rect 248469 19961 248517 19989
rect 248545 19961 248579 19989
rect 248607 19961 248641 19989
rect 248669 19961 248703 19989
rect 248731 19961 248779 19989
rect 234969 14147 235017 14175
rect 235045 14147 235079 14175
rect 235107 14147 235141 14175
rect 235169 14147 235203 14175
rect 235231 14147 235279 14175
rect 234969 14113 235279 14147
rect 234969 14085 235017 14113
rect 235045 14085 235079 14113
rect 235107 14085 235141 14113
rect 235169 14085 235203 14113
rect 235231 14085 235279 14113
rect 234969 14051 235279 14085
rect 234969 14023 235017 14051
rect 235045 14023 235079 14051
rect 235107 14023 235141 14051
rect 235169 14023 235203 14051
rect 235231 14023 235279 14051
rect 234969 13989 235279 14023
rect 234969 13961 235017 13989
rect 235045 13961 235079 13989
rect 235107 13961 235141 13989
rect 235169 13961 235203 13989
rect 235231 13961 235279 13989
rect 234969 5175 235279 13961
rect 246304 14175 246464 14192
rect 246304 14147 246339 14175
rect 246367 14147 246401 14175
rect 246429 14147 246464 14175
rect 246304 14113 246464 14147
rect 246304 14085 246339 14113
rect 246367 14085 246401 14113
rect 246429 14085 246464 14113
rect 246304 14051 246464 14085
rect 246304 14023 246339 14051
rect 246367 14023 246401 14051
rect 246429 14023 246464 14051
rect 246304 13989 246464 14023
rect 246304 13961 246339 13989
rect 246367 13961 246401 13989
rect 246429 13961 246464 13989
rect 246304 13944 246464 13961
rect 238624 11175 238784 11192
rect 238624 11147 238659 11175
rect 238687 11147 238721 11175
rect 238749 11147 238784 11175
rect 238624 11113 238784 11147
rect 238624 11085 238659 11113
rect 238687 11085 238721 11113
rect 238749 11085 238784 11113
rect 238624 11051 238784 11085
rect 238624 11023 238659 11051
rect 238687 11023 238721 11051
rect 238749 11023 238784 11051
rect 238624 10989 238784 11023
rect 238624 10961 238659 10989
rect 238687 10961 238721 10989
rect 238749 10961 238784 10989
rect 238624 10944 238784 10961
rect 248469 11175 248779 19961
rect 248469 11147 248517 11175
rect 248545 11147 248579 11175
rect 248607 11147 248641 11175
rect 248669 11147 248703 11175
rect 248731 11147 248779 11175
rect 248469 11113 248779 11147
rect 248469 11085 248517 11113
rect 248545 11085 248579 11113
rect 248607 11085 248641 11113
rect 248669 11085 248703 11113
rect 248731 11085 248779 11113
rect 248469 11051 248779 11085
rect 248469 11023 248517 11051
rect 248545 11023 248579 11051
rect 248607 11023 248641 11051
rect 248669 11023 248703 11051
rect 248731 11023 248779 11051
rect 248469 10989 248779 11023
rect 248469 10961 248517 10989
rect 248545 10961 248579 10989
rect 248607 10961 248641 10989
rect 248669 10961 248703 10989
rect 248731 10961 248779 10989
rect 234969 5147 235017 5175
rect 235045 5147 235079 5175
rect 235107 5147 235141 5175
rect 235169 5147 235203 5175
rect 235231 5147 235279 5175
rect 234969 5113 235279 5147
rect 234969 5085 235017 5113
rect 235045 5085 235079 5113
rect 235107 5085 235141 5113
rect 235169 5085 235203 5113
rect 235231 5085 235279 5113
rect 234969 5051 235279 5085
rect 234969 5023 235017 5051
rect 235045 5023 235079 5051
rect 235107 5023 235141 5051
rect 235169 5023 235203 5051
rect 235231 5023 235279 5051
rect 234969 4989 235279 5023
rect 234969 4961 235017 4989
rect 235045 4961 235079 4989
rect 235107 4961 235141 4989
rect 235169 4961 235203 4989
rect 235231 4961 235279 4989
rect 234969 -560 235279 4961
rect 246304 5175 246464 5192
rect 246304 5147 246339 5175
rect 246367 5147 246401 5175
rect 246429 5147 246464 5175
rect 246304 5113 246464 5147
rect 246304 5085 246339 5113
rect 246367 5085 246401 5113
rect 246429 5085 246464 5113
rect 246304 5051 246464 5085
rect 246304 5023 246339 5051
rect 246367 5023 246401 5051
rect 246429 5023 246464 5051
rect 246304 4989 246464 5023
rect 246304 4961 246339 4989
rect 246367 4961 246401 4989
rect 246429 4961 246464 4989
rect 246304 4944 246464 4961
rect 234969 -588 235017 -560
rect 235045 -588 235079 -560
rect 235107 -588 235141 -560
rect 235169 -588 235203 -560
rect 235231 -588 235279 -560
rect 234969 -622 235279 -588
rect 234969 -650 235017 -622
rect 235045 -650 235079 -622
rect 235107 -650 235141 -622
rect 235169 -650 235203 -622
rect 235231 -650 235279 -622
rect 234969 -684 235279 -650
rect 234969 -712 235017 -684
rect 235045 -712 235079 -684
rect 235107 -712 235141 -684
rect 235169 -712 235203 -684
rect 235231 -712 235279 -684
rect 234969 -746 235279 -712
rect 234969 -774 235017 -746
rect 235045 -774 235079 -746
rect 235107 -774 235141 -746
rect 235169 -774 235203 -746
rect 235231 -774 235279 -746
rect 234969 -822 235279 -774
rect 248469 2175 248779 10961
rect 248469 2147 248517 2175
rect 248545 2147 248579 2175
rect 248607 2147 248641 2175
rect 248669 2147 248703 2175
rect 248731 2147 248779 2175
rect 248469 2113 248779 2147
rect 248469 2085 248517 2113
rect 248545 2085 248579 2113
rect 248607 2085 248641 2113
rect 248669 2085 248703 2113
rect 248731 2085 248779 2113
rect 248469 2051 248779 2085
rect 248469 2023 248517 2051
rect 248545 2023 248579 2051
rect 248607 2023 248641 2051
rect 248669 2023 248703 2051
rect 248731 2023 248779 2051
rect 248469 1989 248779 2023
rect 248469 1961 248517 1989
rect 248545 1961 248579 1989
rect 248607 1961 248641 1989
rect 248669 1961 248703 1989
rect 248731 1961 248779 1989
rect 248469 -80 248779 1961
rect 248469 -108 248517 -80
rect 248545 -108 248579 -80
rect 248607 -108 248641 -80
rect 248669 -108 248703 -80
rect 248731 -108 248779 -80
rect 248469 -142 248779 -108
rect 248469 -170 248517 -142
rect 248545 -170 248579 -142
rect 248607 -170 248641 -142
rect 248669 -170 248703 -142
rect 248731 -170 248779 -142
rect 248469 -204 248779 -170
rect 248469 -232 248517 -204
rect 248545 -232 248579 -204
rect 248607 -232 248641 -204
rect 248669 -232 248703 -204
rect 248731 -232 248779 -204
rect 248469 -266 248779 -232
rect 248469 -294 248517 -266
rect 248545 -294 248579 -266
rect 248607 -294 248641 -266
rect 248669 -294 248703 -266
rect 248731 -294 248779 -266
rect 248469 -822 248779 -294
rect 250329 299086 250639 299134
rect 250329 299058 250377 299086
rect 250405 299058 250439 299086
rect 250467 299058 250501 299086
rect 250529 299058 250563 299086
rect 250591 299058 250639 299086
rect 250329 299024 250639 299058
rect 250329 298996 250377 299024
rect 250405 298996 250439 299024
rect 250467 298996 250501 299024
rect 250529 298996 250563 299024
rect 250591 298996 250639 299024
rect 250329 298962 250639 298996
rect 250329 298934 250377 298962
rect 250405 298934 250439 298962
rect 250467 298934 250501 298962
rect 250529 298934 250563 298962
rect 250591 298934 250639 298962
rect 250329 298900 250639 298934
rect 250329 298872 250377 298900
rect 250405 298872 250439 298900
rect 250467 298872 250501 298900
rect 250529 298872 250563 298900
rect 250591 298872 250639 298900
rect 250329 293175 250639 298872
rect 250329 293147 250377 293175
rect 250405 293147 250439 293175
rect 250467 293147 250501 293175
rect 250529 293147 250563 293175
rect 250591 293147 250639 293175
rect 250329 293113 250639 293147
rect 250329 293085 250377 293113
rect 250405 293085 250439 293113
rect 250467 293085 250501 293113
rect 250529 293085 250563 293113
rect 250591 293085 250639 293113
rect 250329 293051 250639 293085
rect 250329 293023 250377 293051
rect 250405 293023 250439 293051
rect 250467 293023 250501 293051
rect 250529 293023 250563 293051
rect 250591 293023 250639 293051
rect 250329 292989 250639 293023
rect 250329 292961 250377 292989
rect 250405 292961 250439 292989
rect 250467 292961 250501 292989
rect 250529 292961 250563 292989
rect 250591 292961 250639 292989
rect 250329 284175 250639 292961
rect 250329 284147 250377 284175
rect 250405 284147 250439 284175
rect 250467 284147 250501 284175
rect 250529 284147 250563 284175
rect 250591 284147 250639 284175
rect 250329 284113 250639 284147
rect 250329 284085 250377 284113
rect 250405 284085 250439 284113
rect 250467 284085 250501 284113
rect 250529 284085 250563 284113
rect 250591 284085 250639 284113
rect 250329 284051 250639 284085
rect 250329 284023 250377 284051
rect 250405 284023 250439 284051
rect 250467 284023 250501 284051
rect 250529 284023 250563 284051
rect 250591 284023 250639 284051
rect 250329 283989 250639 284023
rect 250329 283961 250377 283989
rect 250405 283961 250439 283989
rect 250467 283961 250501 283989
rect 250529 283961 250563 283989
rect 250591 283961 250639 283989
rect 250329 275175 250639 283961
rect 250329 275147 250377 275175
rect 250405 275147 250439 275175
rect 250467 275147 250501 275175
rect 250529 275147 250563 275175
rect 250591 275147 250639 275175
rect 250329 275113 250639 275147
rect 250329 275085 250377 275113
rect 250405 275085 250439 275113
rect 250467 275085 250501 275113
rect 250529 275085 250563 275113
rect 250591 275085 250639 275113
rect 250329 275051 250639 275085
rect 250329 275023 250377 275051
rect 250405 275023 250439 275051
rect 250467 275023 250501 275051
rect 250529 275023 250563 275051
rect 250591 275023 250639 275051
rect 250329 274989 250639 275023
rect 250329 274961 250377 274989
rect 250405 274961 250439 274989
rect 250467 274961 250501 274989
rect 250529 274961 250563 274989
rect 250591 274961 250639 274989
rect 250329 266175 250639 274961
rect 250329 266147 250377 266175
rect 250405 266147 250439 266175
rect 250467 266147 250501 266175
rect 250529 266147 250563 266175
rect 250591 266147 250639 266175
rect 250329 266113 250639 266147
rect 250329 266085 250377 266113
rect 250405 266085 250439 266113
rect 250467 266085 250501 266113
rect 250529 266085 250563 266113
rect 250591 266085 250639 266113
rect 250329 266051 250639 266085
rect 250329 266023 250377 266051
rect 250405 266023 250439 266051
rect 250467 266023 250501 266051
rect 250529 266023 250563 266051
rect 250591 266023 250639 266051
rect 250329 265989 250639 266023
rect 250329 265961 250377 265989
rect 250405 265961 250439 265989
rect 250467 265961 250501 265989
rect 250529 265961 250563 265989
rect 250591 265961 250639 265989
rect 250329 257175 250639 265961
rect 250329 257147 250377 257175
rect 250405 257147 250439 257175
rect 250467 257147 250501 257175
rect 250529 257147 250563 257175
rect 250591 257147 250639 257175
rect 250329 257113 250639 257147
rect 250329 257085 250377 257113
rect 250405 257085 250439 257113
rect 250467 257085 250501 257113
rect 250529 257085 250563 257113
rect 250591 257085 250639 257113
rect 250329 257051 250639 257085
rect 250329 257023 250377 257051
rect 250405 257023 250439 257051
rect 250467 257023 250501 257051
rect 250529 257023 250563 257051
rect 250591 257023 250639 257051
rect 250329 256989 250639 257023
rect 250329 256961 250377 256989
rect 250405 256961 250439 256989
rect 250467 256961 250501 256989
rect 250529 256961 250563 256989
rect 250591 256961 250639 256989
rect 250329 248175 250639 256961
rect 250329 248147 250377 248175
rect 250405 248147 250439 248175
rect 250467 248147 250501 248175
rect 250529 248147 250563 248175
rect 250591 248147 250639 248175
rect 250329 248113 250639 248147
rect 250329 248085 250377 248113
rect 250405 248085 250439 248113
rect 250467 248085 250501 248113
rect 250529 248085 250563 248113
rect 250591 248085 250639 248113
rect 250329 248051 250639 248085
rect 250329 248023 250377 248051
rect 250405 248023 250439 248051
rect 250467 248023 250501 248051
rect 250529 248023 250563 248051
rect 250591 248023 250639 248051
rect 250329 247989 250639 248023
rect 250329 247961 250377 247989
rect 250405 247961 250439 247989
rect 250467 247961 250501 247989
rect 250529 247961 250563 247989
rect 250591 247961 250639 247989
rect 250329 239175 250639 247961
rect 250329 239147 250377 239175
rect 250405 239147 250439 239175
rect 250467 239147 250501 239175
rect 250529 239147 250563 239175
rect 250591 239147 250639 239175
rect 250329 239113 250639 239147
rect 250329 239085 250377 239113
rect 250405 239085 250439 239113
rect 250467 239085 250501 239113
rect 250529 239085 250563 239113
rect 250591 239085 250639 239113
rect 250329 239051 250639 239085
rect 250329 239023 250377 239051
rect 250405 239023 250439 239051
rect 250467 239023 250501 239051
rect 250529 239023 250563 239051
rect 250591 239023 250639 239051
rect 250329 238989 250639 239023
rect 250329 238961 250377 238989
rect 250405 238961 250439 238989
rect 250467 238961 250501 238989
rect 250529 238961 250563 238989
rect 250591 238961 250639 238989
rect 250329 230175 250639 238961
rect 250329 230147 250377 230175
rect 250405 230147 250439 230175
rect 250467 230147 250501 230175
rect 250529 230147 250563 230175
rect 250591 230147 250639 230175
rect 250329 230113 250639 230147
rect 250329 230085 250377 230113
rect 250405 230085 250439 230113
rect 250467 230085 250501 230113
rect 250529 230085 250563 230113
rect 250591 230085 250639 230113
rect 250329 230051 250639 230085
rect 250329 230023 250377 230051
rect 250405 230023 250439 230051
rect 250467 230023 250501 230051
rect 250529 230023 250563 230051
rect 250591 230023 250639 230051
rect 250329 229989 250639 230023
rect 250329 229961 250377 229989
rect 250405 229961 250439 229989
rect 250467 229961 250501 229989
rect 250529 229961 250563 229989
rect 250591 229961 250639 229989
rect 250329 221175 250639 229961
rect 250329 221147 250377 221175
rect 250405 221147 250439 221175
rect 250467 221147 250501 221175
rect 250529 221147 250563 221175
rect 250591 221147 250639 221175
rect 250329 221113 250639 221147
rect 250329 221085 250377 221113
rect 250405 221085 250439 221113
rect 250467 221085 250501 221113
rect 250529 221085 250563 221113
rect 250591 221085 250639 221113
rect 250329 221051 250639 221085
rect 250329 221023 250377 221051
rect 250405 221023 250439 221051
rect 250467 221023 250501 221051
rect 250529 221023 250563 221051
rect 250591 221023 250639 221051
rect 250329 220989 250639 221023
rect 250329 220961 250377 220989
rect 250405 220961 250439 220989
rect 250467 220961 250501 220989
rect 250529 220961 250563 220989
rect 250591 220961 250639 220989
rect 250329 212175 250639 220961
rect 250329 212147 250377 212175
rect 250405 212147 250439 212175
rect 250467 212147 250501 212175
rect 250529 212147 250563 212175
rect 250591 212147 250639 212175
rect 250329 212113 250639 212147
rect 250329 212085 250377 212113
rect 250405 212085 250439 212113
rect 250467 212085 250501 212113
rect 250529 212085 250563 212113
rect 250591 212085 250639 212113
rect 250329 212051 250639 212085
rect 250329 212023 250377 212051
rect 250405 212023 250439 212051
rect 250467 212023 250501 212051
rect 250529 212023 250563 212051
rect 250591 212023 250639 212051
rect 250329 211989 250639 212023
rect 250329 211961 250377 211989
rect 250405 211961 250439 211989
rect 250467 211961 250501 211989
rect 250529 211961 250563 211989
rect 250591 211961 250639 211989
rect 250329 203175 250639 211961
rect 250329 203147 250377 203175
rect 250405 203147 250439 203175
rect 250467 203147 250501 203175
rect 250529 203147 250563 203175
rect 250591 203147 250639 203175
rect 250329 203113 250639 203147
rect 250329 203085 250377 203113
rect 250405 203085 250439 203113
rect 250467 203085 250501 203113
rect 250529 203085 250563 203113
rect 250591 203085 250639 203113
rect 250329 203051 250639 203085
rect 250329 203023 250377 203051
rect 250405 203023 250439 203051
rect 250467 203023 250501 203051
rect 250529 203023 250563 203051
rect 250591 203023 250639 203051
rect 250329 202989 250639 203023
rect 250329 202961 250377 202989
rect 250405 202961 250439 202989
rect 250467 202961 250501 202989
rect 250529 202961 250563 202989
rect 250591 202961 250639 202989
rect 250329 194175 250639 202961
rect 250329 194147 250377 194175
rect 250405 194147 250439 194175
rect 250467 194147 250501 194175
rect 250529 194147 250563 194175
rect 250591 194147 250639 194175
rect 250329 194113 250639 194147
rect 250329 194085 250377 194113
rect 250405 194085 250439 194113
rect 250467 194085 250501 194113
rect 250529 194085 250563 194113
rect 250591 194085 250639 194113
rect 250329 194051 250639 194085
rect 250329 194023 250377 194051
rect 250405 194023 250439 194051
rect 250467 194023 250501 194051
rect 250529 194023 250563 194051
rect 250591 194023 250639 194051
rect 250329 193989 250639 194023
rect 250329 193961 250377 193989
rect 250405 193961 250439 193989
rect 250467 193961 250501 193989
rect 250529 193961 250563 193989
rect 250591 193961 250639 193989
rect 250329 185175 250639 193961
rect 250329 185147 250377 185175
rect 250405 185147 250439 185175
rect 250467 185147 250501 185175
rect 250529 185147 250563 185175
rect 250591 185147 250639 185175
rect 250329 185113 250639 185147
rect 250329 185085 250377 185113
rect 250405 185085 250439 185113
rect 250467 185085 250501 185113
rect 250529 185085 250563 185113
rect 250591 185085 250639 185113
rect 250329 185051 250639 185085
rect 250329 185023 250377 185051
rect 250405 185023 250439 185051
rect 250467 185023 250501 185051
rect 250529 185023 250563 185051
rect 250591 185023 250639 185051
rect 250329 184989 250639 185023
rect 250329 184961 250377 184989
rect 250405 184961 250439 184989
rect 250467 184961 250501 184989
rect 250529 184961 250563 184989
rect 250591 184961 250639 184989
rect 250329 176175 250639 184961
rect 250329 176147 250377 176175
rect 250405 176147 250439 176175
rect 250467 176147 250501 176175
rect 250529 176147 250563 176175
rect 250591 176147 250639 176175
rect 250329 176113 250639 176147
rect 250329 176085 250377 176113
rect 250405 176085 250439 176113
rect 250467 176085 250501 176113
rect 250529 176085 250563 176113
rect 250591 176085 250639 176113
rect 250329 176051 250639 176085
rect 250329 176023 250377 176051
rect 250405 176023 250439 176051
rect 250467 176023 250501 176051
rect 250529 176023 250563 176051
rect 250591 176023 250639 176051
rect 250329 175989 250639 176023
rect 250329 175961 250377 175989
rect 250405 175961 250439 175989
rect 250467 175961 250501 175989
rect 250529 175961 250563 175989
rect 250591 175961 250639 175989
rect 250329 167175 250639 175961
rect 263829 298606 264139 299134
rect 263829 298578 263877 298606
rect 263905 298578 263939 298606
rect 263967 298578 264001 298606
rect 264029 298578 264063 298606
rect 264091 298578 264139 298606
rect 263829 298544 264139 298578
rect 263829 298516 263877 298544
rect 263905 298516 263939 298544
rect 263967 298516 264001 298544
rect 264029 298516 264063 298544
rect 264091 298516 264139 298544
rect 263829 298482 264139 298516
rect 263829 298454 263877 298482
rect 263905 298454 263939 298482
rect 263967 298454 264001 298482
rect 264029 298454 264063 298482
rect 264091 298454 264139 298482
rect 263829 298420 264139 298454
rect 263829 298392 263877 298420
rect 263905 298392 263939 298420
rect 263967 298392 264001 298420
rect 264029 298392 264063 298420
rect 264091 298392 264139 298420
rect 263829 290175 264139 298392
rect 263829 290147 263877 290175
rect 263905 290147 263939 290175
rect 263967 290147 264001 290175
rect 264029 290147 264063 290175
rect 264091 290147 264139 290175
rect 263829 290113 264139 290147
rect 263829 290085 263877 290113
rect 263905 290085 263939 290113
rect 263967 290085 264001 290113
rect 264029 290085 264063 290113
rect 264091 290085 264139 290113
rect 263829 290051 264139 290085
rect 263829 290023 263877 290051
rect 263905 290023 263939 290051
rect 263967 290023 264001 290051
rect 264029 290023 264063 290051
rect 264091 290023 264139 290051
rect 263829 289989 264139 290023
rect 263829 289961 263877 289989
rect 263905 289961 263939 289989
rect 263967 289961 264001 289989
rect 264029 289961 264063 289989
rect 264091 289961 264139 289989
rect 263829 281175 264139 289961
rect 263829 281147 263877 281175
rect 263905 281147 263939 281175
rect 263967 281147 264001 281175
rect 264029 281147 264063 281175
rect 264091 281147 264139 281175
rect 263829 281113 264139 281147
rect 263829 281085 263877 281113
rect 263905 281085 263939 281113
rect 263967 281085 264001 281113
rect 264029 281085 264063 281113
rect 264091 281085 264139 281113
rect 263829 281051 264139 281085
rect 263829 281023 263877 281051
rect 263905 281023 263939 281051
rect 263967 281023 264001 281051
rect 264029 281023 264063 281051
rect 264091 281023 264139 281051
rect 263829 280989 264139 281023
rect 263829 280961 263877 280989
rect 263905 280961 263939 280989
rect 263967 280961 264001 280989
rect 264029 280961 264063 280989
rect 264091 280961 264139 280989
rect 263829 272175 264139 280961
rect 263829 272147 263877 272175
rect 263905 272147 263939 272175
rect 263967 272147 264001 272175
rect 264029 272147 264063 272175
rect 264091 272147 264139 272175
rect 263829 272113 264139 272147
rect 263829 272085 263877 272113
rect 263905 272085 263939 272113
rect 263967 272085 264001 272113
rect 264029 272085 264063 272113
rect 264091 272085 264139 272113
rect 263829 272051 264139 272085
rect 263829 272023 263877 272051
rect 263905 272023 263939 272051
rect 263967 272023 264001 272051
rect 264029 272023 264063 272051
rect 264091 272023 264139 272051
rect 263829 271989 264139 272023
rect 263829 271961 263877 271989
rect 263905 271961 263939 271989
rect 263967 271961 264001 271989
rect 264029 271961 264063 271989
rect 264091 271961 264139 271989
rect 263829 263175 264139 271961
rect 263829 263147 263877 263175
rect 263905 263147 263939 263175
rect 263967 263147 264001 263175
rect 264029 263147 264063 263175
rect 264091 263147 264139 263175
rect 263829 263113 264139 263147
rect 263829 263085 263877 263113
rect 263905 263085 263939 263113
rect 263967 263085 264001 263113
rect 264029 263085 264063 263113
rect 264091 263085 264139 263113
rect 263829 263051 264139 263085
rect 263829 263023 263877 263051
rect 263905 263023 263939 263051
rect 263967 263023 264001 263051
rect 264029 263023 264063 263051
rect 264091 263023 264139 263051
rect 263829 262989 264139 263023
rect 263829 262961 263877 262989
rect 263905 262961 263939 262989
rect 263967 262961 264001 262989
rect 264029 262961 264063 262989
rect 264091 262961 264139 262989
rect 263829 254175 264139 262961
rect 263829 254147 263877 254175
rect 263905 254147 263939 254175
rect 263967 254147 264001 254175
rect 264029 254147 264063 254175
rect 264091 254147 264139 254175
rect 263829 254113 264139 254147
rect 263829 254085 263877 254113
rect 263905 254085 263939 254113
rect 263967 254085 264001 254113
rect 264029 254085 264063 254113
rect 264091 254085 264139 254113
rect 263829 254051 264139 254085
rect 263829 254023 263877 254051
rect 263905 254023 263939 254051
rect 263967 254023 264001 254051
rect 264029 254023 264063 254051
rect 264091 254023 264139 254051
rect 263829 253989 264139 254023
rect 263829 253961 263877 253989
rect 263905 253961 263939 253989
rect 263967 253961 264001 253989
rect 264029 253961 264063 253989
rect 264091 253961 264139 253989
rect 263829 245175 264139 253961
rect 263829 245147 263877 245175
rect 263905 245147 263939 245175
rect 263967 245147 264001 245175
rect 264029 245147 264063 245175
rect 264091 245147 264139 245175
rect 263829 245113 264139 245147
rect 263829 245085 263877 245113
rect 263905 245085 263939 245113
rect 263967 245085 264001 245113
rect 264029 245085 264063 245113
rect 264091 245085 264139 245113
rect 263829 245051 264139 245085
rect 263829 245023 263877 245051
rect 263905 245023 263939 245051
rect 263967 245023 264001 245051
rect 264029 245023 264063 245051
rect 264091 245023 264139 245051
rect 263829 244989 264139 245023
rect 263829 244961 263877 244989
rect 263905 244961 263939 244989
rect 263967 244961 264001 244989
rect 264029 244961 264063 244989
rect 264091 244961 264139 244989
rect 263829 236175 264139 244961
rect 263829 236147 263877 236175
rect 263905 236147 263939 236175
rect 263967 236147 264001 236175
rect 264029 236147 264063 236175
rect 264091 236147 264139 236175
rect 263829 236113 264139 236147
rect 263829 236085 263877 236113
rect 263905 236085 263939 236113
rect 263967 236085 264001 236113
rect 264029 236085 264063 236113
rect 264091 236085 264139 236113
rect 263829 236051 264139 236085
rect 263829 236023 263877 236051
rect 263905 236023 263939 236051
rect 263967 236023 264001 236051
rect 264029 236023 264063 236051
rect 264091 236023 264139 236051
rect 263829 235989 264139 236023
rect 263829 235961 263877 235989
rect 263905 235961 263939 235989
rect 263967 235961 264001 235989
rect 264029 235961 264063 235989
rect 264091 235961 264139 235989
rect 263829 227175 264139 235961
rect 263829 227147 263877 227175
rect 263905 227147 263939 227175
rect 263967 227147 264001 227175
rect 264029 227147 264063 227175
rect 264091 227147 264139 227175
rect 263829 227113 264139 227147
rect 263829 227085 263877 227113
rect 263905 227085 263939 227113
rect 263967 227085 264001 227113
rect 264029 227085 264063 227113
rect 264091 227085 264139 227113
rect 263829 227051 264139 227085
rect 263829 227023 263877 227051
rect 263905 227023 263939 227051
rect 263967 227023 264001 227051
rect 264029 227023 264063 227051
rect 264091 227023 264139 227051
rect 263829 226989 264139 227023
rect 263829 226961 263877 226989
rect 263905 226961 263939 226989
rect 263967 226961 264001 226989
rect 264029 226961 264063 226989
rect 264091 226961 264139 226989
rect 263829 218175 264139 226961
rect 263829 218147 263877 218175
rect 263905 218147 263939 218175
rect 263967 218147 264001 218175
rect 264029 218147 264063 218175
rect 264091 218147 264139 218175
rect 263829 218113 264139 218147
rect 263829 218085 263877 218113
rect 263905 218085 263939 218113
rect 263967 218085 264001 218113
rect 264029 218085 264063 218113
rect 264091 218085 264139 218113
rect 263829 218051 264139 218085
rect 263829 218023 263877 218051
rect 263905 218023 263939 218051
rect 263967 218023 264001 218051
rect 264029 218023 264063 218051
rect 264091 218023 264139 218051
rect 263829 217989 264139 218023
rect 263829 217961 263877 217989
rect 263905 217961 263939 217989
rect 263967 217961 264001 217989
rect 264029 217961 264063 217989
rect 264091 217961 264139 217989
rect 263829 209175 264139 217961
rect 263829 209147 263877 209175
rect 263905 209147 263939 209175
rect 263967 209147 264001 209175
rect 264029 209147 264063 209175
rect 264091 209147 264139 209175
rect 263829 209113 264139 209147
rect 263829 209085 263877 209113
rect 263905 209085 263939 209113
rect 263967 209085 264001 209113
rect 264029 209085 264063 209113
rect 264091 209085 264139 209113
rect 263829 209051 264139 209085
rect 263829 209023 263877 209051
rect 263905 209023 263939 209051
rect 263967 209023 264001 209051
rect 264029 209023 264063 209051
rect 264091 209023 264139 209051
rect 263829 208989 264139 209023
rect 263829 208961 263877 208989
rect 263905 208961 263939 208989
rect 263967 208961 264001 208989
rect 264029 208961 264063 208989
rect 264091 208961 264139 208989
rect 263829 200175 264139 208961
rect 263829 200147 263877 200175
rect 263905 200147 263939 200175
rect 263967 200147 264001 200175
rect 264029 200147 264063 200175
rect 264091 200147 264139 200175
rect 263829 200113 264139 200147
rect 263829 200085 263877 200113
rect 263905 200085 263939 200113
rect 263967 200085 264001 200113
rect 264029 200085 264063 200113
rect 264091 200085 264139 200113
rect 263829 200051 264139 200085
rect 263829 200023 263877 200051
rect 263905 200023 263939 200051
rect 263967 200023 264001 200051
rect 264029 200023 264063 200051
rect 264091 200023 264139 200051
rect 263829 199989 264139 200023
rect 263829 199961 263877 199989
rect 263905 199961 263939 199989
rect 263967 199961 264001 199989
rect 264029 199961 264063 199989
rect 264091 199961 264139 199989
rect 263829 191175 264139 199961
rect 263829 191147 263877 191175
rect 263905 191147 263939 191175
rect 263967 191147 264001 191175
rect 264029 191147 264063 191175
rect 264091 191147 264139 191175
rect 263829 191113 264139 191147
rect 263829 191085 263877 191113
rect 263905 191085 263939 191113
rect 263967 191085 264001 191113
rect 264029 191085 264063 191113
rect 264091 191085 264139 191113
rect 263829 191051 264139 191085
rect 263829 191023 263877 191051
rect 263905 191023 263939 191051
rect 263967 191023 264001 191051
rect 264029 191023 264063 191051
rect 264091 191023 264139 191051
rect 263829 190989 264139 191023
rect 263829 190961 263877 190989
rect 263905 190961 263939 190989
rect 263967 190961 264001 190989
rect 264029 190961 264063 190989
rect 264091 190961 264139 190989
rect 263829 182175 264139 190961
rect 263829 182147 263877 182175
rect 263905 182147 263939 182175
rect 263967 182147 264001 182175
rect 264029 182147 264063 182175
rect 264091 182147 264139 182175
rect 263829 182113 264139 182147
rect 263829 182085 263877 182113
rect 263905 182085 263939 182113
rect 263967 182085 264001 182113
rect 264029 182085 264063 182113
rect 264091 182085 264139 182113
rect 263829 182051 264139 182085
rect 263829 182023 263877 182051
rect 263905 182023 263939 182051
rect 263967 182023 264001 182051
rect 264029 182023 264063 182051
rect 264091 182023 264139 182051
rect 263829 181989 264139 182023
rect 263829 181961 263877 181989
rect 263905 181961 263939 181989
rect 263967 181961 264001 181989
rect 264029 181961 264063 181989
rect 264091 181961 264139 181989
rect 253984 173175 254144 173192
rect 253984 173147 254019 173175
rect 254047 173147 254081 173175
rect 254109 173147 254144 173175
rect 253984 173113 254144 173147
rect 253984 173085 254019 173113
rect 254047 173085 254081 173113
rect 254109 173085 254144 173113
rect 253984 173051 254144 173085
rect 253984 173023 254019 173051
rect 254047 173023 254081 173051
rect 254109 173023 254144 173051
rect 253984 172989 254144 173023
rect 253984 172961 254019 172989
rect 254047 172961 254081 172989
rect 254109 172961 254144 172989
rect 253984 172944 254144 172961
rect 263829 173175 264139 181961
rect 263829 173147 263877 173175
rect 263905 173147 263939 173175
rect 263967 173147 264001 173175
rect 264029 173147 264063 173175
rect 264091 173147 264139 173175
rect 263829 173113 264139 173147
rect 263829 173085 263877 173113
rect 263905 173085 263939 173113
rect 263967 173085 264001 173113
rect 264029 173085 264063 173113
rect 264091 173085 264139 173113
rect 263829 173051 264139 173085
rect 263829 173023 263877 173051
rect 263905 173023 263939 173051
rect 263967 173023 264001 173051
rect 264029 173023 264063 173051
rect 264091 173023 264139 173051
rect 263829 172989 264139 173023
rect 263829 172961 263877 172989
rect 263905 172961 263939 172989
rect 263967 172961 264001 172989
rect 264029 172961 264063 172989
rect 264091 172961 264139 172989
rect 250329 167147 250377 167175
rect 250405 167147 250439 167175
rect 250467 167147 250501 167175
rect 250529 167147 250563 167175
rect 250591 167147 250639 167175
rect 250329 167113 250639 167147
rect 250329 167085 250377 167113
rect 250405 167085 250439 167113
rect 250467 167085 250501 167113
rect 250529 167085 250563 167113
rect 250591 167085 250639 167113
rect 250329 167051 250639 167085
rect 250329 167023 250377 167051
rect 250405 167023 250439 167051
rect 250467 167023 250501 167051
rect 250529 167023 250563 167051
rect 250591 167023 250639 167051
rect 250329 166989 250639 167023
rect 250329 166961 250377 166989
rect 250405 166961 250439 166989
rect 250467 166961 250501 166989
rect 250529 166961 250563 166989
rect 250591 166961 250639 166989
rect 250329 158175 250639 166961
rect 261664 167175 261824 167192
rect 261664 167147 261699 167175
rect 261727 167147 261761 167175
rect 261789 167147 261824 167175
rect 261664 167113 261824 167147
rect 261664 167085 261699 167113
rect 261727 167085 261761 167113
rect 261789 167085 261824 167113
rect 261664 167051 261824 167085
rect 261664 167023 261699 167051
rect 261727 167023 261761 167051
rect 261789 167023 261824 167051
rect 261664 166989 261824 167023
rect 261664 166961 261699 166989
rect 261727 166961 261761 166989
rect 261789 166961 261824 166989
rect 261664 166944 261824 166961
rect 253984 164175 254144 164192
rect 253984 164147 254019 164175
rect 254047 164147 254081 164175
rect 254109 164147 254144 164175
rect 253984 164113 254144 164147
rect 253984 164085 254019 164113
rect 254047 164085 254081 164113
rect 254109 164085 254144 164113
rect 253984 164051 254144 164085
rect 253984 164023 254019 164051
rect 254047 164023 254081 164051
rect 254109 164023 254144 164051
rect 253984 163989 254144 164023
rect 253984 163961 254019 163989
rect 254047 163961 254081 163989
rect 254109 163961 254144 163989
rect 253984 163944 254144 163961
rect 263829 164175 264139 172961
rect 263829 164147 263877 164175
rect 263905 164147 263939 164175
rect 263967 164147 264001 164175
rect 264029 164147 264063 164175
rect 264091 164147 264139 164175
rect 263829 164113 264139 164147
rect 263829 164085 263877 164113
rect 263905 164085 263939 164113
rect 263967 164085 264001 164113
rect 264029 164085 264063 164113
rect 264091 164085 264139 164113
rect 263829 164051 264139 164085
rect 263829 164023 263877 164051
rect 263905 164023 263939 164051
rect 263967 164023 264001 164051
rect 264029 164023 264063 164051
rect 264091 164023 264139 164051
rect 263829 163989 264139 164023
rect 263829 163961 263877 163989
rect 263905 163961 263939 163989
rect 263967 163961 264001 163989
rect 264029 163961 264063 163989
rect 264091 163961 264139 163989
rect 250329 158147 250377 158175
rect 250405 158147 250439 158175
rect 250467 158147 250501 158175
rect 250529 158147 250563 158175
rect 250591 158147 250639 158175
rect 250329 158113 250639 158147
rect 250329 158085 250377 158113
rect 250405 158085 250439 158113
rect 250467 158085 250501 158113
rect 250529 158085 250563 158113
rect 250591 158085 250639 158113
rect 250329 158051 250639 158085
rect 250329 158023 250377 158051
rect 250405 158023 250439 158051
rect 250467 158023 250501 158051
rect 250529 158023 250563 158051
rect 250591 158023 250639 158051
rect 250329 157989 250639 158023
rect 250329 157961 250377 157989
rect 250405 157961 250439 157989
rect 250467 157961 250501 157989
rect 250529 157961 250563 157989
rect 250591 157961 250639 157989
rect 250329 149175 250639 157961
rect 261664 158175 261824 158192
rect 261664 158147 261699 158175
rect 261727 158147 261761 158175
rect 261789 158147 261824 158175
rect 261664 158113 261824 158147
rect 261664 158085 261699 158113
rect 261727 158085 261761 158113
rect 261789 158085 261824 158113
rect 261664 158051 261824 158085
rect 261664 158023 261699 158051
rect 261727 158023 261761 158051
rect 261789 158023 261824 158051
rect 261664 157989 261824 158023
rect 261664 157961 261699 157989
rect 261727 157961 261761 157989
rect 261789 157961 261824 157989
rect 261664 157944 261824 157961
rect 253984 155175 254144 155192
rect 253984 155147 254019 155175
rect 254047 155147 254081 155175
rect 254109 155147 254144 155175
rect 253984 155113 254144 155147
rect 253984 155085 254019 155113
rect 254047 155085 254081 155113
rect 254109 155085 254144 155113
rect 253984 155051 254144 155085
rect 253984 155023 254019 155051
rect 254047 155023 254081 155051
rect 254109 155023 254144 155051
rect 253984 154989 254144 155023
rect 253984 154961 254019 154989
rect 254047 154961 254081 154989
rect 254109 154961 254144 154989
rect 253984 154944 254144 154961
rect 263829 155175 264139 163961
rect 263829 155147 263877 155175
rect 263905 155147 263939 155175
rect 263967 155147 264001 155175
rect 264029 155147 264063 155175
rect 264091 155147 264139 155175
rect 263829 155113 264139 155147
rect 263829 155085 263877 155113
rect 263905 155085 263939 155113
rect 263967 155085 264001 155113
rect 264029 155085 264063 155113
rect 264091 155085 264139 155113
rect 263829 155051 264139 155085
rect 263829 155023 263877 155051
rect 263905 155023 263939 155051
rect 263967 155023 264001 155051
rect 264029 155023 264063 155051
rect 264091 155023 264139 155051
rect 263829 154989 264139 155023
rect 263829 154961 263877 154989
rect 263905 154961 263939 154989
rect 263967 154961 264001 154989
rect 264029 154961 264063 154989
rect 264091 154961 264139 154989
rect 250329 149147 250377 149175
rect 250405 149147 250439 149175
rect 250467 149147 250501 149175
rect 250529 149147 250563 149175
rect 250591 149147 250639 149175
rect 250329 149113 250639 149147
rect 250329 149085 250377 149113
rect 250405 149085 250439 149113
rect 250467 149085 250501 149113
rect 250529 149085 250563 149113
rect 250591 149085 250639 149113
rect 250329 149051 250639 149085
rect 250329 149023 250377 149051
rect 250405 149023 250439 149051
rect 250467 149023 250501 149051
rect 250529 149023 250563 149051
rect 250591 149023 250639 149051
rect 250329 148989 250639 149023
rect 250329 148961 250377 148989
rect 250405 148961 250439 148989
rect 250467 148961 250501 148989
rect 250529 148961 250563 148989
rect 250591 148961 250639 148989
rect 250329 140175 250639 148961
rect 261664 149175 261824 149192
rect 261664 149147 261699 149175
rect 261727 149147 261761 149175
rect 261789 149147 261824 149175
rect 261664 149113 261824 149147
rect 261664 149085 261699 149113
rect 261727 149085 261761 149113
rect 261789 149085 261824 149113
rect 261664 149051 261824 149085
rect 261664 149023 261699 149051
rect 261727 149023 261761 149051
rect 261789 149023 261824 149051
rect 261664 148989 261824 149023
rect 261664 148961 261699 148989
rect 261727 148961 261761 148989
rect 261789 148961 261824 148989
rect 261664 148944 261824 148961
rect 253984 146175 254144 146192
rect 253984 146147 254019 146175
rect 254047 146147 254081 146175
rect 254109 146147 254144 146175
rect 253984 146113 254144 146147
rect 253984 146085 254019 146113
rect 254047 146085 254081 146113
rect 254109 146085 254144 146113
rect 253984 146051 254144 146085
rect 253984 146023 254019 146051
rect 254047 146023 254081 146051
rect 254109 146023 254144 146051
rect 253984 145989 254144 146023
rect 253984 145961 254019 145989
rect 254047 145961 254081 145989
rect 254109 145961 254144 145989
rect 253984 145944 254144 145961
rect 263829 146175 264139 154961
rect 263829 146147 263877 146175
rect 263905 146147 263939 146175
rect 263967 146147 264001 146175
rect 264029 146147 264063 146175
rect 264091 146147 264139 146175
rect 263829 146113 264139 146147
rect 263829 146085 263877 146113
rect 263905 146085 263939 146113
rect 263967 146085 264001 146113
rect 264029 146085 264063 146113
rect 264091 146085 264139 146113
rect 263829 146051 264139 146085
rect 263829 146023 263877 146051
rect 263905 146023 263939 146051
rect 263967 146023 264001 146051
rect 264029 146023 264063 146051
rect 264091 146023 264139 146051
rect 263829 145989 264139 146023
rect 263829 145961 263877 145989
rect 263905 145961 263939 145989
rect 263967 145961 264001 145989
rect 264029 145961 264063 145989
rect 264091 145961 264139 145989
rect 250329 140147 250377 140175
rect 250405 140147 250439 140175
rect 250467 140147 250501 140175
rect 250529 140147 250563 140175
rect 250591 140147 250639 140175
rect 250329 140113 250639 140147
rect 250329 140085 250377 140113
rect 250405 140085 250439 140113
rect 250467 140085 250501 140113
rect 250529 140085 250563 140113
rect 250591 140085 250639 140113
rect 250329 140051 250639 140085
rect 250329 140023 250377 140051
rect 250405 140023 250439 140051
rect 250467 140023 250501 140051
rect 250529 140023 250563 140051
rect 250591 140023 250639 140051
rect 250329 139989 250639 140023
rect 250329 139961 250377 139989
rect 250405 139961 250439 139989
rect 250467 139961 250501 139989
rect 250529 139961 250563 139989
rect 250591 139961 250639 139989
rect 250329 131175 250639 139961
rect 261664 140175 261824 140192
rect 261664 140147 261699 140175
rect 261727 140147 261761 140175
rect 261789 140147 261824 140175
rect 261664 140113 261824 140147
rect 261664 140085 261699 140113
rect 261727 140085 261761 140113
rect 261789 140085 261824 140113
rect 261664 140051 261824 140085
rect 261664 140023 261699 140051
rect 261727 140023 261761 140051
rect 261789 140023 261824 140051
rect 261664 139989 261824 140023
rect 261664 139961 261699 139989
rect 261727 139961 261761 139989
rect 261789 139961 261824 139989
rect 261664 139944 261824 139961
rect 253984 137175 254144 137192
rect 253984 137147 254019 137175
rect 254047 137147 254081 137175
rect 254109 137147 254144 137175
rect 253984 137113 254144 137147
rect 253984 137085 254019 137113
rect 254047 137085 254081 137113
rect 254109 137085 254144 137113
rect 253984 137051 254144 137085
rect 253984 137023 254019 137051
rect 254047 137023 254081 137051
rect 254109 137023 254144 137051
rect 253984 136989 254144 137023
rect 253984 136961 254019 136989
rect 254047 136961 254081 136989
rect 254109 136961 254144 136989
rect 253984 136944 254144 136961
rect 263829 137175 264139 145961
rect 263829 137147 263877 137175
rect 263905 137147 263939 137175
rect 263967 137147 264001 137175
rect 264029 137147 264063 137175
rect 264091 137147 264139 137175
rect 263829 137113 264139 137147
rect 263829 137085 263877 137113
rect 263905 137085 263939 137113
rect 263967 137085 264001 137113
rect 264029 137085 264063 137113
rect 264091 137085 264139 137113
rect 263829 137051 264139 137085
rect 263829 137023 263877 137051
rect 263905 137023 263939 137051
rect 263967 137023 264001 137051
rect 264029 137023 264063 137051
rect 264091 137023 264139 137051
rect 263829 136989 264139 137023
rect 263829 136961 263877 136989
rect 263905 136961 263939 136989
rect 263967 136961 264001 136989
rect 264029 136961 264063 136989
rect 264091 136961 264139 136989
rect 250329 131147 250377 131175
rect 250405 131147 250439 131175
rect 250467 131147 250501 131175
rect 250529 131147 250563 131175
rect 250591 131147 250639 131175
rect 250329 131113 250639 131147
rect 250329 131085 250377 131113
rect 250405 131085 250439 131113
rect 250467 131085 250501 131113
rect 250529 131085 250563 131113
rect 250591 131085 250639 131113
rect 250329 131051 250639 131085
rect 250329 131023 250377 131051
rect 250405 131023 250439 131051
rect 250467 131023 250501 131051
rect 250529 131023 250563 131051
rect 250591 131023 250639 131051
rect 250329 130989 250639 131023
rect 250329 130961 250377 130989
rect 250405 130961 250439 130989
rect 250467 130961 250501 130989
rect 250529 130961 250563 130989
rect 250591 130961 250639 130989
rect 250329 122175 250639 130961
rect 261664 131175 261824 131192
rect 261664 131147 261699 131175
rect 261727 131147 261761 131175
rect 261789 131147 261824 131175
rect 261664 131113 261824 131147
rect 261664 131085 261699 131113
rect 261727 131085 261761 131113
rect 261789 131085 261824 131113
rect 261664 131051 261824 131085
rect 261664 131023 261699 131051
rect 261727 131023 261761 131051
rect 261789 131023 261824 131051
rect 261664 130989 261824 131023
rect 261664 130961 261699 130989
rect 261727 130961 261761 130989
rect 261789 130961 261824 130989
rect 261664 130944 261824 130961
rect 253984 128175 254144 128192
rect 253984 128147 254019 128175
rect 254047 128147 254081 128175
rect 254109 128147 254144 128175
rect 253984 128113 254144 128147
rect 253984 128085 254019 128113
rect 254047 128085 254081 128113
rect 254109 128085 254144 128113
rect 253984 128051 254144 128085
rect 253984 128023 254019 128051
rect 254047 128023 254081 128051
rect 254109 128023 254144 128051
rect 253984 127989 254144 128023
rect 253984 127961 254019 127989
rect 254047 127961 254081 127989
rect 254109 127961 254144 127989
rect 253984 127944 254144 127961
rect 263829 128175 264139 136961
rect 263829 128147 263877 128175
rect 263905 128147 263939 128175
rect 263967 128147 264001 128175
rect 264029 128147 264063 128175
rect 264091 128147 264139 128175
rect 263829 128113 264139 128147
rect 263829 128085 263877 128113
rect 263905 128085 263939 128113
rect 263967 128085 264001 128113
rect 264029 128085 264063 128113
rect 264091 128085 264139 128113
rect 263829 128051 264139 128085
rect 263829 128023 263877 128051
rect 263905 128023 263939 128051
rect 263967 128023 264001 128051
rect 264029 128023 264063 128051
rect 264091 128023 264139 128051
rect 263829 127989 264139 128023
rect 263829 127961 263877 127989
rect 263905 127961 263939 127989
rect 263967 127961 264001 127989
rect 264029 127961 264063 127989
rect 264091 127961 264139 127989
rect 250329 122147 250377 122175
rect 250405 122147 250439 122175
rect 250467 122147 250501 122175
rect 250529 122147 250563 122175
rect 250591 122147 250639 122175
rect 250329 122113 250639 122147
rect 250329 122085 250377 122113
rect 250405 122085 250439 122113
rect 250467 122085 250501 122113
rect 250529 122085 250563 122113
rect 250591 122085 250639 122113
rect 250329 122051 250639 122085
rect 250329 122023 250377 122051
rect 250405 122023 250439 122051
rect 250467 122023 250501 122051
rect 250529 122023 250563 122051
rect 250591 122023 250639 122051
rect 250329 121989 250639 122023
rect 250329 121961 250377 121989
rect 250405 121961 250439 121989
rect 250467 121961 250501 121989
rect 250529 121961 250563 121989
rect 250591 121961 250639 121989
rect 250329 113175 250639 121961
rect 261664 122175 261824 122192
rect 261664 122147 261699 122175
rect 261727 122147 261761 122175
rect 261789 122147 261824 122175
rect 261664 122113 261824 122147
rect 261664 122085 261699 122113
rect 261727 122085 261761 122113
rect 261789 122085 261824 122113
rect 261664 122051 261824 122085
rect 261664 122023 261699 122051
rect 261727 122023 261761 122051
rect 261789 122023 261824 122051
rect 261664 121989 261824 122023
rect 261664 121961 261699 121989
rect 261727 121961 261761 121989
rect 261789 121961 261824 121989
rect 261664 121944 261824 121961
rect 253984 119175 254144 119192
rect 253984 119147 254019 119175
rect 254047 119147 254081 119175
rect 254109 119147 254144 119175
rect 253984 119113 254144 119147
rect 253984 119085 254019 119113
rect 254047 119085 254081 119113
rect 254109 119085 254144 119113
rect 253984 119051 254144 119085
rect 253984 119023 254019 119051
rect 254047 119023 254081 119051
rect 254109 119023 254144 119051
rect 253984 118989 254144 119023
rect 253984 118961 254019 118989
rect 254047 118961 254081 118989
rect 254109 118961 254144 118989
rect 253984 118944 254144 118961
rect 263829 119175 264139 127961
rect 263829 119147 263877 119175
rect 263905 119147 263939 119175
rect 263967 119147 264001 119175
rect 264029 119147 264063 119175
rect 264091 119147 264139 119175
rect 263829 119113 264139 119147
rect 263829 119085 263877 119113
rect 263905 119085 263939 119113
rect 263967 119085 264001 119113
rect 264029 119085 264063 119113
rect 264091 119085 264139 119113
rect 263829 119051 264139 119085
rect 263829 119023 263877 119051
rect 263905 119023 263939 119051
rect 263967 119023 264001 119051
rect 264029 119023 264063 119051
rect 264091 119023 264139 119051
rect 263829 118989 264139 119023
rect 263829 118961 263877 118989
rect 263905 118961 263939 118989
rect 263967 118961 264001 118989
rect 264029 118961 264063 118989
rect 264091 118961 264139 118989
rect 250329 113147 250377 113175
rect 250405 113147 250439 113175
rect 250467 113147 250501 113175
rect 250529 113147 250563 113175
rect 250591 113147 250639 113175
rect 250329 113113 250639 113147
rect 250329 113085 250377 113113
rect 250405 113085 250439 113113
rect 250467 113085 250501 113113
rect 250529 113085 250563 113113
rect 250591 113085 250639 113113
rect 250329 113051 250639 113085
rect 250329 113023 250377 113051
rect 250405 113023 250439 113051
rect 250467 113023 250501 113051
rect 250529 113023 250563 113051
rect 250591 113023 250639 113051
rect 250329 112989 250639 113023
rect 250329 112961 250377 112989
rect 250405 112961 250439 112989
rect 250467 112961 250501 112989
rect 250529 112961 250563 112989
rect 250591 112961 250639 112989
rect 250329 104175 250639 112961
rect 261664 113175 261824 113192
rect 261664 113147 261699 113175
rect 261727 113147 261761 113175
rect 261789 113147 261824 113175
rect 261664 113113 261824 113147
rect 261664 113085 261699 113113
rect 261727 113085 261761 113113
rect 261789 113085 261824 113113
rect 261664 113051 261824 113085
rect 261664 113023 261699 113051
rect 261727 113023 261761 113051
rect 261789 113023 261824 113051
rect 261664 112989 261824 113023
rect 261664 112961 261699 112989
rect 261727 112961 261761 112989
rect 261789 112961 261824 112989
rect 261664 112944 261824 112961
rect 253984 110175 254144 110192
rect 253984 110147 254019 110175
rect 254047 110147 254081 110175
rect 254109 110147 254144 110175
rect 253984 110113 254144 110147
rect 253984 110085 254019 110113
rect 254047 110085 254081 110113
rect 254109 110085 254144 110113
rect 253984 110051 254144 110085
rect 253984 110023 254019 110051
rect 254047 110023 254081 110051
rect 254109 110023 254144 110051
rect 253984 109989 254144 110023
rect 253984 109961 254019 109989
rect 254047 109961 254081 109989
rect 254109 109961 254144 109989
rect 253984 109944 254144 109961
rect 263829 110175 264139 118961
rect 263829 110147 263877 110175
rect 263905 110147 263939 110175
rect 263967 110147 264001 110175
rect 264029 110147 264063 110175
rect 264091 110147 264139 110175
rect 263829 110113 264139 110147
rect 263829 110085 263877 110113
rect 263905 110085 263939 110113
rect 263967 110085 264001 110113
rect 264029 110085 264063 110113
rect 264091 110085 264139 110113
rect 263829 110051 264139 110085
rect 263829 110023 263877 110051
rect 263905 110023 263939 110051
rect 263967 110023 264001 110051
rect 264029 110023 264063 110051
rect 264091 110023 264139 110051
rect 263829 109989 264139 110023
rect 263829 109961 263877 109989
rect 263905 109961 263939 109989
rect 263967 109961 264001 109989
rect 264029 109961 264063 109989
rect 264091 109961 264139 109989
rect 250329 104147 250377 104175
rect 250405 104147 250439 104175
rect 250467 104147 250501 104175
rect 250529 104147 250563 104175
rect 250591 104147 250639 104175
rect 250329 104113 250639 104147
rect 250329 104085 250377 104113
rect 250405 104085 250439 104113
rect 250467 104085 250501 104113
rect 250529 104085 250563 104113
rect 250591 104085 250639 104113
rect 250329 104051 250639 104085
rect 250329 104023 250377 104051
rect 250405 104023 250439 104051
rect 250467 104023 250501 104051
rect 250529 104023 250563 104051
rect 250591 104023 250639 104051
rect 250329 103989 250639 104023
rect 250329 103961 250377 103989
rect 250405 103961 250439 103989
rect 250467 103961 250501 103989
rect 250529 103961 250563 103989
rect 250591 103961 250639 103989
rect 250329 95175 250639 103961
rect 261664 104175 261824 104192
rect 261664 104147 261699 104175
rect 261727 104147 261761 104175
rect 261789 104147 261824 104175
rect 261664 104113 261824 104147
rect 261664 104085 261699 104113
rect 261727 104085 261761 104113
rect 261789 104085 261824 104113
rect 261664 104051 261824 104085
rect 261664 104023 261699 104051
rect 261727 104023 261761 104051
rect 261789 104023 261824 104051
rect 261664 103989 261824 104023
rect 261664 103961 261699 103989
rect 261727 103961 261761 103989
rect 261789 103961 261824 103989
rect 261664 103944 261824 103961
rect 253984 101175 254144 101192
rect 253984 101147 254019 101175
rect 254047 101147 254081 101175
rect 254109 101147 254144 101175
rect 253984 101113 254144 101147
rect 253984 101085 254019 101113
rect 254047 101085 254081 101113
rect 254109 101085 254144 101113
rect 253984 101051 254144 101085
rect 253984 101023 254019 101051
rect 254047 101023 254081 101051
rect 254109 101023 254144 101051
rect 253984 100989 254144 101023
rect 253984 100961 254019 100989
rect 254047 100961 254081 100989
rect 254109 100961 254144 100989
rect 253984 100944 254144 100961
rect 263829 101175 264139 109961
rect 263829 101147 263877 101175
rect 263905 101147 263939 101175
rect 263967 101147 264001 101175
rect 264029 101147 264063 101175
rect 264091 101147 264139 101175
rect 263829 101113 264139 101147
rect 263829 101085 263877 101113
rect 263905 101085 263939 101113
rect 263967 101085 264001 101113
rect 264029 101085 264063 101113
rect 264091 101085 264139 101113
rect 263829 101051 264139 101085
rect 263829 101023 263877 101051
rect 263905 101023 263939 101051
rect 263967 101023 264001 101051
rect 264029 101023 264063 101051
rect 264091 101023 264139 101051
rect 263829 100989 264139 101023
rect 263829 100961 263877 100989
rect 263905 100961 263939 100989
rect 263967 100961 264001 100989
rect 264029 100961 264063 100989
rect 264091 100961 264139 100989
rect 250329 95147 250377 95175
rect 250405 95147 250439 95175
rect 250467 95147 250501 95175
rect 250529 95147 250563 95175
rect 250591 95147 250639 95175
rect 250329 95113 250639 95147
rect 250329 95085 250377 95113
rect 250405 95085 250439 95113
rect 250467 95085 250501 95113
rect 250529 95085 250563 95113
rect 250591 95085 250639 95113
rect 250329 95051 250639 95085
rect 250329 95023 250377 95051
rect 250405 95023 250439 95051
rect 250467 95023 250501 95051
rect 250529 95023 250563 95051
rect 250591 95023 250639 95051
rect 250329 94989 250639 95023
rect 250329 94961 250377 94989
rect 250405 94961 250439 94989
rect 250467 94961 250501 94989
rect 250529 94961 250563 94989
rect 250591 94961 250639 94989
rect 250329 86175 250639 94961
rect 261664 95175 261824 95192
rect 261664 95147 261699 95175
rect 261727 95147 261761 95175
rect 261789 95147 261824 95175
rect 261664 95113 261824 95147
rect 261664 95085 261699 95113
rect 261727 95085 261761 95113
rect 261789 95085 261824 95113
rect 261664 95051 261824 95085
rect 261664 95023 261699 95051
rect 261727 95023 261761 95051
rect 261789 95023 261824 95051
rect 261664 94989 261824 95023
rect 261664 94961 261699 94989
rect 261727 94961 261761 94989
rect 261789 94961 261824 94989
rect 261664 94944 261824 94961
rect 253984 92175 254144 92192
rect 253984 92147 254019 92175
rect 254047 92147 254081 92175
rect 254109 92147 254144 92175
rect 253984 92113 254144 92147
rect 253984 92085 254019 92113
rect 254047 92085 254081 92113
rect 254109 92085 254144 92113
rect 253984 92051 254144 92085
rect 253984 92023 254019 92051
rect 254047 92023 254081 92051
rect 254109 92023 254144 92051
rect 253984 91989 254144 92023
rect 253984 91961 254019 91989
rect 254047 91961 254081 91989
rect 254109 91961 254144 91989
rect 253984 91944 254144 91961
rect 263829 92175 264139 100961
rect 263829 92147 263877 92175
rect 263905 92147 263939 92175
rect 263967 92147 264001 92175
rect 264029 92147 264063 92175
rect 264091 92147 264139 92175
rect 263829 92113 264139 92147
rect 263829 92085 263877 92113
rect 263905 92085 263939 92113
rect 263967 92085 264001 92113
rect 264029 92085 264063 92113
rect 264091 92085 264139 92113
rect 263829 92051 264139 92085
rect 263829 92023 263877 92051
rect 263905 92023 263939 92051
rect 263967 92023 264001 92051
rect 264029 92023 264063 92051
rect 264091 92023 264139 92051
rect 263829 91989 264139 92023
rect 263829 91961 263877 91989
rect 263905 91961 263939 91989
rect 263967 91961 264001 91989
rect 264029 91961 264063 91989
rect 264091 91961 264139 91989
rect 250329 86147 250377 86175
rect 250405 86147 250439 86175
rect 250467 86147 250501 86175
rect 250529 86147 250563 86175
rect 250591 86147 250639 86175
rect 250329 86113 250639 86147
rect 250329 86085 250377 86113
rect 250405 86085 250439 86113
rect 250467 86085 250501 86113
rect 250529 86085 250563 86113
rect 250591 86085 250639 86113
rect 250329 86051 250639 86085
rect 250329 86023 250377 86051
rect 250405 86023 250439 86051
rect 250467 86023 250501 86051
rect 250529 86023 250563 86051
rect 250591 86023 250639 86051
rect 250329 85989 250639 86023
rect 250329 85961 250377 85989
rect 250405 85961 250439 85989
rect 250467 85961 250501 85989
rect 250529 85961 250563 85989
rect 250591 85961 250639 85989
rect 250329 77175 250639 85961
rect 261664 86175 261824 86192
rect 261664 86147 261699 86175
rect 261727 86147 261761 86175
rect 261789 86147 261824 86175
rect 261664 86113 261824 86147
rect 261664 86085 261699 86113
rect 261727 86085 261761 86113
rect 261789 86085 261824 86113
rect 261664 86051 261824 86085
rect 261664 86023 261699 86051
rect 261727 86023 261761 86051
rect 261789 86023 261824 86051
rect 261664 85989 261824 86023
rect 261664 85961 261699 85989
rect 261727 85961 261761 85989
rect 261789 85961 261824 85989
rect 261664 85944 261824 85961
rect 253984 83175 254144 83192
rect 253984 83147 254019 83175
rect 254047 83147 254081 83175
rect 254109 83147 254144 83175
rect 253984 83113 254144 83147
rect 253984 83085 254019 83113
rect 254047 83085 254081 83113
rect 254109 83085 254144 83113
rect 253984 83051 254144 83085
rect 253984 83023 254019 83051
rect 254047 83023 254081 83051
rect 254109 83023 254144 83051
rect 253984 82989 254144 83023
rect 253984 82961 254019 82989
rect 254047 82961 254081 82989
rect 254109 82961 254144 82989
rect 253984 82944 254144 82961
rect 263829 83175 264139 91961
rect 263829 83147 263877 83175
rect 263905 83147 263939 83175
rect 263967 83147 264001 83175
rect 264029 83147 264063 83175
rect 264091 83147 264139 83175
rect 263829 83113 264139 83147
rect 263829 83085 263877 83113
rect 263905 83085 263939 83113
rect 263967 83085 264001 83113
rect 264029 83085 264063 83113
rect 264091 83085 264139 83113
rect 263829 83051 264139 83085
rect 263829 83023 263877 83051
rect 263905 83023 263939 83051
rect 263967 83023 264001 83051
rect 264029 83023 264063 83051
rect 264091 83023 264139 83051
rect 263829 82989 264139 83023
rect 263829 82961 263877 82989
rect 263905 82961 263939 82989
rect 263967 82961 264001 82989
rect 264029 82961 264063 82989
rect 264091 82961 264139 82989
rect 250329 77147 250377 77175
rect 250405 77147 250439 77175
rect 250467 77147 250501 77175
rect 250529 77147 250563 77175
rect 250591 77147 250639 77175
rect 250329 77113 250639 77147
rect 250329 77085 250377 77113
rect 250405 77085 250439 77113
rect 250467 77085 250501 77113
rect 250529 77085 250563 77113
rect 250591 77085 250639 77113
rect 250329 77051 250639 77085
rect 250329 77023 250377 77051
rect 250405 77023 250439 77051
rect 250467 77023 250501 77051
rect 250529 77023 250563 77051
rect 250591 77023 250639 77051
rect 250329 76989 250639 77023
rect 250329 76961 250377 76989
rect 250405 76961 250439 76989
rect 250467 76961 250501 76989
rect 250529 76961 250563 76989
rect 250591 76961 250639 76989
rect 250329 68175 250639 76961
rect 261664 77175 261824 77192
rect 261664 77147 261699 77175
rect 261727 77147 261761 77175
rect 261789 77147 261824 77175
rect 261664 77113 261824 77147
rect 261664 77085 261699 77113
rect 261727 77085 261761 77113
rect 261789 77085 261824 77113
rect 261664 77051 261824 77085
rect 261664 77023 261699 77051
rect 261727 77023 261761 77051
rect 261789 77023 261824 77051
rect 261664 76989 261824 77023
rect 261664 76961 261699 76989
rect 261727 76961 261761 76989
rect 261789 76961 261824 76989
rect 261664 76944 261824 76961
rect 253984 74175 254144 74192
rect 253984 74147 254019 74175
rect 254047 74147 254081 74175
rect 254109 74147 254144 74175
rect 253984 74113 254144 74147
rect 253984 74085 254019 74113
rect 254047 74085 254081 74113
rect 254109 74085 254144 74113
rect 253984 74051 254144 74085
rect 253984 74023 254019 74051
rect 254047 74023 254081 74051
rect 254109 74023 254144 74051
rect 253984 73989 254144 74023
rect 253984 73961 254019 73989
rect 254047 73961 254081 73989
rect 254109 73961 254144 73989
rect 253984 73944 254144 73961
rect 263829 74175 264139 82961
rect 263829 74147 263877 74175
rect 263905 74147 263939 74175
rect 263967 74147 264001 74175
rect 264029 74147 264063 74175
rect 264091 74147 264139 74175
rect 263829 74113 264139 74147
rect 263829 74085 263877 74113
rect 263905 74085 263939 74113
rect 263967 74085 264001 74113
rect 264029 74085 264063 74113
rect 264091 74085 264139 74113
rect 263829 74051 264139 74085
rect 263829 74023 263877 74051
rect 263905 74023 263939 74051
rect 263967 74023 264001 74051
rect 264029 74023 264063 74051
rect 264091 74023 264139 74051
rect 263829 73989 264139 74023
rect 263829 73961 263877 73989
rect 263905 73961 263939 73989
rect 263967 73961 264001 73989
rect 264029 73961 264063 73989
rect 264091 73961 264139 73989
rect 250329 68147 250377 68175
rect 250405 68147 250439 68175
rect 250467 68147 250501 68175
rect 250529 68147 250563 68175
rect 250591 68147 250639 68175
rect 250329 68113 250639 68147
rect 250329 68085 250377 68113
rect 250405 68085 250439 68113
rect 250467 68085 250501 68113
rect 250529 68085 250563 68113
rect 250591 68085 250639 68113
rect 250329 68051 250639 68085
rect 250329 68023 250377 68051
rect 250405 68023 250439 68051
rect 250467 68023 250501 68051
rect 250529 68023 250563 68051
rect 250591 68023 250639 68051
rect 250329 67989 250639 68023
rect 250329 67961 250377 67989
rect 250405 67961 250439 67989
rect 250467 67961 250501 67989
rect 250529 67961 250563 67989
rect 250591 67961 250639 67989
rect 250329 59175 250639 67961
rect 261664 68175 261824 68192
rect 261664 68147 261699 68175
rect 261727 68147 261761 68175
rect 261789 68147 261824 68175
rect 261664 68113 261824 68147
rect 261664 68085 261699 68113
rect 261727 68085 261761 68113
rect 261789 68085 261824 68113
rect 261664 68051 261824 68085
rect 261664 68023 261699 68051
rect 261727 68023 261761 68051
rect 261789 68023 261824 68051
rect 261664 67989 261824 68023
rect 261664 67961 261699 67989
rect 261727 67961 261761 67989
rect 261789 67961 261824 67989
rect 261664 67944 261824 67961
rect 253984 65175 254144 65192
rect 253984 65147 254019 65175
rect 254047 65147 254081 65175
rect 254109 65147 254144 65175
rect 253984 65113 254144 65147
rect 253984 65085 254019 65113
rect 254047 65085 254081 65113
rect 254109 65085 254144 65113
rect 253984 65051 254144 65085
rect 253984 65023 254019 65051
rect 254047 65023 254081 65051
rect 254109 65023 254144 65051
rect 253984 64989 254144 65023
rect 253984 64961 254019 64989
rect 254047 64961 254081 64989
rect 254109 64961 254144 64989
rect 253984 64944 254144 64961
rect 263829 65175 264139 73961
rect 263829 65147 263877 65175
rect 263905 65147 263939 65175
rect 263967 65147 264001 65175
rect 264029 65147 264063 65175
rect 264091 65147 264139 65175
rect 263829 65113 264139 65147
rect 263829 65085 263877 65113
rect 263905 65085 263939 65113
rect 263967 65085 264001 65113
rect 264029 65085 264063 65113
rect 264091 65085 264139 65113
rect 263829 65051 264139 65085
rect 263829 65023 263877 65051
rect 263905 65023 263939 65051
rect 263967 65023 264001 65051
rect 264029 65023 264063 65051
rect 264091 65023 264139 65051
rect 263829 64989 264139 65023
rect 263829 64961 263877 64989
rect 263905 64961 263939 64989
rect 263967 64961 264001 64989
rect 264029 64961 264063 64989
rect 264091 64961 264139 64989
rect 250329 59147 250377 59175
rect 250405 59147 250439 59175
rect 250467 59147 250501 59175
rect 250529 59147 250563 59175
rect 250591 59147 250639 59175
rect 250329 59113 250639 59147
rect 250329 59085 250377 59113
rect 250405 59085 250439 59113
rect 250467 59085 250501 59113
rect 250529 59085 250563 59113
rect 250591 59085 250639 59113
rect 250329 59051 250639 59085
rect 250329 59023 250377 59051
rect 250405 59023 250439 59051
rect 250467 59023 250501 59051
rect 250529 59023 250563 59051
rect 250591 59023 250639 59051
rect 250329 58989 250639 59023
rect 250329 58961 250377 58989
rect 250405 58961 250439 58989
rect 250467 58961 250501 58989
rect 250529 58961 250563 58989
rect 250591 58961 250639 58989
rect 250329 50175 250639 58961
rect 261664 59175 261824 59192
rect 261664 59147 261699 59175
rect 261727 59147 261761 59175
rect 261789 59147 261824 59175
rect 261664 59113 261824 59147
rect 261664 59085 261699 59113
rect 261727 59085 261761 59113
rect 261789 59085 261824 59113
rect 261664 59051 261824 59085
rect 261664 59023 261699 59051
rect 261727 59023 261761 59051
rect 261789 59023 261824 59051
rect 261664 58989 261824 59023
rect 261664 58961 261699 58989
rect 261727 58961 261761 58989
rect 261789 58961 261824 58989
rect 261664 58944 261824 58961
rect 253984 56175 254144 56192
rect 253984 56147 254019 56175
rect 254047 56147 254081 56175
rect 254109 56147 254144 56175
rect 253984 56113 254144 56147
rect 253984 56085 254019 56113
rect 254047 56085 254081 56113
rect 254109 56085 254144 56113
rect 253984 56051 254144 56085
rect 253984 56023 254019 56051
rect 254047 56023 254081 56051
rect 254109 56023 254144 56051
rect 253984 55989 254144 56023
rect 253984 55961 254019 55989
rect 254047 55961 254081 55989
rect 254109 55961 254144 55989
rect 253984 55944 254144 55961
rect 263829 56175 264139 64961
rect 263829 56147 263877 56175
rect 263905 56147 263939 56175
rect 263967 56147 264001 56175
rect 264029 56147 264063 56175
rect 264091 56147 264139 56175
rect 263829 56113 264139 56147
rect 263829 56085 263877 56113
rect 263905 56085 263939 56113
rect 263967 56085 264001 56113
rect 264029 56085 264063 56113
rect 264091 56085 264139 56113
rect 263829 56051 264139 56085
rect 263829 56023 263877 56051
rect 263905 56023 263939 56051
rect 263967 56023 264001 56051
rect 264029 56023 264063 56051
rect 264091 56023 264139 56051
rect 263829 55989 264139 56023
rect 263829 55961 263877 55989
rect 263905 55961 263939 55989
rect 263967 55961 264001 55989
rect 264029 55961 264063 55989
rect 264091 55961 264139 55989
rect 250329 50147 250377 50175
rect 250405 50147 250439 50175
rect 250467 50147 250501 50175
rect 250529 50147 250563 50175
rect 250591 50147 250639 50175
rect 250329 50113 250639 50147
rect 250329 50085 250377 50113
rect 250405 50085 250439 50113
rect 250467 50085 250501 50113
rect 250529 50085 250563 50113
rect 250591 50085 250639 50113
rect 250329 50051 250639 50085
rect 250329 50023 250377 50051
rect 250405 50023 250439 50051
rect 250467 50023 250501 50051
rect 250529 50023 250563 50051
rect 250591 50023 250639 50051
rect 250329 49989 250639 50023
rect 250329 49961 250377 49989
rect 250405 49961 250439 49989
rect 250467 49961 250501 49989
rect 250529 49961 250563 49989
rect 250591 49961 250639 49989
rect 250329 41175 250639 49961
rect 261664 50175 261824 50192
rect 261664 50147 261699 50175
rect 261727 50147 261761 50175
rect 261789 50147 261824 50175
rect 261664 50113 261824 50147
rect 261664 50085 261699 50113
rect 261727 50085 261761 50113
rect 261789 50085 261824 50113
rect 261664 50051 261824 50085
rect 261664 50023 261699 50051
rect 261727 50023 261761 50051
rect 261789 50023 261824 50051
rect 261664 49989 261824 50023
rect 261664 49961 261699 49989
rect 261727 49961 261761 49989
rect 261789 49961 261824 49989
rect 261664 49944 261824 49961
rect 253984 47175 254144 47192
rect 253984 47147 254019 47175
rect 254047 47147 254081 47175
rect 254109 47147 254144 47175
rect 253984 47113 254144 47147
rect 253984 47085 254019 47113
rect 254047 47085 254081 47113
rect 254109 47085 254144 47113
rect 253984 47051 254144 47085
rect 253984 47023 254019 47051
rect 254047 47023 254081 47051
rect 254109 47023 254144 47051
rect 253984 46989 254144 47023
rect 253984 46961 254019 46989
rect 254047 46961 254081 46989
rect 254109 46961 254144 46989
rect 253984 46944 254144 46961
rect 263829 47175 264139 55961
rect 263829 47147 263877 47175
rect 263905 47147 263939 47175
rect 263967 47147 264001 47175
rect 264029 47147 264063 47175
rect 264091 47147 264139 47175
rect 263829 47113 264139 47147
rect 263829 47085 263877 47113
rect 263905 47085 263939 47113
rect 263967 47085 264001 47113
rect 264029 47085 264063 47113
rect 264091 47085 264139 47113
rect 263829 47051 264139 47085
rect 263829 47023 263877 47051
rect 263905 47023 263939 47051
rect 263967 47023 264001 47051
rect 264029 47023 264063 47051
rect 264091 47023 264139 47051
rect 263829 46989 264139 47023
rect 263829 46961 263877 46989
rect 263905 46961 263939 46989
rect 263967 46961 264001 46989
rect 264029 46961 264063 46989
rect 264091 46961 264139 46989
rect 250329 41147 250377 41175
rect 250405 41147 250439 41175
rect 250467 41147 250501 41175
rect 250529 41147 250563 41175
rect 250591 41147 250639 41175
rect 250329 41113 250639 41147
rect 250329 41085 250377 41113
rect 250405 41085 250439 41113
rect 250467 41085 250501 41113
rect 250529 41085 250563 41113
rect 250591 41085 250639 41113
rect 250329 41051 250639 41085
rect 250329 41023 250377 41051
rect 250405 41023 250439 41051
rect 250467 41023 250501 41051
rect 250529 41023 250563 41051
rect 250591 41023 250639 41051
rect 250329 40989 250639 41023
rect 250329 40961 250377 40989
rect 250405 40961 250439 40989
rect 250467 40961 250501 40989
rect 250529 40961 250563 40989
rect 250591 40961 250639 40989
rect 250329 32175 250639 40961
rect 261664 41175 261824 41192
rect 261664 41147 261699 41175
rect 261727 41147 261761 41175
rect 261789 41147 261824 41175
rect 261664 41113 261824 41147
rect 261664 41085 261699 41113
rect 261727 41085 261761 41113
rect 261789 41085 261824 41113
rect 261664 41051 261824 41085
rect 261664 41023 261699 41051
rect 261727 41023 261761 41051
rect 261789 41023 261824 41051
rect 261664 40989 261824 41023
rect 261664 40961 261699 40989
rect 261727 40961 261761 40989
rect 261789 40961 261824 40989
rect 261664 40944 261824 40961
rect 253984 38175 254144 38192
rect 253984 38147 254019 38175
rect 254047 38147 254081 38175
rect 254109 38147 254144 38175
rect 253984 38113 254144 38147
rect 253984 38085 254019 38113
rect 254047 38085 254081 38113
rect 254109 38085 254144 38113
rect 253984 38051 254144 38085
rect 253984 38023 254019 38051
rect 254047 38023 254081 38051
rect 254109 38023 254144 38051
rect 253984 37989 254144 38023
rect 253984 37961 254019 37989
rect 254047 37961 254081 37989
rect 254109 37961 254144 37989
rect 253984 37944 254144 37961
rect 263829 38175 264139 46961
rect 263829 38147 263877 38175
rect 263905 38147 263939 38175
rect 263967 38147 264001 38175
rect 264029 38147 264063 38175
rect 264091 38147 264139 38175
rect 263829 38113 264139 38147
rect 263829 38085 263877 38113
rect 263905 38085 263939 38113
rect 263967 38085 264001 38113
rect 264029 38085 264063 38113
rect 264091 38085 264139 38113
rect 263829 38051 264139 38085
rect 263829 38023 263877 38051
rect 263905 38023 263939 38051
rect 263967 38023 264001 38051
rect 264029 38023 264063 38051
rect 264091 38023 264139 38051
rect 263829 37989 264139 38023
rect 263829 37961 263877 37989
rect 263905 37961 263939 37989
rect 263967 37961 264001 37989
rect 264029 37961 264063 37989
rect 264091 37961 264139 37989
rect 250329 32147 250377 32175
rect 250405 32147 250439 32175
rect 250467 32147 250501 32175
rect 250529 32147 250563 32175
rect 250591 32147 250639 32175
rect 250329 32113 250639 32147
rect 250329 32085 250377 32113
rect 250405 32085 250439 32113
rect 250467 32085 250501 32113
rect 250529 32085 250563 32113
rect 250591 32085 250639 32113
rect 250329 32051 250639 32085
rect 250329 32023 250377 32051
rect 250405 32023 250439 32051
rect 250467 32023 250501 32051
rect 250529 32023 250563 32051
rect 250591 32023 250639 32051
rect 250329 31989 250639 32023
rect 250329 31961 250377 31989
rect 250405 31961 250439 31989
rect 250467 31961 250501 31989
rect 250529 31961 250563 31989
rect 250591 31961 250639 31989
rect 250329 23175 250639 31961
rect 261664 32175 261824 32192
rect 261664 32147 261699 32175
rect 261727 32147 261761 32175
rect 261789 32147 261824 32175
rect 261664 32113 261824 32147
rect 261664 32085 261699 32113
rect 261727 32085 261761 32113
rect 261789 32085 261824 32113
rect 261664 32051 261824 32085
rect 261664 32023 261699 32051
rect 261727 32023 261761 32051
rect 261789 32023 261824 32051
rect 261664 31989 261824 32023
rect 261664 31961 261699 31989
rect 261727 31961 261761 31989
rect 261789 31961 261824 31989
rect 261664 31944 261824 31961
rect 253984 29175 254144 29192
rect 253984 29147 254019 29175
rect 254047 29147 254081 29175
rect 254109 29147 254144 29175
rect 253984 29113 254144 29147
rect 253984 29085 254019 29113
rect 254047 29085 254081 29113
rect 254109 29085 254144 29113
rect 253984 29051 254144 29085
rect 253984 29023 254019 29051
rect 254047 29023 254081 29051
rect 254109 29023 254144 29051
rect 253984 28989 254144 29023
rect 253984 28961 254019 28989
rect 254047 28961 254081 28989
rect 254109 28961 254144 28989
rect 253984 28944 254144 28961
rect 263829 29175 264139 37961
rect 263829 29147 263877 29175
rect 263905 29147 263939 29175
rect 263967 29147 264001 29175
rect 264029 29147 264063 29175
rect 264091 29147 264139 29175
rect 263829 29113 264139 29147
rect 263829 29085 263877 29113
rect 263905 29085 263939 29113
rect 263967 29085 264001 29113
rect 264029 29085 264063 29113
rect 264091 29085 264139 29113
rect 263829 29051 264139 29085
rect 263829 29023 263877 29051
rect 263905 29023 263939 29051
rect 263967 29023 264001 29051
rect 264029 29023 264063 29051
rect 264091 29023 264139 29051
rect 263829 28989 264139 29023
rect 263829 28961 263877 28989
rect 263905 28961 263939 28989
rect 263967 28961 264001 28989
rect 264029 28961 264063 28989
rect 264091 28961 264139 28989
rect 250329 23147 250377 23175
rect 250405 23147 250439 23175
rect 250467 23147 250501 23175
rect 250529 23147 250563 23175
rect 250591 23147 250639 23175
rect 250329 23113 250639 23147
rect 250329 23085 250377 23113
rect 250405 23085 250439 23113
rect 250467 23085 250501 23113
rect 250529 23085 250563 23113
rect 250591 23085 250639 23113
rect 250329 23051 250639 23085
rect 250329 23023 250377 23051
rect 250405 23023 250439 23051
rect 250467 23023 250501 23051
rect 250529 23023 250563 23051
rect 250591 23023 250639 23051
rect 250329 22989 250639 23023
rect 250329 22961 250377 22989
rect 250405 22961 250439 22989
rect 250467 22961 250501 22989
rect 250529 22961 250563 22989
rect 250591 22961 250639 22989
rect 250329 14175 250639 22961
rect 261664 23175 261824 23192
rect 261664 23147 261699 23175
rect 261727 23147 261761 23175
rect 261789 23147 261824 23175
rect 261664 23113 261824 23147
rect 261664 23085 261699 23113
rect 261727 23085 261761 23113
rect 261789 23085 261824 23113
rect 261664 23051 261824 23085
rect 261664 23023 261699 23051
rect 261727 23023 261761 23051
rect 261789 23023 261824 23051
rect 261664 22989 261824 23023
rect 261664 22961 261699 22989
rect 261727 22961 261761 22989
rect 261789 22961 261824 22989
rect 261664 22944 261824 22961
rect 253984 20175 254144 20192
rect 253984 20147 254019 20175
rect 254047 20147 254081 20175
rect 254109 20147 254144 20175
rect 253984 20113 254144 20147
rect 253984 20085 254019 20113
rect 254047 20085 254081 20113
rect 254109 20085 254144 20113
rect 253984 20051 254144 20085
rect 253984 20023 254019 20051
rect 254047 20023 254081 20051
rect 254109 20023 254144 20051
rect 253984 19989 254144 20023
rect 253984 19961 254019 19989
rect 254047 19961 254081 19989
rect 254109 19961 254144 19989
rect 253984 19944 254144 19961
rect 263829 20175 264139 28961
rect 263829 20147 263877 20175
rect 263905 20147 263939 20175
rect 263967 20147 264001 20175
rect 264029 20147 264063 20175
rect 264091 20147 264139 20175
rect 263829 20113 264139 20147
rect 263829 20085 263877 20113
rect 263905 20085 263939 20113
rect 263967 20085 264001 20113
rect 264029 20085 264063 20113
rect 264091 20085 264139 20113
rect 263829 20051 264139 20085
rect 263829 20023 263877 20051
rect 263905 20023 263939 20051
rect 263967 20023 264001 20051
rect 264029 20023 264063 20051
rect 264091 20023 264139 20051
rect 263829 19989 264139 20023
rect 263829 19961 263877 19989
rect 263905 19961 263939 19989
rect 263967 19961 264001 19989
rect 264029 19961 264063 19989
rect 264091 19961 264139 19989
rect 250329 14147 250377 14175
rect 250405 14147 250439 14175
rect 250467 14147 250501 14175
rect 250529 14147 250563 14175
rect 250591 14147 250639 14175
rect 250329 14113 250639 14147
rect 250329 14085 250377 14113
rect 250405 14085 250439 14113
rect 250467 14085 250501 14113
rect 250529 14085 250563 14113
rect 250591 14085 250639 14113
rect 250329 14051 250639 14085
rect 250329 14023 250377 14051
rect 250405 14023 250439 14051
rect 250467 14023 250501 14051
rect 250529 14023 250563 14051
rect 250591 14023 250639 14051
rect 250329 13989 250639 14023
rect 250329 13961 250377 13989
rect 250405 13961 250439 13989
rect 250467 13961 250501 13989
rect 250529 13961 250563 13989
rect 250591 13961 250639 13989
rect 250329 5175 250639 13961
rect 261664 14175 261824 14192
rect 261664 14147 261699 14175
rect 261727 14147 261761 14175
rect 261789 14147 261824 14175
rect 261664 14113 261824 14147
rect 261664 14085 261699 14113
rect 261727 14085 261761 14113
rect 261789 14085 261824 14113
rect 261664 14051 261824 14085
rect 261664 14023 261699 14051
rect 261727 14023 261761 14051
rect 261789 14023 261824 14051
rect 261664 13989 261824 14023
rect 261664 13961 261699 13989
rect 261727 13961 261761 13989
rect 261789 13961 261824 13989
rect 261664 13944 261824 13961
rect 253984 11175 254144 11192
rect 253984 11147 254019 11175
rect 254047 11147 254081 11175
rect 254109 11147 254144 11175
rect 253984 11113 254144 11147
rect 253984 11085 254019 11113
rect 254047 11085 254081 11113
rect 254109 11085 254144 11113
rect 253984 11051 254144 11085
rect 253984 11023 254019 11051
rect 254047 11023 254081 11051
rect 254109 11023 254144 11051
rect 253984 10989 254144 11023
rect 253984 10961 254019 10989
rect 254047 10961 254081 10989
rect 254109 10961 254144 10989
rect 253984 10944 254144 10961
rect 263829 11175 264139 19961
rect 263829 11147 263877 11175
rect 263905 11147 263939 11175
rect 263967 11147 264001 11175
rect 264029 11147 264063 11175
rect 264091 11147 264139 11175
rect 263829 11113 264139 11147
rect 263829 11085 263877 11113
rect 263905 11085 263939 11113
rect 263967 11085 264001 11113
rect 264029 11085 264063 11113
rect 264091 11085 264139 11113
rect 263829 11051 264139 11085
rect 263829 11023 263877 11051
rect 263905 11023 263939 11051
rect 263967 11023 264001 11051
rect 264029 11023 264063 11051
rect 264091 11023 264139 11051
rect 263829 10989 264139 11023
rect 263829 10961 263877 10989
rect 263905 10961 263939 10989
rect 263967 10961 264001 10989
rect 264029 10961 264063 10989
rect 264091 10961 264139 10989
rect 250329 5147 250377 5175
rect 250405 5147 250439 5175
rect 250467 5147 250501 5175
rect 250529 5147 250563 5175
rect 250591 5147 250639 5175
rect 250329 5113 250639 5147
rect 250329 5085 250377 5113
rect 250405 5085 250439 5113
rect 250467 5085 250501 5113
rect 250529 5085 250563 5113
rect 250591 5085 250639 5113
rect 250329 5051 250639 5085
rect 250329 5023 250377 5051
rect 250405 5023 250439 5051
rect 250467 5023 250501 5051
rect 250529 5023 250563 5051
rect 250591 5023 250639 5051
rect 250329 4989 250639 5023
rect 250329 4961 250377 4989
rect 250405 4961 250439 4989
rect 250467 4961 250501 4989
rect 250529 4961 250563 4989
rect 250591 4961 250639 4989
rect 250329 -560 250639 4961
rect 261664 5175 261824 5192
rect 261664 5147 261699 5175
rect 261727 5147 261761 5175
rect 261789 5147 261824 5175
rect 261664 5113 261824 5147
rect 261664 5085 261699 5113
rect 261727 5085 261761 5113
rect 261789 5085 261824 5113
rect 261664 5051 261824 5085
rect 261664 5023 261699 5051
rect 261727 5023 261761 5051
rect 261789 5023 261824 5051
rect 261664 4989 261824 5023
rect 261664 4961 261699 4989
rect 261727 4961 261761 4989
rect 261789 4961 261824 4989
rect 261664 4944 261824 4961
rect 250329 -588 250377 -560
rect 250405 -588 250439 -560
rect 250467 -588 250501 -560
rect 250529 -588 250563 -560
rect 250591 -588 250639 -560
rect 250329 -622 250639 -588
rect 250329 -650 250377 -622
rect 250405 -650 250439 -622
rect 250467 -650 250501 -622
rect 250529 -650 250563 -622
rect 250591 -650 250639 -622
rect 250329 -684 250639 -650
rect 250329 -712 250377 -684
rect 250405 -712 250439 -684
rect 250467 -712 250501 -684
rect 250529 -712 250563 -684
rect 250591 -712 250639 -684
rect 250329 -746 250639 -712
rect 250329 -774 250377 -746
rect 250405 -774 250439 -746
rect 250467 -774 250501 -746
rect 250529 -774 250563 -746
rect 250591 -774 250639 -746
rect 250329 -822 250639 -774
rect 263829 2175 264139 10961
rect 263829 2147 263877 2175
rect 263905 2147 263939 2175
rect 263967 2147 264001 2175
rect 264029 2147 264063 2175
rect 264091 2147 264139 2175
rect 263829 2113 264139 2147
rect 263829 2085 263877 2113
rect 263905 2085 263939 2113
rect 263967 2085 264001 2113
rect 264029 2085 264063 2113
rect 264091 2085 264139 2113
rect 263829 2051 264139 2085
rect 263829 2023 263877 2051
rect 263905 2023 263939 2051
rect 263967 2023 264001 2051
rect 264029 2023 264063 2051
rect 264091 2023 264139 2051
rect 263829 1989 264139 2023
rect 263829 1961 263877 1989
rect 263905 1961 263939 1989
rect 263967 1961 264001 1989
rect 264029 1961 264063 1989
rect 264091 1961 264139 1989
rect 263829 -80 264139 1961
rect 263829 -108 263877 -80
rect 263905 -108 263939 -80
rect 263967 -108 264001 -80
rect 264029 -108 264063 -80
rect 264091 -108 264139 -80
rect 263829 -142 264139 -108
rect 263829 -170 263877 -142
rect 263905 -170 263939 -142
rect 263967 -170 264001 -142
rect 264029 -170 264063 -142
rect 264091 -170 264139 -142
rect 263829 -204 264139 -170
rect 263829 -232 263877 -204
rect 263905 -232 263939 -204
rect 263967 -232 264001 -204
rect 264029 -232 264063 -204
rect 264091 -232 264139 -204
rect 263829 -266 264139 -232
rect 263829 -294 263877 -266
rect 263905 -294 263939 -266
rect 263967 -294 264001 -266
rect 264029 -294 264063 -266
rect 264091 -294 264139 -266
rect 263829 -822 264139 -294
rect 265689 299086 265999 299134
rect 265689 299058 265737 299086
rect 265765 299058 265799 299086
rect 265827 299058 265861 299086
rect 265889 299058 265923 299086
rect 265951 299058 265999 299086
rect 265689 299024 265999 299058
rect 265689 298996 265737 299024
rect 265765 298996 265799 299024
rect 265827 298996 265861 299024
rect 265889 298996 265923 299024
rect 265951 298996 265999 299024
rect 265689 298962 265999 298996
rect 265689 298934 265737 298962
rect 265765 298934 265799 298962
rect 265827 298934 265861 298962
rect 265889 298934 265923 298962
rect 265951 298934 265999 298962
rect 265689 298900 265999 298934
rect 265689 298872 265737 298900
rect 265765 298872 265799 298900
rect 265827 298872 265861 298900
rect 265889 298872 265923 298900
rect 265951 298872 265999 298900
rect 265689 293175 265999 298872
rect 265689 293147 265737 293175
rect 265765 293147 265799 293175
rect 265827 293147 265861 293175
rect 265889 293147 265923 293175
rect 265951 293147 265999 293175
rect 265689 293113 265999 293147
rect 265689 293085 265737 293113
rect 265765 293085 265799 293113
rect 265827 293085 265861 293113
rect 265889 293085 265923 293113
rect 265951 293085 265999 293113
rect 265689 293051 265999 293085
rect 265689 293023 265737 293051
rect 265765 293023 265799 293051
rect 265827 293023 265861 293051
rect 265889 293023 265923 293051
rect 265951 293023 265999 293051
rect 265689 292989 265999 293023
rect 265689 292961 265737 292989
rect 265765 292961 265799 292989
rect 265827 292961 265861 292989
rect 265889 292961 265923 292989
rect 265951 292961 265999 292989
rect 265689 284175 265999 292961
rect 265689 284147 265737 284175
rect 265765 284147 265799 284175
rect 265827 284147 265861 284175
rect 265889 284147 265923 284175
rect 265951 284147 265999 284175
rect 265689 284113 265999 284147
rect 265689 284085 265737 284113
rect 265765 284085 265799 284113
rect 265827 284085 265861 284113
rect 265889 284085 265923 284113
rect 265951 284085 265999 284113
rect 265689 284051 265999 284085
rect 265689 284023 265737 284051
rect 265765 284023 265799 284051
rect 265827 284023 265861 284051
rect 265889 284023 265923 284051
rect 265951 284023 265999 284051
rect 265689 283989 265999 284023
rect 265689 283961 265737 283989
rect 265765 283961 265799 283989
rect 265827 283961 265861 283989
rect 265889 283961 265923 283989
rect 265951 283961 265999 283989
rect 265689 275175 265999 283961
rect 265689 275147 265737 275175
rect 265765 275147 265799 275175
rect 265827 275147 265861 275175
rect 265889 275147 265923 275175
rect 265951 275147 265999 275175
rect 265689 275113 265999 275147
rect 265689 275085 265737 275113
rect 265765 275085 265799 275113
rect 265827 275085 265861 275113
rect 265889 275085 265923 275113
rect 265951 275085 265999 275113
rect 265689 275051 265999 275085
rect 265689 275023 265737 275051
rect 265765 275023 265799 275051
rect 265827 275023 265861 275051
rect 265889 275023 265923 275051
rect 265951 275023 265999 275051
rect 265689 274989 265999 275023
rect 265689 274961 265737 274989
rect 265765 274961 265799 274989
rect 265827 274961 265861 274989
rect 265889 274961 265923 274989
rect 265951 274961 265999 274989
rect 265689 266175 265999 274961
rect 265689 266147 265737 266175
rect 265765 266147 265799 266175
rect 265827 266147 265861 266175
rect 265889 266147 265923 266175
rect 265951 266147 265999 266175
rect 265689 266113 265999 266147
rect 265689 266085 265737 266113
rect 265765 266085 265799 266113
rect 265827 266085 265861 266113
rect 265889 266085 265923 266113
rect 265951 266085 265999 266113
rect 265689 266051 265999 266085
rect 265689 266023 265737 266051
rect 265765 266023 265799 266051
rect 265827 266023 265861 266051
rect 265889 266023 265923 266051
rect 265951 266023 265999 266051
rect 265689 265989 265999 266023
rect 265689 265961 265737 265989
rect 265765 265961 265799 265989
rect 265827 265961 265861 265989
rect 265889 265961 265923 265989
rect 265951 265961 265999 265989
rect 265689 257175 265999 265961
rect 265689 257147 265737 257175
rect 265765 257147 265799 257175
rect 265827 257147 265861 257175
rect 265889 257147 265923 257175
rect 265951 257147 265999 257175
rect 265689 257113 265999 257147
rect 265689 257085 265737 257113
rect 265765 257085 265799 257113
rect 265827 257085 265861 257113
rect 265889 257085 265923 257113
rect 265951 257085 265999 257113
rect 265689 257051 265999 257085
rect 265689 257023 265737 257051
rect 265765 257023 265799 257051
rect 265827 257023 265861 257051
rect 265889 257023 265923 257051
rect 265951 257023 265999 257051
rect 265689 256989 265999 257023
rect 265689 256961 265737 256989
rect 265765 256961 265799 256989
rect 265827 256961 265861 256989
rect 265889 256961 265923 256989
rect 265951 256961 265999 256989
rect 265689 248175 265999 256961
rect 265689 248147 265737 248175
rect 265765 248147 265799 248175
rect 265827 248147 265861 248175
rect 265889 248147 265923 248175
rect 265951 248147 265999 248175
rect 265689 248113 265999 248147
rect 265689 248085 265737 248113
rect 265765 248085 265799 248113
rect 265827 248085 265861 248113
rect 265889 248085 265923 248113
rect 265951 248085 265999 248113
rect 265689 248051 265999 248085
rect 265689 248023 265737 248051
rect 265765 248023 265799 248051
rect 265827 248023 265861 248051
rect 265889 248023 265923 248051
rect 265951 248023 265999 248051
rect 265689 247989 265999 248023
rect 265689 247961 265737 247989
rect 265765 247961 265799 247989
rect 265827 247961 265861 247989
rect 265889 247961 265923 247989
rect 265951 247961 265999 247989
rect 265689 239175 265999 247961
rect 265689 239147 265737 239175
rect 265765 239147 265799 239175
rect 265827 239147 265861 239175
rect 265889 239147 265923 239175
rect 265951 239147 265999 239175
rect 265689 239113 265999 239147
rect 265689 239085 265737 239113
rect 265765 239085 265799 239113
rect 265827 239085 265861 239113
rect 265889 239085 265923 239113
rect 265951 239085 265999 239113
rect 265689 239051 265999 239085
rect 265689 239023 265737 239051
rect 265765 239023 265799 239051
rect 265827 239023 265861 239051
rect 265889 239023 265923 239051
rect 265951 239023 265999 239051
rect 265689 238989 265999 239023
rect 265689 238961 265737 238989
rect 265765 238961 265799 238989
rect 265827 238961 265861 238989
rect 265889 238961 265923 238989
rect 265951 238961 265999 238989
rect 265689 230175 265999 238961
rect 265689 230147 265737 230175
rect 265765 230147 265799 230175
rect 265827 230147 265861 230175
rect 265889 230147 265923 230175
rect 265951 230147 265999 230175
rect 265689 230113 265999 230147
rect 265689 230085 265737 230113
rect 265765 230085 265799 230113
rect 265827 230085 265861 230113
rect 265889 230085 265923 230113
rect 265951 230085 265999 230113
rect 265689 230051 265999 230085
rect 265689 230023 265737 230051
rect 265765 230023 265799 230051
rect 265827 230023 265861 230051
rect 265889 230023 265923 230051
rect 265951 230023 265999 230051
rect 265689 229989 265999 230023
rect 265689 229961 265737 229989
rect 265765 229961 265799 229989
rect 265827 229961 265861 229989
rect 265889 229961 265923 229989
rect 265951 229961 265999 229989
rect 265689 221175 265999 229961
rect 265689 221147 265737 221175
rect 265765 221147 265799 221175
rect 265827 221147 265861 221175
rect 265889 221147 265923 221175
rect 265951 221147 265999 221175
rect 265689 221113 265999 221147
rect 265689 221085 265737 221113
rect 265765 221085 265799 221113
rect 265827 221085 265861 221113
rect 265889 221085 265923 221113
rect 265951 221085 265999 221113
rect 265689 221051 265999 221085
rect 265689 221023 265737 221051
rect 265765 221023 265799 221051
rect 265827 221023 265861 221051
rect 265889 221023 265923 221051
rect 265951 221023 265999 221051
rect 265689 220989 265999 221023
rect 265689 220961 265737 220989
rect 265765 220961 265799 220989
rect 265827 220961 265861 220989
rect 265889 220961 265923 220989
rect 265951 220961 265999 220989
rect 265689 212175 265999 220961
rect 265689 212147 265737 212175
rect 265765 212147 265799 212175
rect 265827 212147 265861 212175
rect 265889 212147 265923 212175
rect 265951 212147 265999 212175
rect 265689 212113 265999 212147
rect 265689 212085 265737 212113
rect 265765 212085 265799 212113
rect 265827 212085 265861 212113
rect 265889 212085 265923 212113
rect 265951 212085 265999 212113
rect 265689 212051 265999 212085
rect 265689 212023 265737 212051
rect 265765 212023 265799 212051
rect 265827 212023 265861 212051
rect 265889 212023 265923 212051
rect 265951 212023 265999 212051
rect 265689 211989 265999 212023
rect 265689 211961 265737 211989
rect 265765 211961 265799 211989
rect 265827 211961 265861 211989
rect 265889 211961 265923 211989
rect 265951 211961 265999 211989
rect 265689 203175 265999 211961
rect 265689 203147 265737 203175
rect 265765 203147 265799 203175
rect 265827 203147 265861 203175
rect 265889 203147 265923 203175
rect 265951 203147 265999 203175
rect 265689 203113 265999 203147
rect 265689 203085 265737 203113
rect 265765 203085 265799 203113
rect 265827 203085 265861 203113
rect 265889 203085 265923 203113
rect 265951 203085 265999 203113
rect 265689 203051 265999 203085
rect 265689 203023 265737 203051
rect 265765 203023 265799 203051
rect 265827 203023 265861 203051
rect 265889 203023 265923 203051
rect 265951 203023 265999 203051
rect 265689 202989 265999 203023
rect 265689 202961 265737 202989
rect 265765 202961 265799 202989
rect 265827 202961 265861 202989
rect 265889 202961 265923 202989
rect 265951 202961 265999 202989
rect 265689 194175 265999 202961
rect 265689 194147 265737 194175
rect 265765 194147 265799 194175
rect 265827 194147 265861 194175
rect 265889 194147 265923 194175
rect 265951 194147 265999 194175
rect 265689 194113 265999 194147
rect 265689 194085 265737 194113
rect 265765 194085 265799 194113
rect 265827 194085 265861 194113
rect 265889 194085 265923 194113
rect 265951 194085 265999 194113
rect 265689 194051 265999 194085
rect 265689 194023 265737 194051
rect 265765 194023 265799 194051
rect 265827 194023 265861 194051
rect 265889 194023 265923 194051
rect 265951 194023 265999 194051
rect 265689 193989 265999 194023
rect 265689 193961 265737 193989
rect 265765 193961 265799 193989
rect 265827 193961 265861 193989
rect 265889 193961 265923 193989
rect 265951 193961 265999 193989
rect 265689 185175 265999 193961
rect 265689 185147 265737 185175
rect 265765 185147 265799 185175
rect 265827 185147 265861 185175
rect 265889 185147 265923 185175
rect 265951 185147 265999 185175
rect 265689 185113 265999 185147
rect 265689 185085 265737 185113
rect 265765 185085 265799 185113
rect 265827 185085 265861 185113
rect 265889 185085 265923 185113
rect 265951 185085 265999 185113
rect 265689 185051 265999 185085
rect 265689 185023 265737 185051
rect 265765 185023 265799 185051
rect 265827 185023 265861 185051
rect 265889 185023 265923 185051
rect 265951 185023 265999 185051
rect 265689 184989 265999 185023
rect 265689 184961 265737 184989
rect 265765 184961 265799 184989
rect 265827 184961 265861 184989
rect 265889 184961 265923 184989
rect 265951 184961 265999 184989
rect 265689 176175 265999 184961
rect 265689 176147 265737 176175
rect 265765 176147 265799 176175
rect 265827 176147 265861 176175
rect 265889 176147 265923 176175
rect 265951 176147 265999 176175
rect 265689 176113 265999 176147
rect 265689 176085 265737 176113
rect 265765 176085 265799 176113
rect 265827 176085 265861 176113
rect 265889 176085 265923 176113
rect 265951 176085 265999 176113
rect 265689 176051 265999 176085
rect 265689 176023 265737 176051
rect 265765 176023 265799 176051
rect 265827 176023 265861 176051
rect 265889 176023 265923 176051
rect 265951 176023 265999 176051
rect 265689 175989 265999 176023
rect 265689 175961 265737 175989
rect 265765 175961 265799 175989
rect 265827 175961 265861 175989
rect 265889 175961 265923 175989
rect 265951 175961 265999 175989
rect 265689 167175 265999 175961
rect 279189 298606 279499 299134
rect 279189 298578 279237 298606
rect 279265 298578 279299 298606
rect 279327 298578 279361 298606
rect 279389 298578 279423 298606
rect 279451 298578 279499 298606
rect 279189 298544 279499 298578
rect 279189 298516 279237 298544
rect 279265 298516 279299 298544
rect 279327 298516 279361 298544
rect 279389 298516 279423 298544
rect 279451 298516 279499 298544
rect 279189 298482 279499 298516
rect 279189 298454 279237 298482
rect 279265 298454 279299 298482
rect 279327 298454 279361 298482
rect 279389 298454 279423 298482
rect 279451 298454 279499 298482
rect 279189 298420 279499 298454
rect 279189 298392 279237 298420
rect 279265 298392 279299 298420
rect 279327 298392 279361 298420
rect 279389 298392 279423 298420
rect 279451 298392 279499 298420
rect 279189 290175 279499 298392
rect 279189 290147 279237 290175
rect 279265 290147 279299 290175
rect 279327 290147 279361 290175
rect 279389 290147 279423 290175
rect 279451 290147 279499 290175
rect 279189 290113 279499 290147
rect 279189 290085 279237 290113
rect 279265 290085 279299 290113
rect 279327 290085 279361 290113
rect 279389 290085 279423 290113
rect 279451 290085 279499 290113
rect 279189 290051 279499 290085
rect 279189 290023 279237 290051
rect 279265 290023 279299 290051
rect 279327 290023 279361 290051
rect 279389 290023 279423 290051
rect 279451 290023 279499 290051
rect 279189 289989 279499 290023
rect 279189 289961 279237 289989
rect 279265 289961 279299 289989
rect 279327 289961 279361 289989
rect 279389 289961 279423 289989
rect 279451 289961 279499 289989
rect 279189 281175 279499 289961
rect 279189 281147 279237 281175
rect 279265 281147 279299 281175
rect 279327 281147 279361 281175
rect 279389 281147 279423 281175
rect 279451 281147 279499 281175
rect 279189 281113 279499 281147
rect 279189 281085 279237 281113
rect 279265 281085 279299 281113
rect 279327 281085 279361 281113
rect 279389 281085 279423 281113
rect 279451 281085 279499 281113
rect 279189 281051 279499 281085
rect 279189 281023 279237 281051
rect 279265 281023 279299 281051
rect 279327 281023 279361 281051
rect 279389 281023 279423 281051
rect 279451 281023 279499 281051
rect 279189 280989 279499 281023
rect 279189 280961 279237 280989
rect 279265 280961 279299 280989
rect 279327 280961 279361 280989
rect 279389 280961 279423 280989
rect 279451 280961 279499 280989
rect 279189 272175 279499 280961
rect 279189 272147 279237 272175
rect 279265 272147 279299 272175
rect 279327 272147 279361 272175
rect 279389 272147 279423 272175
rect 279451 272147 279499 272175
rect 279189 272113 279499 272147
rect 279189 272085 279237 272113
rect 279265 272085 279299 272113
rect 279327 272085 279361 272113
rect 279389 272085 279423 272113
rect 279451 272085 279499 272113
rect 279189 272051 279499 272085
rect 279189 272023 279237 272051
rect 279265 272023 279299 272051
rect 279327 272023 279361 272051
rect 279389 272023 279423 272051
rect 279451 272023 279499 272051
rect 279189 271989 279499 272023
rect 279189 271961 279237 271989
rect 279265 271961 279299 271989
rect 279327 271961 279361 271989
rect 279389 271961 279423 271989
rect 279451 271961 279499 271989
rect 279189 263175 279499 271961
rect 279189 263147 279237 263175
rect 279265 263147 279299 263175
rect 279327 263147 279361 263175
rect 279389 263147 279423 263175
rect 279451 263147 279499 263175
rect 279189 263113 279499 263147
rect 279189 263085 279237 263113
rect 279265 263085 279299 263113
rect 279327 263085 279361 263113
rect 279389 263085 279423 263113
rect 279451 263085 279499 263113
rect 279189 263051 279499 263085
rect 279189 263023 279237 263051
rect 279265 263023 279299 263051
rect 279327 263023 279361 263051
rect 279389 263023 279423 263051
rect 279451 263023 279499 263051
rect 279189 262989 279499 263023
rect 279189 262961 279237 262989
rect 279265 262961 279299 262989
rect 279327 262961 279361 262989
rect 279389 262961 279423 262989
rect 279451 262961 279499 262989
rect 279189 254175 279499 262961
rect 279189 254147 279237 254175
rect 279265 254147 279299 254175
rect 279327 254147 279361 254175
rect 279389 254147 279423 254175
rect 279451 254147 279499 254175
rect 279189 254113 279499 254147
rect 279189 254085 279237 254113
rect 279265 254085 279299 254113
rect 279327 254085 279361 254113
rect 279389 254085 279423 254113
rect 279451 254085 279499 254113
rect 279189 254051 279499 254085
rect 279189 254023 279237 254051
rect 279265 254023 279299 254051
rect 279327 254023 279361 254051
rect 279389 254023 279423 254051
rect 279451 254023 279499 254051
rect 279189 253989 279499 254023
rect 279189 253961 279237 253989
rect 279265 253961 279299 253989
rect 279327 253961 279361 253989
rect 279389 253961 279423 253989
rect 279451 253961 279499 253989
rect 279189 245175 279499 253961
rect 279189 245147 279237 245175
rect 279265 245147 279299 245175
rect 279327 245147 279361 245175
rect 279389 245147 279423 245175
rect 279451 245147 279499 245175
rect 279189 245113 279499 245147
rect 279189 245085 279237 245113
rect 279265 245085 279299 245113
rect 279327 245085 279361 245113
rect 279389 245085 279423 245113
rect 279451 245085 279499 245113
rect 279189 245051 279499 245085
rect 279189 245023 279237 245051
rect 279265 245023 279299 245051
rect 279327 245023 279361 245051
rect 279389 245023 279423 245051
rect 279451 245023 279499 245051
rect 279189 244989 279499 245023
rect 279189 244961 279237 244989
rect 279265 244961 279299 244989
rect 279327 244961 279361 244989
rect 279389 244961 279423 244989
rect 279451 244961 279499 244989
rect 279189 236175 279499 244961
rect 279189 236147 279237 236175
rect 279265 236147 279299 236175
rect 279327 236147 279361 236175
rect 279389 236147 279423 236175
rect 279451 236147 279499 236175
rect 279189 236113 279499 236147
rect 279189 236085 279237 236113
rect 279265 236085 279299 236113
rect 279327 236085 279361 236113
rect 279389 236085 279423 236113
rect 279451 236085 279499 236113
rect 279189 236051 279499 236085
rect 279189 236023 279237 236051
rect 279265 236023 279299 236051
rect 279327 236023 279361 236051
rect 279389 236023 279423 236051
rect 279451 236023 279499 236051
rect 279189 235989 279499 236023
rect 279189 235961 279237 235989
rect 279265 235961 279299 235989
rect 279327 235961 279361 235989
rect 279389 235961 279423 235989
rect 279451 235961 279499 235989
rect 279189 227175 279499 235961
rect 279189 227147 279237 227175
rect 279265 227147 279299 227175
rect 279327 227147 279361 227175
rect 279389 227147 279423 227175
rect 279451 227147 279499 227175
rect 279189 227113 279499 227147
rect 279189 227085 279237 227113
rect 279265 227085 279299 227113
rect 279327 227085 279361 227113
rect 279389 227085 279423 227113
rect 279451 227085 279499 227113
rect 279189 227051 279499 227085
rect 279189 227023 279237 227051
rect 279265 227023 279299 227051
rect 279327 227023 279361 227051
rect 279389 227023 279423 227051
rect 279451 227023 279499 227051
rect 279189 226989 279499 227023
rect 279189 226961 279237 226989
rect 279265 226961 279299 226989
rect 279327 226961 279361 226989
rect 279389 226961 279423 226989
rect 279451 226961 279499 226989
rect 279189 218175 279499 226961
rect 279189 218147 279237 218175
rect 279265 218147 279299 218175
rect 279327 218147 279361 218175
rect 279389 218147 279423 218175
rect 279451 218147 279499 218175
rect 279189 218113 279499 218147
rect 279189 218085 279237 218113
rect 279265 218085 279299 218113
rect 279327 218085 279361 218113
rect 279389 218085 279423 218113
rect 279451 218085 279499 218113
rect 279189 218051 279499 218085
rect 279189 218023 279237 218051
rect 279265 218023 279299 218051
rect 279327 218023 279361 218051
rect 279389 218023 279423 218051
rect 279451 218023 279499 218051
rect 279189 217989 279499 218023
rect 279189 217961 279237 217989
rect 279265 217961 279299 217989
rect 279327 217961 279361 217989
rect 279389 217961 279423 217989
rect 279451 217961 279499 217989
rect 279189 209175 279499 217961
rect 279189 209147 279237 209175
rect 279265 209147 279299 209175
rect 279327 209147 279361 209175
rect 279389 209147 279423 209175
rect 279451 209147 279499 209175
rect 279189 209113 279499 209147
rect 279189 209085 279237 209113
rect 279265 209085 279299 209113
rect 279327 209085 279361 209113
rect 279389 209085 279423 209113
rect 279451 209085 279499 209113
rect 279189 209051 279499 209085
rect 279189 209023 279237 209051
rect 279265 209023 279299 209051
rect 279327 209023 279361 209051
rect 279389 209023 279423 209051
rect 279451 209023 279499 209051
rect 279189 208989 279499 209023
rect 279189 208961 279237 208989
rect 279265 208961 279299 208989
rect 279327 208961 279361 208989
rect 279389 208961 279423 208989
rect 279451 208961 279499 208989
rect 279189 200175 279499 208961
rect 279189 200147 279237 200175
rect 279265 200147 279299 200175
rect 279327 200147 279361 200175
rect 279389 200147 279423 200175
rect 279451 200147 279499 200175
rect 279189 200113 279499 200147
rect 279189 200085 279237 200113
rect 279265 200085 279299 200113
rect 279327 200085 279361 200113
rect 279389 200085 279423 200113
rect 279451 200085 279499 200113
rect 279189 200051 279499 200085
rect 279189 200023 279237 200051
rect 279265 200023 279299 200051
rect 279327 200023 279361 200051
rect 279389 200023 279423 200051
rect 279451 200023 279499 200051
rect 279189 199989 279499 200023
rect 279189 199961 279237 199989
rect 279265 199961 279299 199989
rect 279327 199961 279361 199989
rect 279389 199961 279423 199989
rect 279451 199961 279499 199989
rect 279189 191175 279499 199961
rect 279189 191147 279237 191175
rect 279265 191147 279299 191175
rect 279327 191147 279361 191175
rect 279389 191147 279423 191175
rect 279451 191147 279499 191175
rect 279189 191113 279499 191147
rect 279189 191085 279237 191113
rect 279265 191085 279299 191113
rect 279327 191085 279361 191113
rect 279389 191085 279423 191113
rect 279451 191085 279499 191113
rect 279189 191051 279499 191085
rect 279189 191023 279237 191051
rect 279265 191023 279299 191051
rect 279327 191023 279361 191051
rect 279389 191023 279423 191051
rect 279451 191023 279499 191051
rect 279189 190989 279499 191023
rect 279189 190961 279237 190989
rect 279265 190961 279299 190989
rect 279327 190961 279361 190989
rect 279389 190961 279423 190989
rect 279451 190961 279499 190989
rect 279189 182175 279499 190961
rect 279189 182147 279237 182175
rect 279265 182147 279299 182175
rect 279327 182147 279361 182175
rect 279389 182147 279423 182175
rect 279451 182147 279499 182175
rect 279189 182113 279499 182147
rect 279189 182085 279237 182113
rect 279265 182085 279299 182113
rect 279327 182085 279361 182113
rect 279389 182085 279423 182113
rect 279451 182085 279499 182113
rect 279189 182051 279499 182085
rect 279189 182023 279237 182051
rect 279265 182023 279299 182051
rect 279327 182023 279361 182051
rect 279389 182023 279423 182051
rect 279451 182023 279499 182051
rect 279189 181989 279499 182023
rect 279189 181961 279237 181989
rect 279265 181961 279299 181989
rect 279327 181961 279361 181989
rect 279389 181961 279423 181989
rect 279451 181961 279499 181989
rect 269344 173175 269504 173192
rect 269344 173147 269379 173175
rect 269407 173147 269441 173175
rect 269469 173147 269504 173175
rect 269344 173113 269504 173147
rect 269344 173085 269379 173113
rect 269407 173085 269441 173113
rect 269469 173085 269504 173113
rect 269344 173051 269504 173085
rect 269344 173023 269379 173051
rect 269407 173023 269441 173051
rect 269469 173023 269504 173051
rect 269344 172989 269504 173023
rect 269344 172961 269379 172989
rect 269407 172961 269441 172989
rect 269469 172961 269504 172989
rect 269344 172944 269504 172961
rect 279189 173175 279499 181961
rect 279189 173147 279237 173175
rect 279265 173147 279299 173175
rect 279327 173147 279361 173175
rect 279389 173147 279423 173175
rect 279451 173147 279499 173175
rect 279189 173113 279499 173147
rect 279189 173085 279237 173113
rect 279265 173085 279299 173113
rect 279327 173085 279361 173113
rect 279389 173085 279423 173113
rect 279451 173085 279499 173113
rect 279189 173051 279499 173085
rect 279189 173023 279237 173051
rect 279265 173023 279299 173051
rect 279327 173023 279361 173051
rect 279389 173023 279423 173051
rect 279451 173023 279499 173051
rect 279189 172989 279499 173023
rect 279189 172961 279237 172989
rect 279265 172961 279299 172989
rect 279327 172961 279361 172989
rect 279389 172961 279423 172989
rect 279451 172961 279499 172989
rect 265689 167147 265737 167175
rect 265765 167147 265799 167175
rect 265827 167147 265861 167175
rect 265889 167147 265923 167175
rect 265951 167147 265999 167175
rect 265689 167113 265999 167147
rect 265689 167085 265737 167113
rect 265765 167085 265799 167113
rect 265827 167085 265861 167113
rect 265889 167085 265923 167113
rect 265951 167085 265999 167113
rect 265689 167051 265999 167085
rect 265689 167023 265737 167051
rect 265765 167023 265799 167051
rect 265827 167023 265861 167051
rect 265889 167023 265923 167051
rect 265951 167023 265999 167051
rect 265689 166989 265999 167023
rect 265689 166961 265737 166989
rect 265765 166961 265799 166989
rect 265827 166961 265861 166989
rect 265889 166961 265923 166989
rect 265951 166961 265999 166989
rect 265689 158175 265999 166961
rect 277024 167175 277184 167192
rect 277024 167147 277059 167175
rect 277087 167147 277121 167175
rect 277149 167147 277184 167175
rect 277024 167113 277184 167147
rect 277024 167085 277059 167113
rect 277087 167085 277121 167113
rect 277149 167085 277184 167113
rect 277024 167051 277184 167085
rect 277024 167023 277059 167051
rect 277087 167023 277121 167051
rect 277149 167023 277184 167051
rect 277024 166989 277184 167023
rect 277024 166961 277059 166989
rect 277087 166961 277121 166989
rect 277149 166961 277184 166989
rect 277024 166944 277184 166961
rect 269344 164175 269504 164192
rect 269344 164147 269379 164175
rect 269407 164147 269441 164175
rect 269469 164147 269504 164175
rect 269344 164113 269504 164147
rect 269344 164085 269379 164113
rect 269407 164085 269441 164113
rect 269469 164085 269504 164113
rect 269344 164051 269504 164085
rect 269344 164023 269379 164051
rect 269407 164023 269441 164051
rect 269469 164023 269504 164051
rect 269344 163989 269504 164023
rect 269344 163961 269379 163989
rect 269407 163961 269441 163989
rect 269469 163961 269504 163989
rect 269344 163944 269504 163961
rect 279189 164175 279499 172961
rect 279189 164147 279237 164175
rect 279265 164147 279299 164175
rect 279327 164147 279361 164175
rect 279389 164147 279423 164175
rect 279451 164147 279499 164175
rect 279189 164113 279499 164147
rect 279189 164085 279237 164113
rect 279265 164085 279299 164113
rect 279327 164085 279361 164113
rect 279389 164085 279423 164113
rect 279451 164085 279499 164113
rect 279189 164051 279499 164085
rect 279189 164023 279237 164051
rect 279265 164023 279299 164051
rect 279327 164023 279361 164051
rect 279389 164023 279423 164051
rect 279451 164023 279499 164051
rect 279189 163989 279499 164023
rect 279189 163961 279237 163989
rect 279265 163961 279299 163989
rect 279327 163961 279361 163989
rect 279389 163961 279423 163989
rect 279451 163961 279499 163989
rect 265689 158147 265737 158175
rect 265765 158147 265799 158175
rect 265827 158147 265861 158175
rect 265889 158147 265923 158175
rect 265951 158147 265999 158175
rect 265689 158113 265999 158147
rect 265689 158085 265737 158113
rect 265765 158085 265799 158113
rect 265827 158085 265861 158113
rect 265889 158085 265923 158113
rect 265951 158085 265999 158113
rect 265689 158051 265999 158085
rect 265689 158023 265737 158051
rect 265765 158023 265799 158051
rect 265827 158023 265861 158051
rect 265889 158023 265923 158051
rect 265951 158023 265999 158051
rect 265689 157989 265999 158023
rect 265689 157961 265737 157989
rect 265765 157961 265799 157989
rect 265827 157961 265861 157989
rect 265889 157961 265923 157989
rect 265951 157961 265999 157989
rect 265689 149175 265999 157961
rect 277024 158175 277184 158192
rect 277024 158147 277059 158175
rect 277087 158147 277121 158175
rect 277149 158147 277184 158175
rect 277024 158113 277184 158147
rect 277024 158085 277059 158113
rect 277087 158085 277121 158113
rect 277149 158085 277184 158113
rect 277024 158051 277184 158085
rect 277024 158023 277059 158051
rect 277087 158023 277121 158051
rect 277149 158023 277184 158051
rect 277024 157989 277184 158023
rect 277024 157961 277059 157989
rect 277087 157961 277121 157989
rect 277149 157961 277184 157989
rect 277024 157944 277184 157961
rect 269344 155175 269504 155192
rect 269344 155147 269379 155175
rect 269407 155147 269441 155175
rect 269469 155147 269504 155175
rect 269344 155113 269504 155147
rect 269344 155085 269379 155113
rect 269407 155085 269441 155113
rect 269469 155085 269504 155113
rect 269344 155051 269504 155085
rect 269344 155023 269379 155051
rect 269407 155023 269441 155051
rect 269469 155023 269504 155051
rect 269344 154989 269504 155023
rect 269344 154961 269379 154989
rect 269407 154961 269441 154989
rect 269469 154961 269504 154989
rect 269344 154944 269504 154961
rect 279189 155175 279499 163961
rect 279189 155147 279237 155175
rect 279265 155147 279299 155175
rect 279327 155147 279361 155175
rect 279389 155147 279423 155175
rect 279451 155147 279499 155175
rect 279189 155113 279499 155147
rect 279189 155085 279237 155113
rect 279265 155085 279299 155113
rect 279327 155085 279361 155113
rect 279389 155085 279423 155113
rect 279451 155085 279499 155113
rect 279189 155051 279499 155085
rect 279189 155023 279237 155051
rect 279265 155023 279299 155051
rect 279327 155023 279361 155051
rect 279389 155023 279423 155051
rect 279451 155023 279499 155051
rect 279189 154989 279499 155023
rect 279189 154961 279237 154989
rect 279265 154961 279299 154989
rect 279327 154961 279361 154989
rect 279389 154961 279423 154989
rect 279451 154961 279499 154989
rect 265689 149147 265737 149175
rect 265765 149147 265799 149175
rect 265827 149147 265861 149175
rect 265889 149147 265923 149175
rect 265951 149147 265999 149175
rect 265689 149113 265999 149147
rect 265689 149085 265737 149113
rect 265765 149085 265799 149113
rect 265827 149085 265861 149113
rect 265889 149085 265923 149113
rect 265951 149085 265999 149113
rect 265689 149051 265999 149085
rect 265689 149023 265737 149051
rect 265765 149023 265799 149051
rect 265827 149023 265861 149051
rect 265889 149023 265923 149051
rect 265951 149023 265999 149051
rect 265689 148989 265999 149023
rect 265689 148961 265737 148989
rect 265765 148961 265799 148989
rect 265827 148961 265861 148989
rect 265889 148961 265923 148989
rect 265951 148961 265999 148989
rect 265689 140175 265999 148961
rect 277024 149175 277184 149192
rect 277024 149147 277059 149175
rect 277087 149147 277121 149175
rect 277149 149147 277184 149175
rect 277024 149113 277184 149147
rect 277024 149085 277059 149113
rect 277087 149085 277121 149113
rect 277149 149085 277184 149113
rect 277024 149051 277184 149085
rect 277024 149023 277059 149051
rect 277087 149023 277121 149051
rect 277149 149023 277184 149051
rect 277024 148989 277184 149023
rect 277024 148961 277059 148989
rect 277087 148961 277121 148989
rect 277149 148961 277184 148989
rect 277024 148944 277184 148961
rect 269344 146175 269504 146192
rect 269344 146147 269379 146175
rect 269407 146147 269441 146175
rect 269469 146147 269504 146175
rect 269344 146113 269504 146147
rect 269344 146085 269379 146113
rect 269407 146085 269441 146113
rect 269469 146085 269504 146113
rect 269344 146051 269504 146085
rect 269344 146023 269379 146051
rect 269407 146023 269441 146051
rect 269469 146023 269504 146051
rect 269344 145989 269504 146023
rect 269344 145961 269379 145989
rect 269407 145961 269441 145989
rect 269469 145961 269504 145989
rect 269344 145944 269504 145961
rect 279189 146175 279499 154961
rect 279189 146147 279237 146175
rect 279265 146147 279299 146175
rect 279327 146147 279361 146175
rect 279389 146147 279423 146175
rect 279451 146147 279499 146175
rect 279189 146113 279499 146147
rect 279189 146085 279237 146113
rect 279265 146085 279299 146113
rect 279327 146085 279361 146113
rect 279389 146085 279423 146113
rect 279451 146085 279499 146113
rect 279189 146051 279499 146085
rect 279189 146023 279237 146051
rect 279265 146023 279299 146051
rect 279327 146023 279361 146051
rect 279389 146023 279423 146051
rect 279451 146023 279499 146051
rect 279189 145989 279499 146023
rect 279189 145961 279237 145989
rect 279265 145961 279299 145989
rect 279327 145961 279361 145989
rect 279389 145961 279423 145989
rect 279451 145961 279499 145989
rect 265689 140147 265737 140175
rect 265765 140147 265799 140175
rect 265827 140147 265861 140175
rect 265889 140147 265923 140175
rect 265951 140147 265999 140175
rect 265689 140113 265999 140147
rect 265689 140085 265737 140113
rect 265765 140085 265799 140113
rect 265827 140085 265861 140113
rect 265889 140085 265923 140113
rect 265951 140085 265999 140113
rect 265689 140051 265999 140085
rect 265689 140023 265737 140051
rect 265765 140023 265799 140051
rect 265827 140023 265861 140051
rect 265889 140023 265923 140051
rect 265951 140023 265999 140051
rect 265689 139989 265999 140023
rect 265689 139961 265737 139989
rect 265765 139961 265799 139989
rect 265827 139961 265861 139989
rect 265889 139961 265923 139989
rect 265951 139961 265999 139989
rect 265689 131175 265999 139961
rect 277024 140175 277184 140192
rect 277024 140147 277059 140175
rect 277087 140147 277121 140175
rect 277149 140147 277184 140175
rect 277024 140113 277184 140147
rect 277024 140085 277059 140113
rect 277087 140085 277121 140113
rect 277149 140085 277184 140113
rect 277024 140051 277184 140085
rect 277024 140023 277059 140051
rect 277087 140023 277121 140051
rect 277149 140023 277184 140051
rect 277024 139989 277184 140023
rect 277024 139961 277059 139989
rect 277087 139961 277121 139989
rect 277149 139961 277184 139989
rect 277024 139944 277184 139961
rect 269344 137175 269504 137192
rect 269344 137147 269379 137175
rect 269407 137147 269441 137175
rect 269469 137147 269504 137175
rect 269344 137113 269504 137147
rect 269344 137085 269379 137113
rect 269407 137085 269441 137113
rect 269469 137085 269504 137113
rect 269344 137051 269504 137085
rect 269344 137023 269379 137051
rect 269407 137023 269441 137051
rect 269469 137023 269504 137051
rect 269344 136989 269504 137023
rect 269344 136961 269379 136989
rect 269407 136961 269441 136989
rect 269469 136961 269504 136989
rect 269344 136944 269504 136961
rect 279189 137175 279499 145961
rect 279189 137147 279237 137175
rect 279265 137147 279299 137175
rect 279327 137147 279361 137175
rect 279389 137147 279423 137175
rect 279451 137147 279499 137175
rect 279189 137113 279499 137147
rect 279189 137085 279237 137113
rect 279265 137085 279299 137113
rect 279327 137085 279361 137113
rect 279389 137085 279423 137113
rect 279451 137085 279499 137113
rect 279189 137051 279499 137085
rect 279189 137023 279237 137051
rect 279265 137023 279299 137051
rect 279327 137023 279361 137051
rect 279389 137023 279423 137051
rect 279451 137023 279499 137051
rect 279189 136989 279499 137023
rect 279189 136961 279237 136989
rect 279265 136961 279299 136989
rect 279327 136961 279361 136989
rect 279389 136961 279423 136989
rect 279451 136961 279499 136989
rect 265689 131147 265737 131175
rect 265765 131147 265799 131175
rect 265827 131147 265861 131175
rect 265889 131147 265923 131175
rect 265951 131147 265999 131175
rect 265689 131113 265999 131147
rect 265689 131085 265737 131113
rect 265765 131085 265799 131113
rect 265827 131085 265861 131113
rect 265889 131085 265923 131113
rect 265951 131085 265999 131113
rect 265689 131051 265999 131085
rect 265689 131023 265737 131051
rect 265765 131023 265799 131051
rect 265827 131023 265861 131051
rect 265889 131023 265923 131051
rect 265951 131023 265999 131051
rect 265689 130989 265999 131023
rect 265689 130961 265737 130989
rect 265765 130961 265799 130989
rect 265827 130961 265861 130989
rect 265889 130961 265923 130989
rect 265951 130961 265999 130989
rect 265689 122175 265999 130961
rect 277024 131175 277184 131192
rect 277024 131147 277059 131175
rect 277087 131147 277121 131175
rect 277149 131147 277184 131175
rect 277024 131113 277184 131147
rect 277024 131085 277059 131113
rect 277087 131085 277121 131113
rect 277149 131085 277184 131113
rect 277024 131051 277184 131085
rect 277024 131023 277059 131051
rect 277087 131023 277121 131051
rect 277149 131023 277184 131051
rect 277024 130989 277184 131023
rect 277024 130961 277059 130989
rect 277087 130961 277121 130989
rect 277149 130961 277184 130989
rect 277024 130944 277184 130961
rect 269344 128175 269504 128192
rect 269344 128147 269379 128175
rect 269407 128147 269441 128175
rect 269469 128147 269504 128175
rect 269344 128113 269504 128147
rect 269344 128085 269379 128113
rect 269407 128085 269441 128113
rect 269469 128085 269504 128113
rect 269344 128051 269504 128085
rect 269344 128023 269379 128051
rect 269407 128023 269441 128051
rect 269469 128023 269504 128051
rect 269344 127989 269504 128023
rect 269344 127961 269379 127989
rect 269407 127961 269441 127989
rect 269469 127961 269504 127989
rect 269344 127944 269504 127961
rect 279189 128175 279499 136961
rect 279189 128147 279237 128175
rect 279265 128147 279299 128175
rect 279327 128147 279361 128175
rect 279389 128147 279423 128175
rect 279451 128147 279499 128175
rect 279189 128113 279499 128147
rect 279189 128085 279237 128113
rect 279265 128085 279299 128113
rect 279327 128085 279361 128113
rect 279389 128085 279423 128113
rect 279451 128085 279499 128113
rect 279189 128051 279499 128085
rect 279189 128023 279237 128051
rect 279265 128023 279299 128051
rect 279327 128023 279361 128051
rect 279389 128023 279423 128051
rect 279451 128023 279499 128051
rect 279189 127989 279499 128023
rect 279189 127961 279237 127989
rect 279265 127961 279299 127989
rect 279327 127961 279361 127989
rect 279389 127961 279423 127989
rect 279451 127961 279499 127989
rect 265689 122147 265737 122175
rect 265765 122147 265799 122175
rect 265827 122147 265861 122175
rect 265889 122147 265923 122175
rect 265951 122147 265999 122175
rect 265689 122113 265999 122147
rect 265689 122085 265737 122113
rect 265765 122085 265799 122113
rect 265827 122085 265861 122113
rect 265889 122085 265923 122113
rect 265951 122085 265999 122113
rect 265689 122051 265999 122085
rect 265689 122023 265737 122051
rect 265765 122023 265799 122051
rect 265827 122023 265861 122051
rect 265889 122023 265923 122051
rect 265951 122023 265999 122051
rect 265689 121989 265999 122023
rect 265689 121961 265737 121989
rect 265765 121961 265799 121989
rect 265827 121961 265861 121989
rect 265889 121961 265923 121989
rect 265951 121961 265999 121989
rect 265689 113175 265999 121961
rect 277024 122175 277184 122192
rect 277024 122147 277059 122175
rect 277087 122147 277121 122175
rect 277149 122147 277184 122175
rect 277024 122113 277184 122147
rect 277024 122085 277059 122113
rect 277087 122085 277121 122113
rect 277149 122085 277184 122113
rect 277024 122051 277184 122085
rect 277024 122023 277059 122051
rect 277087 122023 277121 122051
rect 277149 122023 277184 122051
rect 277024 121989 277184 122023
rect 277024 121961 277059 121989
rect 277087 121961 277121 121989
rect 277149 121961 277184 121989
rect 277024 121944 277184 121961
rect 269344 119175 269504 119192
rect 269344 119147 269379 119175
rect 269407 119147 269441 119175
rect 269469 119147 269504 119175
rect 269344 119113 269504 119147
rect 269344 119085 269379 119113
rect 269407 119085 269441 119113
rect 269469 119085 269504 119113
rect 269344 119051 269504 119085
rect 269344 119023 269379 119051
rect 269407 119023 269441 119051
rect 269469 119023 269504 119051
rect 269344 118989 269504 119023
rect 269344 118961 269379 118989
rect 269407 118961 269441 118989
rect 269469 118961 269504 118989
rect 269344 118944 269504 118961
rect 279189 119175 279499 127961
rect 279189 119147 279237 119175
rect 279265 119147 279299 119175
rect 279327 119147 279361 119175
rect 279389 119147 279423 119175
rect 279451 119147 279499 119175
rect 279189 119113 279499 119147
rect 279189 119085 279237 119113
rect 279265 119085 279299 119113
rect 279327 119085 279361 119113
rect 279389 119085 279423 119113
rect 279451 119085 279499 119113
rect 279189 119051 279499 119085
rect 279189 119023 279237 119051
rect 279265 119023 279299 119051
rect 279327 119023 279361 119051
rect 279389 119023 279423 119051
rect 279451 119023 279499 119051
rect 279189 118989 279499 119023
rect 279189 118961 279237 118989
rect 279265 118961 279299 118989
rect 279327 118961 279361 118989
rect 279389 118961 279423 118989
rect 279451 118961 279499 118989
rect 265689 113147 265737 113175
rect 265765 113147 265799 113175
rect 265827 113147 265861 113175
rect 265889 113147 265923 113175
rect 265951 113147 265999 113175
rect 265689 113113 265999 113147
rect 265689 113085 265737 113113
rect 265765 113085 265799 113113
rect 265827 113085 265861 113113
rect 265889 113085 265923 113113
rect 265951 113085 265999 113113
rect 265689 113051 265999 113085
rect 265689 113023 265737 113051
rect 265765 113023 265799 113051
rect 265827 113023 265861 113051
rect 265889 113023 265923 113051
rect 265951 113023 265999 113051
rect 265689 112989 265999 113023
rect 265689 112961 265737 112989
rect 265765 112961 265799 112989
rect 265827 112961 265861 112989
rect 265889 112961 265923 112989
rect 265951 112961 265999 112989
rect 265689 104175 265999 112961
rect 277024 113175 277184 113192
rect 277024 113147 277059 113175
rect 277087 113147 277121 113175
rect 277149 113147 277184 113175
rect 277024 113113 277184 113147
rect 277024 113085 277059 113113
rect 277087 113085 277121 113113
rect 277149 113085 277184 113113
rect 277024 113051 277184 113085
rect 277024 113023 277059 113051
rect 277087 113023 277121 113051
rect 277149 113023 277184 113051
rect 277024 112989 277184 113023
rect 277024 112961 277059 112989
rect 277087 112961 277121 112989
rect 277149 112961 277184 112989
rect 277024 112944 277184 112961
rect 269344 110175 269504 110192
rect 269344 110147 269379 110175
rect 269407 110147 269441 110175
rect 269469 110147 269504 110175
rect 269344 110113 269504 110147
rect 269344 110085 269379 110113
rect 269407 110085 269441 110113
rect 269469 110085 269504 110113
rect 269344 110051 269504 110085
rect 269344 110023 269379 110051
rect 269407 110023 269441 110051
rect 269469 110023 269504 110051
rect 269344 109989 269504 110023
rect 269344 109961 269379 109989
rect 269407 109961 269441 109989
rect 269469 109961 269504 109989
rect 269344 109944 269504 109961
rect 279189 110175 279499 118961
rect 279189 110147 279237 110175
rect 279265 110147 279299 110175
rect 279327 110147 279361 110175
rect 279389 110147 279423 110175
rect 279451 110147 279499 110175
rect 279189 110113 279499 110147
rect 279189 110085 279237 110113
rect 279265 110085 279299 110113
rect 279327 110085 279361 110113
rect 279389 110085 279423 110113
rect 279451 110085 279499 110113
rect 279189 110051 279499 110085
rect 279189 110023 279237 110051
rect 279265 110023 279299 110051
rect 279327 110023 279361 110051
rect 279389 110023 279423 110051
rect 279451 110023 279499 110051
rect 279189 109989 279499 110023
rect 279189 109961 279237 109989
rect 279265 109961 279299 109989
rect 279327 109961 279361 109989
rect 279389 109961 279423 109989
rect 279451 109961 279499 109989
rect 265689 104147 265737 104175
rect 265765 104147 265799 104175
rect 265827 104147 265861 104175
rect 265889 104147 265923 104175
rect 265951 104147 265999 104175
rect 265689 104113 265999 104147
rect 265689 104085 265737 104113
rect 265765 104085 265799 104113
rect 265827 104085 265861 104113
rect 265889 104085 265923 104113
rect 265951 104085 265999 104113
rect 265689 104051 265999 104085
rect 265689 104023 265737 104051
rect 265765 104023 265799 104051
rect 265827 104023 265861 104051
rect 265889 104023 265923 104051
rect 265951 104023 265999 104051
rect 265689 103989 265999 104023
rect 265689 103961 265737 103989
rect 265765 103961 265799 103989
rect 265827 103961 265861 103989
rect 265889 103961 265923 103989
rect 265951 103961 265999 103989
rect 265689 95175 265999 103961
rect 277024 104175 277184 104192
rect 277024 104147 277059 104175
rect 277087 104147 277121 104175
rect 277149 104147 277184 104175
rect 277024 104113 277184 104147
rect 277024 104085 277059 104113
rect 277087 104085 277121 104113
rect 277149 104085 277184 104113
rect 277024 104051 277184 104085
rect 277024 104023 277059 104051
rect 277087 104023 277121 104051
rect 277149 104023 277184 104051
rect 277024 103989 277184 104023
rect 277024 103961 277059 103989
rect 277087 103961 277121 103989
rect 277149 103961 277184 103989
rect 277024 103944 277184 103961
rect 269344 101175 269504 101192
rect 269344 101147 269379 101175
rect 269407 101147 269441 101175
rect 269469 101147 269504 101175
rect 269344 101113 269504 101147
rect 269344 101085 269379 101113
rect 269407 101085 269441 101113
rect 269469 101085 269504 101113
rect 269344 101051 269504 101085
rect 269344 101023 269379 101051
rect 269407 101023 269441 101051
rect 269469 101023 269504 101051
rect 269344 100989 269504 101023
rect 269344 100961 269379 100989
rect 269407 100961 269441 100989
rect 269469 100961 269504 100989
rect 269344 100944 269504 100961
rect 279189 101175 279499 109961
rect 279189 101147 279237 101175
rect 279265 101147 279299 101175
rect 279327 101147 279361 101175
rect 279389 101147 279423 101175
rect 279451 101147 279499 101175
rect 279189 101113 279499 101147
rect 279189 101085 279237 101113
rect 279265 101085 279299 101113
rect 279327 101085 279361 101113
rect 279389 101085 279423 101113
rect 279451 101085 279499 101113
rect 279189 101051 279499 101085
rect 279189 101023 279237 101051
rect 279265 101023 279299 101051
rect 279327 101023 279361 101051
rect 279389 101023 279423 101051
rect 279451 101023 279499 101051
rect 279189 100989 279499 101023
rect 279189 100961 279237 100989
rect 279265 100961 279299 100989
rect 279327 100961 279361 100989
rect 279389 100961 279423 100989
rect 279451 100961 279499 100989
rect 265689 95147 265737 95175
rect 265765 95147 265799 95175
rect 265827 95147 265861 95175
rect 265889 95147 265923 95175
rect 265951 95147 265999 95175
rect 265689 95113 265999 95147
rect 265689 95085 265737 95113
rect 265765 95085 265799 95113
rect 265827 95085 265861 95113
rect 265889 95085 265923 95113
rect 265951 95085 265999 95113
rect 265689 95051 265999 95085
rect 265689 95023 265737 95051
rect 265765 95023 265799 95051
rect 265827 95023 265861 95051
rect 265889 95023 265923 95051
rect 265951 95023 265999 95051
rect 265689 94989 265999 95023
rect 265689 94961 265737 94989
rect 265765 94961 265799 94989
rect 265827 94961 265861 94989
rect 265889 94961 265923 94989
rect 265951 94961 265999 94989
rect 265689 86175 265999 94961
rect 277024 95175 277184 95192
rect 277024 95147 277059 95175
rect 277087 95147 277121 95175
rect 277149 95147 277184 95175
rect 277024 95113 277184 95147
rect 277024 95085 277059 95113
rect 277087 95085 277121 95113
rect 277149 95085 277184 95113
rect 277024 95051 277184 95085
rect 277024 95023 277059 95051
rect 277087 95023 277121 95051
rect 277149 95023 277184 95051
rect 277024 94989 277184 95023
rect 277024 94961 277059 94989
rect 277087 94961 277121 94989
rect 277149 94961 277184 94989
rect 277024 94944 277184 94961
rect 269344 92175 269504 92192
rect 269344 92147 269379 92175
rect 269407 92147 269441 92175
rect 269469 92147 269504 92175
rect 269344 92113 269504 92147
rect 269344 92085 269379 92113
rect 269407 92085 269441 92113
rect 269469 92085 269504 92113
rect 269344 92051 269504 92085
rect 269344 92023 269379 92051
rect 269407 92023 269441 92051
rect 269469 92023 269504 92051
rect 269344 91989 269504 92023
rect 269344 91961 269379 91989
rect 269407 91961 269441 91989
rect 269469 91961 269504 91989
rect 269344 91944 269504 91961
rect 279189 92175 279499 100961
rect 279189 92147 279237 92175
rect 279265 92147 279299 92175
rect 279327 92147 279361 92175
rect 279389 92147 279423 92175
rect 279451 92147 279499 92175
rect 279189 92113 279499 92147
rect 279189 92085 279237 92113
rect 279265 92085 279299 92113
rect 279327 92085 279361 92113
rect 279389 92085 279423 92113
rect 279451 92085 279499 92113
rect 279189 92051 279499 92085
rect 279189 92023 279237 92051
rect 279265 92023 279299 92051
rect 279327 92023 279361 92051
rect 279389 92023 279423 92051
rect 279451 92023 279499 92051
rect 279189 91989 279499 92023
rect 279189 91961 279237 91989
rect 279265 91961 279299 91989
rect 279327 91961 279361 91989
rect 279389 91961 279423 91989
rect 279451 91961 279499 91989
rect 265689 86147 265737 86175
rect 265765 86147 265799 86175
rect 265827 86147 265861 86175
rect 265889 86147 265923 86175
rect 265951 86147 265999 86175
rect 265689 86113 265999 86147
rect 265689 86085 265737 86113
rect 265765 86085 265799 86113
rect 265827 86085 265861 86113
rect 265889 86085 265923 86113
rect 265951 86085 265999 86113
rect 265689 86051 265999 86085
rect 265689 86023 265737 86051
rect 265765 86023 265799 86051
rect 265827 86023 265861 86051
rect 265889 86023 265923 86051
rect 265951 86023 265999 86051
rect 265689 85989 265999 86023
rect 265689 85961 265737 85989
rect 265765 85961 265799 85989
rect 265827 85961 265861 85989
rect 265889 85961 265923 85989
rect 265951 85961 265999 85989
rect 265689 77175 265999 85961
rect 277024 86175 277184 86192
rect 277024 86147 277059 86175
rect 277087 86147 277121 86175
rect 277149 86147 277184 86175
rect 277024 86113 277184 86147
rect 277024 86085 277059 86113
rect 277087 86085 277121 86113
rect 277149 86085 277184 86113
rect 277024 86051 277184 86085
rect 277024 86023 277059 86051
rect 277087 86023 277121 86051
rect 277149 86023 277184 86051
rect 277024 85989 277184 86023
rect 277024 85961 277059 85989
rect 277087 85961 277121 85989
rect 277149 85961 277184 85989
rect 277024 85944 277184 85961
rect 269344 83175 269504 83192
rect 269344 83147 269379 83175
rect 269407 83147 269441 83175
rect 269469 83147 269504 83175
rect 269344 83113 269504 83147
rect 269344 83085 269379 83113
rect 269407 83085 269441 83113
rect 269469 83085 269504 83113
rect 269344 83051 269504 83085
rect 269344 83023 269379 83051
rect 269407 83023 269441 83051
rect 269469 83023 269504 83051
rect 269344 82989 269504 83023
rect 269344 82961 269379 82989
rect 269407 82961 269441 82989
rect 269469 82961 269504 82989
rect 269344 82944 269504 82961
rect 279189 83175 279499 91961
rect 279189 83147 279237 83175
rect 279265 83147 279299 83175
rect 279327 83147 279361 83175
rect 279389 83147 279423 83175
rect 279451 83147 279499 83175
rect 279189 83113 279499 83147
rect 279189 83085 279237 83113
rect 279265 83085 279299 83113
rect 279327 83085 279361 83113
rect 279389 83085 279423 83113
rect 279451 83085 279499 83113
rect 279189 83051 279499 83085
rect 279189 83023 279237 83051
rect 279265 83023 279299 83051
rect 279327 83023 279361 83051
rect 279389 83023 279423 83051
rect 279451 83023 279499 83051
rect 279189 82989 279499 83023
rect 279189 82961 279237 82989
rect 279265 82961 279299 82989
rect 279327 82961 279361 82989
rect 279389 82961 279423 82989
rect 279451 82961 279499 82989
rect 265689 77147 265737 77175
rect 265765 77147 265799 77175
rect 265827 77147 265861 77175
rect 265889 77147 265923 77175
rect 265951 77147 265999 77175
rect 265689 77113 265999 77147
rect 265689 77085 265737 77113
rect 265765 77085 265799 77113
rect 265827 77085 265861 77113
rect 265889 77085 265923 77113
rect 265951 77085 265999 77113
rect 265689 77051 265999 77085
rect 265689 77023 265737 77051
rect 265765 77023 265799 77051
rect 265827 77023 265861 77051
rect 265889 77023 265923 77051
rect 265951 77023 265999 77051
rect 265689 76989 265999 77023
rect 265689 76961 265737 76989
rect 265765 76961 265799 76989
rect 265827 76961 265861 76989
rect 265889 76961 265923 76989
rect 265951 76961 265999 76989
rect 265689 68175 265999 76961
rect 277024 77175 277184 77192
rect 277024 77147 277059 77175
rect 277087 77147 277121 77175
rect 277149 77147 277184 77175
rect 277024 77113 277184 77147
rect 277024 77085 277059 77113
rect 277087 77085 277121 77113
rect 277149 77085 277184 77113
rect 277024 77051 277184 77085
rect 277024 77023 277059 77051
rect 277087 77023 277121 77051
rect 277149 77023 277184 77051
rect 277024 76989 277184 77023
rect 277024 76961 277059 76989
rect 277087 76961 277121 76989
rect 277149 76961 277184 76989
rect 277024 76944 277184 76961
rect 269344 74175 269504 74192
rect 269344 74147 269379 74175
rect 269407 74147 269441 74175
rect 269469 74147 269504 74175
rect 269344 74113 269504 74147
rect 269344 74085 269379 74113
rect 269407 74085 269441 74113
rect 269469 74085 269504 74113
rect 269344 74051 269504 74085
rect 269344 74023 269379 74051
rect 269407 74023 269441 74051
rect 269469 74023 269504 74051
rect 269344 73989 269504 74023
rect 269344 73961 269379 73989
rect 269407 73961 269441 73989
rect 269469 73961 269504 73989
rect 269344 73944 269504 73961
rect 279189 74175 279499 82961
rect 279189 74147 279237 74175
rect 279265 74147 279299 74175
rect 279327 74147 279361 74175
rect 279389 74147 279423 74175
rect 279451 74147 279499 74175
rect 279189 74113 279499 74147
rect 279189 74085 279237 74113
rect 279265 74085 279299 74113
rect 279327 74085 279361 74113
rect 279389 74085 279423 74113
rect 279451 74085 279499 74113
rect 279189 74051 279499 74085
rect 279189 74023 279237 74051
rect 279265 74023 279299 74051
rect 279327 74023 279361 74051
rect 279389 74023 279423 74051
rect 279451 74023 279499 74051
rect 279189 73989 279499 74023
rect 279189 73961 279237 73989
rect 279265 73961 279299 73989
rect 279327 73961 279361 73989
rect 279389 73961 279423 73989
rect 279451 73961 279499 73989
rect 265689 68147 265737 68175
rect 265765 68147 265799 68175
rect 265827 68147 265861 68175
rect 265889 68147 265923 68175
rect 265951 68147 265999 68175
rect 265689 68113 265999 68147
rect 265689 68085 265737 68113
rect 265765 68085 265799 68113
rect 265827 68085 265861 68113
rect 265889 68085 265923 68113
rect 265951 68085 265999 68113
rect 265689 68051 265999 68085
rect 265689 68023 265737 68051
rect 265765 68023 265799 68051
rect 265827 68023 265861 68051
rect 265889 68023 265923 68051
rect 265951 68023 265999 68051
rect 265689 67989 265999 68023
rect 265689 67961 265737 67989
rect 265765 67961 265799 67989
rect 265827 67961 265861 67989
rect 265889 67961 265923 67989
rect 265951 67961 265999 67989
rect 265689 59175 265999 67961
rect 277024 68175 277184 68192
rect 277024 68147 277059 68175
rect 277087 68147 277121 68175
rect 277149 68147 277184 68175
rect 277024 68113 277184 68147
rect 277024 68085 277059 68113
rect 277087 68085 277121 68113
rect 277149 68085 277184 68113
rect 277024 68051 277184 68085
rect 277024 68023 277059 68051
rect 277087 68023 277121 68051
rect 277149 68023 277184 68051
rect 277024 67989 277184 68023
rect 277024 67961 277059 67989
rect 277087 67961 277121 67989
rect 277149 67961 277184 67989
rect 277024 67944 277184 67961
rect 269344 65175 269504 65192
rect 269344 65147 269379 65175
rect 269407 65147 269441 65175
rect 269469 65147 269504 65175
rect 269344 65113 269504 65147
rect 269344 65085 269379 65113
rect 269407 65085 269441 65113
rect 269469 65085 269504 65113
rect 269344 65051 269504 65085
rect 269344 65023 269379 65051
rect 269407 65023 269441 65051
rect 269469 65023 269504 65051
rect 269344 64989 269504 65023
rect 269344 64961 269379 64989
rect 269407 64961 269441 64989
rect 269469 64961 269504 64989
rect 269344 64944 269504 64961
rect 279189 65175 279499 73961
rect 279189 65147 279237 65175
rect 279265 65147 279299 65175
rect 279327 65147 279361 65175
rect 279389 65147 279423 65175
rect 279451 65147 279499 65175
rect 279189 65113 279499 65147
rect 279189 65085 279237 65113
rect 279265 65085 279299 65113
rect 279327 65085 279361 65113
rect 279389 65085 279423 65113
rect 279451 65085 279499 65113
rect 279189 65051 279499 65085
rect 279189 65023 279237 65051
rect 279265 65023 279299 65051
rect 279327 65023 279361 65051
rect 279389 65023 279423 65051
rect 279451 65023 279499 65051
rect 279189 64989 279499 65023
rect 279189 64961 279237 64989
rect 279265 64961 279299 64989
rect 279327 64961 279361 64989
rect 279389 64961 279423 64989
rect 279451 64961 279499 64989
rect 265689 59147 265737 59175
rect 265765 59147 265799 59175
rect 265827 59147 265861 59175
rect 265889 59147 265923 59175
rect 265951 59147 265999 59175
rect 265689 59113 265999 59147
rect 265689 59085 265737 59113
rect 265765 59085 265799 59113
rect 265827 59085 265861 59113
rect 265889 59085 265923 59113
rect 265951 59085 265999 59113
rect 265689 59051 265999 59085
rect 265689 59023 265737 59051
rect 265765 59023 265799 59051
rect 265827 59023 265861 59051
rect 265889 59023 265923 59051
rect 265951 59023 265999 59051
rect 265689 58989 265999 59023
rect 265689 58961 265737 58989
rect 265765 58961 265799 58989
rect 265827 58961 265861 58989
rect 265889 58961 265923 58989
rect 265951 58961 265999 58989
rect 265689 50175 265999 58961
rect 277024 59175 277184 59192
rect 277024 59147 277059 59175
rect 277087 59147 277121 59175
rect 277149 59147 277184 59175
rect 277024 59113 277184 59147
rect 277024 59085 277059 59113
rect 277087 59085 277121 59113
rect 277149 59085 277184 59113
rect 277024 59051 277184 59085
rect 277024 59023 277059 59051
rect 277087 59023 277121 59051
rect 277149 59023 277184 59051
rect 277024 58989 277184 59023
rect 277024 58961 277059 58989
rect 277087 58961 277121 58989
rect 277149 58961 277184 58989
rect 277024 58944 277184 58961
rect 269344 56175 269504 56192
rect 269344 56147 269379 56175
rect 269407 56147 269441 56175
rect 269469 56147 269504 56175
rect 269344 56113 269504 56147
rect 269344 56085 269379 56113
rect 269407 56085 269441 56113
rect 269469 56085 269504 56113
rect 269344 56051 269504 56085
rect 269344 56023 269379 56051
rect 269407 56023 269441 56051
rect 269469 56023 269504 56051
rect 269344 55989 269504 56023
rect 269344 55961 269379 55989
rect 269407 55961 269441 55989
rect 269469 55961 269504 55989
rect 269344 55944 269504 55961
rect 279189 56175 279499 64961
rect 279189 56147 279237 56175
rect 279265 56147 279299 56175
rect 279327 56147 279361 56175
rect 279389 56147 279423 56175
rect 279451 56147 279499 56175
rect 279189 56113 279499 56147
rect 279189 56085 279237 56113
rect 279265 56085 279299 56113
rect 279327 56085 279361 56113
rect 279389 56085 279423 56113
rect 279451 56085 279499 56113
rect 279189 56051 279499 56085
rect 279189 56023 279237 56051
rect 279265 56023 279299 56051
rect 279327 56023 279361 56051
rect 279389 56023 279423 56051
rect 279451 56023 279499 56051
rect 279189 55989 279499 56023
rect 279189 55961 279237 55989
rect 279265 55961 279299 55989
rect 279327 55961 279361 55989
rect 279389 55961 279423 55989
rect 279451 55961 279499 55989
rect 265689 50147 265737 50175
rect 265765 50147 265799 50175
rect 265827 50147 265861 50175
rect 265889 50147 265923 50175
rect 265951 50147 265999 50175
rect 265689 50113 265999 50147
rect 265689 50085 265737 50113
rect 265765 50085 265799 50113
rect 265827 50085 265861 50113
rect 265889 50085 265923 50113
rect 265951 50085 265999 50113
rect 265689 50051 265999 50085
rect 265689 50023 265737 50051
rect 265765 50023 265799 50051
rect 265827 50023 265861 50051
rect 265889 50023 265923 50051
rect 265951 50023 265999 50051
rect 265689 49989 265999 50023
rect 265689 49961 265737 49989
rect 265765 49961 265799 49989
rect 265827 49961 265861 49989
rect 265889 49961 265923 49989
rect 265951 49961 265999 49989
rect 265689 41175 265999 49961
rect 277024 50175 277184 50192
rect 277024 50147 277059 50175
rect 277087 50147 277121 50175
rect 277149 50147 277184 50175
rect 277024 50113 277184 50147
rect 277024 50085 277059 50113
rect 277087 50085 277121 50113
rect 277149 50085 277184 50113
rect 277024 50051 277184 50085
rect 277024 50023 277059 50051
rect 277087 50023 277121 50051
rect 277149 50023 277184 50051
rect 277024 49989 277184 50023
rect 277024 49961 277059 49989
rect 277087 49961 277121 49989
rect 277149 49961 277184 49989
rect 277024 49944 277184 49961
rect 269344 47175 269504 47192
rect 269344 47147 269379 47175
rect 269407 47147 269441 47175
rect 269469 47147 269504 47175
rect 269344 47113 269504 47147
rect 269344 47085 269379 47113
rect 269407 47085 269441 47113
rect 269469 47085 269504 47113
rect 269344 47051 269504 47085
rect 269344 47023 269379 47051
rect 269407 47023 269441 47051
rect 269469 47023 269504 47051
rect 269344 46989 269504 47023
rect 269344 46961 269379 46989
rect 269407 46961 269441 46989
rect 269469 46961 269504 46989
rect 269344 46944 269504 46961
rect 279189 47175 279499 55961
rect 279189 47147 279237 47175
rect 279265 47147 279299 47175
rect 279327 47147 279361 47175
rect 279389 47147 279423 47175
rect 279451 47147 279499 47175
rect 279189 47113 279499 47147
rect 279189 47085 279237 47113
rect 279265 47085 279299 47113
rect 279327 47085 279361 47113
rect 279389 47085 279423 47113
rect 279451 47085 279499 47113
rect 279189 47051 279499 47085
rect 279189 47023 279237 47051
rect 279265 47023 279299 47051
rect 279327 47023 279361 47051
rect 279389 47023 279423 47051
rect 279451 47023 279499 47051
rect 279189 46989 279499 47023
rect 279189 46961 279237 46989
rect 279265 46961 279299 46989
rect 279327 46961 279361 46989
rect 279389 46961 279423 46989
rect 279451 46961 279499 46989
rect 265689 41147 265737 41175
rect 265765 41147 265799 41175
rect 265827 41147 265861 41175
rect 265889 41147 265923 41175
rect 265951 41147 265999 41175
rect 265689 41113 265999 41147
rect 265689 41085 265737 41113
rect 265765 41085 265799 41113
rect 265827 41085 265861 41113
rect 265889 41085 265923 41113
rect 265951 41085 265999 41113
rect 265689 41051 265999 41085
rect 265689 41023 265737 41051
rect 265765 41023 265799 41051
rect 265827 41023 265861 41051
rect 265889 41023 265923 41051
rect 265951 41023 265999 41051
rect 265689 40989 265999 41023
rect 265689 40961 265737 40989
rect 265765 40961 265799 40989
rect 265827 40961 265861 40989
rect 265889 40961 265923 40989
rect 265951 40961 265999 40989
rect 265689 32175 265999 40961
rect 277024 41175 277184 41192
rect 277024 41147 277059 41175
rect 277087 41147 277121 41175
rect 277149 41147 277184 41175
rect 277024 41113 277184 41147
rect 277024 41085 277059 41113
rect 277087 41085 277121 41113
rect 277149 41085 277184 41113
rect 277024 41051 277184 41085
rect 277024 41023 277059 41051
rect 277087 41023 277121 41051
rect 277149 41023 277184 41051
rect 277024 40989 277184 41023
rect 277024 40961 277059 40989
rect 277087 40961 277121 40989
rect 277149 40961 277184 40989
rect 277024 40944 277184 40961
rect 269344 38175 269504 38192
rect 269344 38147 269379 38175
rect 269407 38147 269441 38175
rect 269469 38147 269504 38175
rect 269344 38113 269504 38147
rect 269344 38085 269379 38113
rect 269407 38085 269441 38113
rect 269469 38085 269504 38113
rect 269344 38051 269504 38085
rect 269344 38023 269379 38051
rect 269407 38023 269441 38051
rect 269469 38023 269504 38051
rect 269344 37989 269504 38023
rect 269344 37961 269379 37989
rect 269407 37961 269441 37989
rect 269469 37961 269504 37989
rect 269344 37944 269504 37961
rect 279189 38175 279499 46961
rect 279189 38147 279237 38175
rect 279265 38147 279299 38175
rect 279327 38147 279361 38175
rect 279389 38147 279423 38175
rect 279451 38147 279499 38175
rect 279189 38113 279499 38147
rect 279189 38085 279237 38113
rect 279265 38085 279299 38113
rect 279327 38085 279361 38113
rect 279389 38085 279423 38113
rect 279451 38085 279499 38113
rect 279189 38051 279499 38085
rect 279189 38023 279237 38051
rect 279265 38023 279299 38051
rect 279327 38023 279361 38051
rect 279389 38023 279423 38051
rect 279451 38023 279499 38051
rect 279189 37989 279499 38023
rect 279189 37961 279237 37989
rect 279265 37961 279299 37989
rect 279327 37961 279361 37989
rect 279389 37961 279423 37989
rect 279451 37961 279499 37989
rect 265689 32147 265737 32175
rect 265765 32147 265799 32175
rect 265827 32147 265861 32175
rect 265889 32147 265923 32175
rect 265951 32147 265999 32175
rect 265689 32113 265999 32147
rect 265689 32085 265737 32113
rect 265765 32085 265799 32113
rect 265827 32085 265861 32113
rect 265889 32085 265923 32113
rect 265951 32085 265999 32113
rect 265689 32051 265999 32085
rect 265689 32023 265737 32051
rect 265765 32023 265799 32051
rect 265827 32023 265861 32051
rect 265889 32023 265923 32051
rect 265951 32023 265999 32051
rect 265689 31989 265999 32023
rect 265689 31961 265737 31989
rect 265765 31961 265799 31989
rect 265827 31961 265861 31989
rect 265889 31961 265923 31989
rect 265951 31961 265999 31989
rect 265689 23175 265999 31961
rect 277024 32175 277184 32192
rect 277024 32147 277059 32175
rect 277087 32147 277121 32175
rect 277149 32147 277184 32175
rect 277024 32113 277184 32147
rect 277024 32085 277059 32113
rect 277087 32085 277121 32113
rect 277149 32085 277184 32113
rect 277024 32051 277184 32085
rect 277024 32023 277059 32051
rect 277087 32023 277121 32051
rect 277149 32023 277184 32051
rect 277024 31989 277184 32023
rect 277024 31961 277059 31989
rect 277087 31961 277121 31989
rect 277149 31961 277184 31989
rect 277024 31944 277184 31961
rect 269344 29175 269504 29192
rect 269344 29147 269379 29175
rect 269407 29147 269441 29175
rect 269469 29147 269504 29175
rect 269344 29113 269504 29147
rect 269344 29085 269379 29113
rect 269407 29085 269441 29113
rect 269469 29085 269504 29113
rect 269344 29051 269504 29085
rect 269344 29023 269379 29051
rect 269407 29023 269441 29051
rect 269469 29023 269504 29051
rect 269344 28989 269504 29023
rect 269344 28961 269379 28989
rect 269407 28961 269441 28989
rect 269469 28961 269504 28989
rect 269344 28944 269504 28961
rect 279189 29175 279499 37961
rect 279189 29147 279237 29175
rect 279265 29147 279299 29175
rect 279327 29147 279361 29175
rect 279389 29147 279423 29175
rect 279451 29147 279499 29175
rect 279189 29113 279499 29147
rect 279189 29085 279237 29113
rect 279265 29085 279299 29113
rect 279327 29085 279361 29113
rect 279389 29085 279423 29113
rect 279451 29085 279499 29113
rect 279189 29051 279499 29085
rect 279189 29023 279237 29051
rect 279265 29023 279299 29051
rect 279327 29023 279361 29051
rect 279389 29023 279423 29051
rect 279451 29023 279499 29051
rect 279189 28989 279499 29023
rect 279189 28961 279237 28989
rect 279265 28961 279299 28989
rect 279327 28961 279361 28989
rect 279389 28961 279423 28989
rect 279451 28961 279499 28989
rect 265689 23147 265737 23175
rect 265765 23147 265799 23175
rect 265827 23147 265861 23175
rect 265889 23147 265923 23175
rect 265951 23147 265999 23175
rect 265689 23113 265999 23147
rect 265689 23085 265737 23113
rect 265765 23085 265799 23113
rect 265827 23085 265861 23113
rect 265889 23085 265923 23113
rect 265951 23085 265999 23113
rect 265689 23051 265999 23085
rect 265689 23023 265737 23051
rect 265765 23023 265799 23051
rect 265827 23023 265861 23051
rect 265889 23023 265923 23051
rect 265951 23023 265999 23051
rect 265689 22989 265999 23023
rect 265689 22961 265737 22989
rect 265765 22961 265799 22989
rect 265827 22961 265861 22989
rect 265889 22961 265923 22989
rect 265951 22961 265999 22989
rect 265689 14175 265999 22961
rect 277024 23175 277184 23192
rect 277024 23147 277059 23175
rect 277087 23147 277121 23175
rect 277149 23147 277184 23175
rect 277024 23113 277184 23147
rect 277024 23085 277059 23113
rect 277087 23085 277121 23113
rect 277149 23085 277184 23113
rect 277024 23051 277184 23085
rect 277024 23023 277059 23051
rect 277087 23023 277121 23051
rect 277149 23023 277184 23051
rect 277024 22989 277184 23023
rect 277024 22961 277059 22989
rect 277087 22961 277121 22989
rect 277149 22961 277184 22989
rect 277024 22944 277184 22961
rect 269344 20175 269504 20192
rect 269344 20147 269379 20175
rect 269407 20147 269441 20175
rect 269469 20147 269504 20175
rect 269344 20113 269504 20147
rect 269344 20085 269379 20113
rect 269407 20085 269441 20113
rect 269469 20085 269504 20113
rect 269344 20051 269504 20085
rect 269344 20023 269379 20051
rect 269407 20023 269441 20051
rect 269469 20023 269504 20051
rect 269344 19989 269504 20023
rect 269344 19961 269379 19989
rect 269407 19961 269441 19989
rect 269469 19961 269504 19989
rect 269344 19944 269504 19961
rect 279189 20175 279499 28961
rect 279189 20147 279237 20175
rect 279265 20147 279299 20175
rect 279327 20147 279361 20175
rect 279389 20147 279423 20175
rect 279451 20147 279499 20175
rect 279189 20113 279499 20147
rect 279189 20085 279237 20113
rect 279265 20085 279299 20113
rect 279327 20085 279361 20113
rect 279389 20085 279423 20113
rect 279451 20085 279499 20113
rect 279189 20051 279499 20085
rect 279189 20023 279237 20051
rect 279265 20023 279299 20051
rect 279327 20023 279361 20051
rect 279389 20023 279423 20051
rect 279451 20023 279499 20051
rect 279189 19989 279499 20023
rect 279189 19961 279237 19989
rect 279265 19961 279299 19989
rect 279327 19961 279361 19989
rect 279389 19961 279423 19989
rect 279451 19961 279499 19989
rect 265689 14147 265737 14175
rect 265765 14147 265799 14175
rect 265827 14147 265861 14175
rect 265889 14147 265923 14175
rect 265951 14147 265999 14175
rect 265689 14113 265999 14147
rect 265689 14085 265737 14113
rect 265765 14085 265799 14113
rect 265827 14085 265861 14113
rect 265889 14085 265923 14113
rect 265951 14085 265999 14113
rect 265689 14051 265999 14085
rect 265689 14023 265737 14051
rect 265765 14023 265799 14051
rect 265827 14023 265861 14051
rect 265889 14023 265923 14051
rect 265951 14023 265999 14051
rect 265689 13989 265999 14023
rect 265689 13961 265737 13989
rect 265765 13961 265799 13989
rect 265827 13961 265861 13989
rect 265889 13961 265923 13989
rect 265951 13961 265999 13989
rect 265689 5175 265999 13961
rect 277024 14175 277184 14192
rect 277024 14147 277059 14175
rect 277087 14147 277121 14175
rect 277149 14147 277184 14175
rect 277024 14113 277184 14147
rect 277024 14085 277059 14113
rect 277087 14085 277121 14113
rect 277149 14085 277184 14113
rect 277024 14051 277184 14085
rect 277024 14023 277059 14051
rect 277087 14023 277121 14051
rect 277149 14023 277184 14051
rect 277024 13989 277184 14023
rect 277024 13961 277059 13989
rect 277087 13961 277121 13989
rect 277149 13961 277184 13989
rect 277024 13944 277184 13961
rect 269344 11175 269504 11192
rect 269344 11147 269379 11175
rect 269407 11147 269441 11175
rect 269469 11147 269504 11175
rect 269344 11113 269504 11147
rect 269344 11085 269379 11113
rect 269407 11085 269441 11113
rect 269469 11085 269504 11113
rect 269344 11051 269504 11085
rect 269344 11023 269379 11051
rect 269407 11023 269441 11051
rect 269469 11023 269504 11051
rect 269344 10989 269504 11023
rect 269344 10961 269379 10989
rect 269407 10961 269441 10989
rect 269469 10961 269504 10989
rect 269344 10944 269504 10961
rect 279189 11175 279499 19961
rect 279189 11147 279237 11175
rect 279265 11147 279299 11175
rect 279327 11147 279361 11175
rect 279389 11147 279423 11175
rect 279451 11147 279499 11175
rect 279189 11113 279499 11147
rect 279189 11085 279237 11113
rect 279265 11085 279299 11113
rect 279327 11085 279361 11113
rect 279389 11085 279423 11113
rect 279451 11085 279499 11113
rect 279189 11051 279499 11085
rect 279189 11023 279237 11051
rect 279265 11023 279299 11051
rect 279327 11023 279361 11051
rect 279389 11023 279423 11051
rect 279451 11023 279499 11051
rect 279189 10989 279499 11023
rect 279189 10961 279237 10989
rect 279265 10961 279299 10989
rect 279327 10961 279361 10989
rect 279389 10961 279423 10989
rect 279451 10961 279499 10989
rect 265689 5147 265737 5175
rect 265765 5147 265799 5175
rect 265827 5147 265861 5175
rect 265889 5147 265923 5175
rect 265951 5147 265999 5175
rect 265689 5113 265999 5147
rect 265689 5085 265737 5113
rect 265765 5085 265799 5113
rect 265827 5085 265861 5113
rect 265889 5085 265923 5113
rect 265951 5085 265999 5113
rect 265689 5051 265999 5085
rect 265689 5023 265737 5051
rect 265765 5023 265799 5051
rect 265827 5023 265861 5051
rect 265889 5023 265923 5051
rect 265951 5023 265999 5051
rect 265689 4989 265999 5023
rect 265689 4961 265737 4989
rect 265765 4961 265799 4989
rect 265827 4961 265861 4989
rect 265889 4961 265923 4989
rect 265951 4961 265999 4989
rect 265689 -560 265999 4961
rect 277024 5175 277184 5192
rect 277024 5147 277059 5175
rect 277087 5147 277121 5175
rect 277149 5147 277184 5175
rect 277024 5113 277184 5147
rect 277024 5085 277059 5113
rect 277087 5085 277121 5113
rect 277149 5085 277184 5113
rect 277024 5051 277184 5085
rect 277024 5023 277059 5051
rect 277087 5023 277121 5051
rect 277149 5023 277184 5051
rect 277024 4989 277184 5023
rect 277024 4961 277059 4989
rect 277087 4961 277121 4989
rect 277149 4961 277184 4989
rect 277024 4944 277184 4961
rect 265689 -588 265737 -560
rect 265765 -588 265799 -560
rect 265827 -588 265861 -560
rect 265889 -588 265923 -560
rect 265951 -588 265999 -560
rect 265689 -622 265999 -588
rect 265689 -650 265737 -622
rect 265765 -650 265799 -622
rect 265827 -650 265861 -622
rect 265889 -650 265923 -622
rect 265951 -650 265999 -622
rect 265689 -684 265999 -650
rect 265689 -712 265737 -684
rect 265765 -712 265799 -684
rect 265827 -712 265861 -684
rect 265889 -712 265923 -684
rect 265951 -712 265999 -684
rect 265689 -746 265999 -712
rect 265689 -774 265737 -746
rect 265765 -774 265799 -746
rect 265827 -774 265861 -746
rect 265889 -774 265923 -746
rect 265951 -774 265999 -746
rect 265689 -822 265999 -774
rect 279189 2175 279499 10961
rect 279189 2147 279237 2175
rect 279265 2147 279299 2175
rect 279327 2147 279361 2175
rect 279389 2147 279423 2175
rect 279451 2147 279499 2175
rect 279189 2113 279499 2147
rect 279189 2085 279237 2113
rect 279265 2085 279299 2113
rect 279327 2085 279361 2113
rect 279389 2085 279423 2113
rect 279451 2085 279499 2113
rect 279189 2051 279499 2085
rect 279189 2023 279237 2051
rect 279265 2023 279299 2051
rect 279327 2023 279361 2051
rect 279389 2023 279423 2051
rect 279451 2023 279499 2051
rect 279189 1989 279499 2023
rect 279189 1961 279237 1989
rect 279265 1961 279299 1989
rect 279327 1961 279361 1989
rect 279389 1961 279423 1989
rect 279451 1961 279499 1989
rect 279189 -80 279499 1961
rect 279189 -108 279237 -80
rect 279265 -108 279299 -80
rect 279327 -108 279361 -80
rect 279389 -108 279423 -80
rect 279451 -108 279499 -80
rect 279189 -142 279499 -108
rect 279189 -170 279237 -142
rect 279265 -170 279299 -142
rect 279327 -170 279361 -142
rect 279389 -170 279423 -142
rect 279451 -170 279499 -142
rect 279189 -204 279499 -170
rect 279189 -232 279237 -204
rect 279265 -232 279299 -204
rect 279327 -232 279361 -204
rect 279389 -232 279423 -204
rect 279451 -232 279499 -204
rect 279189 -266 279499 -232
rect 279189 -294 279237 -266
rect 279265 -294 279299 -266
rect 279327 -294 279361 -266
rect 279389 -294 279423 -266
rect 279451 -294 279499 -266
rect 279189 -822 279499 -294
rect 281049 299086 281359 299134
rect 281049 299058 281097 299086
rect 281125 299058 281159 299086
rect 281187 299058 281221 299086
rect 281249 299058 281283 299086
rect 281311 299058 281359 299086
rect 281049 299024 281359 299058
rect 281049 298996 281097 299024
rect 281125 298996 281159 299024
rect 281187 298996 281221 299024
rect 281249 298996 281283 299024
rect 281311 298996 281359 299024
rect 281049 298962 281359 298996
rect 281049 298934 281097 298962
rect 281125 298934 281159 298962
rect 281187 298934 281221 298962
rect 281249 298934 281283 298962
rect 281311 298934 281359 298962
rect 281049 298900 281359 298934
rect 281049 298872 281097 298900
rect 281125 298872 281159 298900
rect 281187 298872 281221 298900
rect 281249 298872 281283 298900
rect 281311 298872 281359 298900
rect 281049 293175 281359 298872
rect 281049 293147 281097 293175
rect 281125 293147 281159 293175
rect 281187 293147 281221 293175
rect 281249 293147 281283 293175
rect 281311 293147 281359 293175
rect 281049 293113 281359 293147
rect 281049 293085 281097 293113
rect 281125 293085 281159 293113
rect 281187 293085 281221 293113
rect 281249 293085 281283 293113
rect 281311 293085 281359 293113
rect 281049 293051 281359 293085
rect 281049 293023 281097 293051
rect 281125 293023 281159 293051
rect 281187 293023 281221 293051
rect 281249 293023 281283 293051
rect 281311 293023 281359 293051
rect 281049 292989 281359 293023
rect 281049 292961 281097 292989
rect 281125 292961 281159 292989
rect 281187 292961 281221 292989
rect 281249 292961 281283 292989
rect 281311 292961 281359 292989
rect 281049 284175 281359 292961
rect 281049 284147 281097 284175
rect 281125 284147 281159 284175
rect 281187 284147 281221 284175
rect 281249 284147 281283 284175
rect 281311 284147 281359 284175
rect 281049 284113 281359 284147
rect 281049 284085 281097 284113
rect 281125 284085 281159 284113
rect 281187 284085 281221 284113
rect 281249 284085 281283 284113
rect 281311 284085 281359 284113
rect 281049 284051 281359 284085
rect 281049 284023 281097 284051
rect 281125 284023 281159 284051
rect 281187 284023 281221 284051
rect 281249 284023 281283 284051
rect 281311 284023 281359 284051
rect 281049 283989 281359 284023
rect 281049 283961 281097 283989
rect 281125 283961 281159 283989
rect 281187 283961 281221 283989
rect 281249 283961 281283 283989
rect 281311 283961 281359 283989
rect 281049 275175 281359 283961
rect 281049 275147 281097 275175
rect 281125 275147 281159 275175
rect 281187 275147 281221 275175
rect 281249 275147 281283 275175
rect 281311 275147 281359 275175
rect 281049 275113 281359 275147
rect 281049 275085 281097 275113
rect 281125 275085 281159 275113
rect 281187 275085 281221 275113
rect 281249 275085 281283 275113
rect 281311 275085 281359 275113
rect 281049 275051 281359 275085
rect 281049 275023 281097 275051
rect 281125 275023 281159 275051
rect 281187 275023 281221 275051
rect 281249 275023 281283 275051
rect 281311 275023 281359 275051
rect 281049 274989 281359 275023
rect 281049 274961 281097 274989
rect 281125 274961 281159 274989
rect 281187 274961 281221 274989
rect 281249 274961 281283 274989
rect 281311 274961 281359 274989
rect 281049 266175 281359 274961
rect 281049 266147 281097 266175
rect 281125 266147 281159 266175
rect 281187 266147 281221 266175
rect 281249 266147 281283 266175
rect 281311 266147 281359 266175
rect 281049 266113 281359 266147
rect 281049 266085 281097 266113
rect 281125 266085 281159 266113
rect 281187 266085 281221 266113
rect 281249 266085 281283 266113
rect 281311 266085 281359 266113
rect 281049 266051 281359 266085
rect 281049 266023 281097 266051
rect 281125 266023 281159 266051
rect 281187 266023 281221 266051
rect 281249 266023 281283 266051
rect 281311 266023 281359 266051
rect 281049 265989 281359 266023
rect 281049 265961 281097 265989
rect 281125 265961 281159 265989
rect 281187 265961 281221 265989
rect 281249 265961 281283 265989
rect 281311 265961 281359 265989
rect 281049 257175 281359 265961
rect 281049 257147 281097 257175
rect 281125 257147 281159 257175
rect 281187 257147 281221 257175
rect 281249 257147 281283 257175
rect 281311 257147 281359 257175
rect 281049 257113 281359 257147
rect 281049 257085 281097 257113
rect 281125 257085 281159 257113
rect 281187 257085 281221 257113
rect 281249 257085 281283 257113
rect 281311 257085 281359 257113
rect 281049 257051 281359 257085
rect 281049 257023 281097 257051
rect 281125 257023 281159 257051
rect 281187 257023 281221 257051
rect 281249 257023 281283 257051
rect 281311 257023 281359 257051
rect 281049 256989 281359 257023
rect 281049 256961 281097 256989
rect 281125 256961 281159 256989
rect 281187 256961 281221 256989
rect 281249 256961 281283 256989
rect 281311 256961 281359 256989
rect 281049 248175 281359 256961
rect 281049 248147 281097 248175
rect 281125 248147 281159 248175
rect 281187 248147 281221 248175
rect 281249 248147 281283 248175
rect 281311 248147 281359 248175
rect 281049 248113 281359 248147
rect 281049 248085 281097 248113
rect 281125 248085 281159 248113
rect 281187 248085 281221 248113
rect 281249 248085 281283 248113
rect 281311 248085 281359 248113
rect 281049 248051 281359 248085
rect 281049 248023 281097 248051
rect 281125 248023 281159 248051
rect 281187 248023 281221 248051
rect 281249 248023 281283 248051
rect 281311 248023 281359 248051
rect 281049 247989 281359 248023
rect 281049 247961 281097 247989
rect 281125 247961 281159 247989
rect 281187 247961 281221 247989
rect 281249 247961 281283 247989
rect 281311 247961 281359 247989
rect 281049 239175 281359 247961
rect 281049 239147 281097 239175
rect 281125 239147 281159 239175
rect 281187 239147 281221 239175
rect 281249 239147 281283 239175
rect 281311 239147 281359 239175
rect 281049 239113 281359 239147
rect 281049 239085 281097 239113
rect 281125 239085 281159 239113
rect 281187 239085 281221 239113
rect 281249 239085 281283 239113
rect 281311 239085 281359 239113
rect 281049 239051 281359 239085
rect 281049 239023 281097 239051
rect 281125 239023 281159 239051
rect 281187 239023 281221 239051
rect 281249 239023 281283 239051
rect 281311 239023 281359 239051
rect 281049 238989 281359 239023
rect 281049 238961 281097 238989
rect 281125 238961 281159 238989
rect 281187 238961 281221 238989
rect 281249 238961 281283 238989
rect 281311 238961 281359 238989
rect 281049 230175 281359 238961
rect 281049 230147 281097 230175
rect 281125 230147 281159 230175
rect 281187 230147 281221 230175
rect 281249 230147 281283 230175
rect 281311 230147 281359 230175
rect 281049 230113 281359 230147
rect 281049 230085 281097 230113
rect 281125 230085 281159 230113
rect 281187 230085 281221 230113
rect 281249 230085 281283 230113
rect 281311 230085 281359 230113
rect 281049 230051 281359 230085
rect 281049 230023 281097 230051
rect 281125 230023 281159 230051
rect 281187 230023 281221 230051
rect 281249 230023 281283 230051
rect 281311 230023 281359 230051
rect 281049 229989 281359 230023
rect 281049 229961 281097 229989
rect 281125 229961 281159 229989
rect 281187 229961 281221 229989
rect 281249 229961 281283 229989
rect 281311 229961 281359 229989
rect 281049 221175 281359 229961
rect 281049 221147 281097 221175
rect 281125 221147 281159 221175
rect 281187 221147 281221 221175
rect 281249 221147 281283 221175
rect 281311 221147 281359 221175
rect 281049 221113 281359 221147
rect 281049 221085 281097 221113
rect 281125 221085 281159 221113
rect 281187 221085 281221 221113
rect 281249 221085 281283 221113
rect 281311 221085 281359 221113
rect 281049 221051 281359 221085
rect 281049 221023 281097 221051
rect 281125 221023 281159 221051
rect 281187 221023 281221 221051
rect 281249 221023 281283 221051
rect 281311 221023 281359 221051
rect 281049 220989 281359 221023
rect 281049 220961 281097 220989
rect 281125 220961 281159 220989
rect 281187 220961 281221 220989
rect 281249 220961 281283 220989
rect 281311 220961 281359 220989
rect 281049 212175 281359 220961
rect 281049 212147 281097 212175
rect 281125 212147 281159 212175
rect 281187 212147 281221 212175
rect 281249 212147 281283 212175
rect 281311 212147 281359 212175
rect 281049 212113 281359 212147
rect 281049 212085 281097 212113
rect 281125 212085 281159 212113
rect 281187 212085 281221 212113
rect 281249 212085 281283 212113
rect 281311 212085 281359 212113
rect 281049 212051 281359 212085
rect 281049 212023 281097 212051
rect 281125 212023 281159 212051
rect 281187 212023 281221 212051
rect 281249 212023 281283 212051
rect 281311 212023 281359 212051
rect 281049 211989 281359 212023
rect 281049 211961 281097 211989
rect 281125 211961 281159 211989
rect 281187 211961 281221 211989
rect 281249 211961 281283 211989
rect 281311 211961 281359 211989
rect 281049 203175 281359 211961
rect 281049 203147 281097 203175
rect 281125 203147 281159 203175
rect 281187 203147 281221 203175
rect 281249 203147 281283 203175
rect 281311 203147 281359 203175
rect 281049 203113 281359 203147
rect 281049 203085 281097 203113
rect 281125 203085 281159 203113
rect 281187 203085 281221 203113
rect 281249 203085 281283 203113
rect 281311 203085 281359 203113
rect 281049 203051 281359 203085
rect 281049 203023 281097 203051
rect 281125 203023 281159 203051
rect 281187 203023 281221 203051
rect 281249 203023 281283 203051
rect 281311 203023 281359 203051
rect 281049 202989 281359 203023
rect 281049 202961 281097 202989
rect 281125 202961 281159 202989
rect 281187 202961 281221 202989
rect 281249 202961 281283 202989
rect 281311 202961 281359 202989
rect 281049 194175 281359 202961
rect 281049 194147 281097 194175
rect 281125 194147 281159 194175
rect 281187 194147 281221 194175
rect 281249 194147 281283 194175
rect 281311 194147 281359 194175
rect 281049 194113 281359 194147
rect 281049 194085 281097 194113
rect 281125 194085 281159 194113
rect 281187 194085 281221 194113
rect 281249 194085 281283 194113
rect 281311 194085 281359 194113
rect 281049 194051 281359 194085
rect 281049 194023 281097 194051
rect 281125 194023 281159 194051
rect 281187 194023 281221 194051
rect 281249 194023 281283 194051
rect 281311 194023 281359 194051
rect 281049 193989 281359 194023
rect 281049 193961 281097 193989
rect 281125 193961 281159 193989
rect 281187 193961 281221 193989
rect 281249 193961 281283 193989
rect 281311 193961 281359 193989
rect 281049 185175 281359 193961
rect 281049 185147 281097 185175
rect 281125 185147 281159 185175
rect 281187 185147 281221 185175
rect 281249 185147 281283 185175
rect 281311 185147 281359 185175
rect 281049 185113 281359 185147
rect 281049 185085 281097 185113
rect 281125 185085 281159 185113
rect 281187 185085 281221 185113
rect 281249 185085 281283 185113
rect 281311 185085 281359 185113
rect 281049 185051 281359 185085
rect 281049 185023 281097 185051
rect 281125 185023 281159 185051
rect 281187 185023 281221 185051
rect 281249 185023 281283 185051
rect 281311 185023 281359 185051
rect 281049 184989 281359 185023
rect 281049 184961 281097 184989
rect 281125 184961 281159 184989
rect 281187 184961 281221 184989
rect 281249 184961 281283 184989
rect 281311 184961 281359 184989
rect 281049 176175 281359 184961
rect 281049 176147 281097 176175
rect 281125 176147 281159 176175
rect 281187 176147 281221 176175
rect 281249 176147 281283 176175
rect 281311 176147 281359 176175
rect 281049 176113 281359 176147
rect 281049 176085 281097 176113
rect 281125 176085 281159 176113
rect 281187 176085 281221 176113
rect 281249 176085 281283 176113
rect 281311 176085 281359 176113
rect 281049 176051 281359 176085
rect 281049 176023 281097 176051
rect 281125 176023 281159 176051
rect 281187 176023 281221 176051
rect 281249 176023 281283 176051
rect 281311 176023 281359 176051
rect 281049 175989 281359 176023
rect 281049 175961 281097 175989
rect 281125 175961 281159 175989
rect 281187 175961 281221 175989
rect 281249 175961 281283 175989
rect 281311 175961 281359 175989
rect 281049 167175 281359 175961
rect 294549 298606 294859 299134
rect 294549 298578 294597 298606
rect 294625 298578 294659 298606
rect 294687 298578 294721 298606
rect 294749 298578 294783 298606
rect 294811 298578 294859 298606
rect 294549 298544 294859 298578
rect 294549 298516 294597 298544
rect 294625 298516 294659 298544
rect 294687 298516 294721 298544
rect 294749 298516 294783 298544
rect 294811 298516 294859 298544
rect 294549 298482 294859 298516
rect 294549 298454 294597 298482
rect 294625 298454 294659 298482
rect 294687 298454 294721 298482
rect 294749 298454 294783 298482
rect 294811 298454 294859 298482
rect 294549 298420 294859 298454
rect 294549 298392 294597 298420
rect 294625 298392 294659 298420
rect 294687 298392 294721 298420
rect 294749 298392 294783 298420
rect 294811 298392 294859 298420
rect 294549 290175 294859 298392
rect 294549 290147 294597 290175
rect 294625 290147 294659 290175
rect 294687 290147 294721 290175
rect 294749 290147 294783 290175
rect 294811 290147 294859 290175
rect 294549 290113 294859 290147
rect 294549 290085 294597 290113
rect 294625 290085 294659 290113
rect 294687 290085 294721 290113
rect 294749 290085 294783 290113
rect 294811 290085 294859 290113
rect 294549 290051 294859 290085
rect 294549 290023 294597 290051
rect 294625 290023 294659 290051
rect 294687 290023 294721 290051
rect 294749 290023 294783 290051
rect 294811 290023 294859 290051
rect 294549 289989 294859 290023
rect 294549 289961 294597 289989
rect 294625 289961 294659 289989
rect 294687 289961 294721 289989
rect 294749 289961 294783 289989
rect 294811 289961 294859 289989
rect 294549 281175 294859 289961
rect 294549 281147 294597 281175
rect 294625 281147 294659 281175
rect 294687 281147 294721 281175
rect 294749 281147 294783 281175
rect 294811 281147 294859 281175
rect 294549 281113 294859 281147
rect 294549 281085 294597 281113
rect 294625 281085 294659 281113
rect 294687 281085 294721 281113
rect 294749 281085 294783 281113
rect 294811 281085 294859 281113
rect 294549 281051 294859 281085
rect 294549 281023 294597 281051
rect 294625 281023 294659 281051
rect 294687 281023 294721 281051
rect 294749 281023 294783 281051
rect 294811 281023 294859 281051
rect 294549 280989 294859 281023
rect 294549 280961 294597 280989
rect 294625 280961 294659 280989
rect 294687 280961 294721 280989
rect 294749 280961 294783 280989
rect 294811 280961 294859 280989
rect 294549 272175 294859 280961
rect 294549 272147 294597 272175
rect 294625 272147 294659 272175
rect 294687 272147 294721 272175
rect 294749 272147 294783 272175
rect 294811 272147 294859 272175
rect 294549 272113 294859 272147
rect 294549 272085 294597 272113
rect 294625 272085 294659 272113
rect 294687 272085 294721 272113
rect 294749 272085 294783 272113
rect 294811 272085 294859 272113
rect 294549 272051 294859 272085
rect 294549 272023 294597 272051
rect 294625 272023 294659 272051
rect 294687 272023 294721 272051
rect 294749 272023 294783 272051
rect 294811 272023 294859 272051
rect 294549 271989 294859 272023
rect 294549 271961 294597 271989
rect 294625 271961 294659 271989
rect 294687 271961 294721 271989
rect 294749 271961 294783 271989
rect 294811 271961 294859 271989
rect 294549 263175 294859 271961
rect 294549 263147 294597 263175
rect 294625 263147 294659 263175
rect 294687 263147 294721 263175
rect 294749 263147 294783 263175
rect 294811 263147 294859 263175
rect 294549 263113 294859 263147
rect 294549 263085 294597 263113
rect 294625 263085 294659 263113
rect 294687 263085 294721 263113
rect 294749 263085 294783 263113
rect 294811 263085 294859 263113
rect 294549 263051 294859 263085
rect 294549 263023 294597 263051
rect 294625 263023 294659 263051
rect 294687 263023 294721 263051
rect 294749 263023 294783 263051
rect 294811 263023 294859 263051
rect 294549 262989 294859 263023
rect 294549 262961 294597 262989
rect 294625 262961 294659 262989
rect 294687 262961 294721 262989
rect 294749 262961 294783 262989
rect 294811 262961 294859 262989
rect 294549 254175 294859 262961
rect 294549 254147 294597 254175
rect 294625 254147 294659 254175
rect 294687 254147 294721 254175
rect 294749 254147 294783 254175
rect 294811 254147 294859 254175
rect 294549 254113 294859 254147
rect 294549 254085 294597 254113
rect 294625 254085 294659 254113
rect 294687 254085 294721 254113
rect 294749 254085 294783 254113
rect 294811 254085 294859 254113
rect 294549 254051 294859 254085
rect 294549 254023 294597 254051
rect 294625 254023 294659 254051
rect 294687 254023 294721 254051
rect 294749 254023 294783 254051
rect 294811 254023 294859 254051
rect 294549 253989 294859 254023
rect 294549 253961 294597 253989
rect 294625 253961 294659 253989
rect 294687 253961 294721 253989
rect 294749 253961 294783 253989
rect 294811 253961 294859 253989
rect 294549 245175 294859 253961
rect 294549 245147 294597 245175
rect 294625 245147 294659 245175
rect 294687 245147 294721 245175
rect 294749 245147 294783 245175
rect 294811 245147 294859 245175
rect 294549 245113 294859 245147
rect 294549 245085 294597 245113
rect 294625 245085 294659 245113
rect 294687 245085 294721 245113
rect 294749 245085 294783 245113
rect 294811 245085 294859 245113
rect 294549 245051 294859 245085
rect 294549 245023 294597 245051
rect 294625 245023 294659 245051
rect 294687 245023 294721 245051
rect 294749 245023 294783 245051
rect 294811 245023 294859 245051
rect 294549 244989 294859 245023
rect 294549 244961 294597 244989
rect 294625 244961 294659 244989
rect 294687 244961 294721 244989
rect 294749 244961 294783 244989
rect 294811 244961 294859 244989
rect 294549 236175 294859 244961
rect 294549 236147 294597 236175
rect 294625 236147 294659 236175
rect 294687 236147 294721 236175
rect 294749 236147 294783 236175
rect 294811 236147 294859 236175
rect 294549 236113 294859 236147
rect 294549 236085 294597 236113
rect 294625 236085 294659 236113
rect 294687 236085 294721 236113
rect 294749 236085 294783 236113
rect 294811 236085 294859 236113
rect 294549 236051 294859 236085
rect 294549 236023 294597 236051
rect 294625 236023 294659 236051
rect 294687 236023 294721 236051
rect 294749 236023 294783 236051
rect 294811 236023 294859 236051
rect 294549 235989 294859 236023
rect 294549 235961 294597 235989
rect 294625 235961 294659 235989
rect 294687 235961 294721 235989
rect 294749 235961 294783 235989
rect 294811 235961 294859 235989
rect 294549 227175 294859 235961
rect 294549 227147 294597 227175
rect 294625 227147 294659 227175
rect 294687 227147 294721 227175
rect 294749 227147 294783 227175
rect 294811 227147 294859 227175
rect 294549 227113 294859 227147
rect 294549 227085 294597 227113
rect 294625 227085 294659 227113
rect 294687 227085 294721 227113
rect 294749 227085 294783 227113
rect 294811 227085 294859 227113
rect 294549 227051 294859 227085
rect 294549 227023 294597 227051
rect 294625 227023 294659 227051
rect 294687 227023 294721 227051
rect 294749 227023 294783 227051
rect 294811 227023 294859 227051
rect 294549 226989 294859 227023
rect 294549 226961 294597 226989
rect 294625 226961 294659 226989
rect 294687 226961 294721 226989
rect 294749 226961 294783 226989
rect 294811 226961 294859 226989
rect 294549 218175 294859 226961
rect 294549 218147 294597 218175
rect 294625 218147 294659 218175
rect 294687 218147 294721 218175
rect 294749 218147 294783 218175
rect 294811 218147 294859 218175
rect 294549 218113 294859 218147
rect 294549 218085 294597 218113
rect 294625 218085 294659 218113
rect 294687 218085 294721 218113
rect 294749 218085 294783 218113
rect 294811 218085 294859 218113
rect 294549 218051 294859 218085
rect 294549 218023 294597 218051
rect 294625 218023 294659 218051
rect 294687 218023 294721 218051
rect 294749 218023 294783 218051
rect 294811 218023 294859 218051
rect 294549 217989 294859 218023
rect 294549 217961 294597 217989
rect 294625 217961 294659 217989
rect 294687 217961 294721 217989
rect 294749 217961 294783 217989
rect 294811 217961 294859 217989
rect 294549 209175 294859 217961
rect 294549 209147 294597 209175
rect 294625 209147 294659 209175
rect 294687 209147 294721 209175
rect 294749 209147 294783 209175
rect 294811 209147 294859 209175
rect 294549 209113 294859 209147
rect 294549 209085 294597 209113
rect 294625 209085 294659 209113
rect 294687 209085 294721 209113
rect 294749 209085 294783 209113
rect 294811 209085 294859 209113
rect 294549 209051 294859 209085
rect 294549 209023 294597 209051
rect 294625 209023 294659 209051
rect 294687 209023 294721 209051
rect 294749 209023 294783 209051
rect 294811 209023 294859 209051
rect 294549 208989 294859 209023
rect 294549 208961 294597 208989
rect 294625 208961 294659 208989
rect 294687 208961 294721 208989
rect 294749 208961 294783 208989
rect 294811 208961 294859 208989
rect 294549 200175 294859 208961
rect 294549 200147 294597 200175
rect 294625 200147 294659 200175
rect 294687 200147 294721 200175
rect 294749 200147 294783 200175
rect 294811 200147 294859 200175
rect 294549 200113 294859 200147
rect 294549 200085 294597 200113
rect 294625 200085 294659 200113
rect 294687 200085 294721 200113
rect 294749 200085 294783 200113
rect 294811 200085 294859 200113
rect 294549 200051 294859 200085
rect 294549 200023 294597 200051
rect 294625 200023 294659 200051
rect 294687 200023 294721 200051
rect 294749 200023 294783 200051
rect 294811 200023 294859 200051
rect 294549 199989 294859 200023
rect 294549 199961 294597 199989
rect 294625 199961 294659 199989
rect 294687 199961 294721 199989
rect 294749 199961 294783 199989
rect 294811 199961 294859 199989
rect 294549 191175 294859 199961
rect 294549 191147 294597 191175
rect 294625 191147 294659 191175
rect 294687 191147 294721 191175
rect 294749 191147 294783 191175
rect 294811 191147 294859 191175
rect 294549 191113 294859 191147
rect 294549 191085 294597 191113
rect 294625 191085 294659 191113
rect 294687 191085 294721 191113
rect 294749 191085 294783 191113
rect 294811 191085 294859 191113
rect 294549 191051 294859 191085
rect 294549 191023 294597 191051
rect 294625 191023 294659 191051
rect 294687 191023 294721 191051
rect 294749 191023 294783 191051
rect 294811 191023 294859 191051
rect 294549 190989 294859 191023
rect 294549 190961 294597 190989
rect 294625 190961 294659 190989
rect 294687 190961 294721 190989
rect 294749 190961 294783 190989
rect 294811 190961 294859 190989
rect 294549 182175 294859 190961
rect 294549 182147 294597 182175
rect 294625 182147 294659 182175
rect 294687 182147 294721 182175
rect 294749 182147 294783 182175
rect 294811 182147 294859 182175
rect 294549 182113 294859 182147
rect 294549 182085 294597 182113
rect 294625 182085 294659 182113
rect 294687 182085 294721 182113
rect 294749 182085 294783 182113
rect 294811 182085 294859 182113
rect 294549 182051 294859 182085
rect 294549 182023 294597 182051
rect 294625 182023 294659 182051
rect 294687 182023 294721 182051
rect 294749 182023 294783 182051
rect 294811 182023 294859 182051
rect 294549 181989 294859 182023
rect 294549 181961 294597 181989
rect 294625 181961 294659 181989
rect 294687 181961 294721 181989
rect 294749 181961 294783 181989
rect 294811 181961 294859 181989
rect 287686 173250 287714 173255
rect 284704 173175 284864 173192
rect 284704 173147 284739 173175
rect 284767 173147 284801 173175
rect 284829 173147 284864 173175
rect 284704 173113 284864 173147
rect 284704 173085 284739 173113
rect 284767 173085 284801 173113
rect 284829 173085 284864 173113
rect 284704 173051 284864 173085
rect 284704 173023 284739 173051
rect 284767 173023 284801 173051
rect 284829 173023 284864 173051
rect 284704 172989 284864 173023
rect 284704 172961 284739 172989
rect 284767 172961 284801 172989
rect 284829 172961 284864 172989
rect 284704 172944 284864 172961
rect 281049 167147 281097 167175
rect 281125 167147 281159 167175
rect 281187 167147 281221 167175
rect 281249 167147 281283 167175
rect 281311 167147 281359 167175
rect 281049 167113 281359 167147
rect 281049 167085 281097 167113
rect 281125 167085 281159 167113
rect 281187 167085 281221 167113
rect 281249 167085 281283 167113
rect 281311 167085 281359 167113
rect 281049 167051 281359 167085
rect 281049 167023 281097 167051
rect 281125 167023 281159 167051
rect 281187 167023 281221 167051
rect 281249 167023 281283 167051
rect 281311 167023 281359 167051
rect 281049 166989 281359 167023
rect 281049 166961 281097 166989
rect 281125 166961 281159 166989
rect 281187 166961 281221 166989
rect 281249 166961 281283 166989
rect 281311 166961 281359 166989
rect 281049 158175 281359 166961
rect 284704 164175 284864 164192
rect 284704 164147 284739 164175
rect 284767 164147 284801 164175
rect 284829 164147 284864 164175
rect 284704 164113 284864 164147
rect 284704 164085 284739 164113
rect 284767 164085 284801 164113
rect 284829 164085 284864 164113
rect 284704 164051 284864 164085
rect 284704 164023 284739 164051
rect 284767 164023 284801 164051
rect 284829 164023 284864 164051
rect 284704 163989 284864 164023
rect 284704 163961 284739 163989
rect 284767 163961 284801 163989
rect 284829 163961 284864 163989
rect 284704 163944 284864 163961
rect 281049 158147 281097 158175
rect 281125 158147 281159 158175
rect 281187 158147 281221 158175
rect 281249 158147 281283 158175
rect 281311 158147 281359 158175
rect 281049 158113 281359 158147
rect 281049 158085 281097 158113
rect 281125 158085 281159 158113
rect 281187 158085 281221 158113
rect 281249 158085 281283 158113
rect 281311 158085 281359 158113
rect 281049 158051 281359 158085
rect 281049 158023 281097 158051
rect 281125 158023 281159 158051
rect 281187 158023 281221 158051
rect 281249 158023 281283 158051
rect 281311 158023 281359 158051
rect 281049 157989 281359 158023
rect 281049 157961 281097 157989
rect 281125 157961 281159 157989
rect 281187 157961 281221 157989
rect 281249 157961 281283 157989
rect 281311 157961 281359 157989
rect 281049 149175 281359 157961
rect 287686 155554 287714 173222
rect 294549 173175 294859 181961
rect 294549 173147 294597 173175
rect 294625 173147 294659 173175
rect 294687 173147 294721 173175
rect 294749 173147 294783 173175
rect 294811 173147 294859 173175
rect 294549 173113 294859 173147
rect 294549 173085 294597 173113
rect 294625 173085 294659 173113
rect 294687 173085 294721 173113
rect 294749 173085 294783 173113
rect 294811 173085 294859 173113
rect 294549 173051 294859 173085
rect 294549 173023 294597 173051
rect 294625 173023 294659 173051
rect 294687 173023 294721 173051
rect 294749 173023 294783 173051
rect 294811 173023 294859 173051
rect 294549 172989 294859 173023
rect 294549 172961 294597 172989
rect 294625 172961 294659 172989
rect 294687 172961 294721 172989
rect 294749 172961 294783 172989
rect 294811 172961 294859 172989
rect 287686 155521 287714 155526
rect 287742 165970 287770 165975
rect 284704 155175 284864 155192
rect 284704 155147 284739 155175
rect 284767 155147 284801 155175
rect 284829 155147 284864 155175
rect 284704 155113 284864 155147
rect 284704 155085 284739 155113
rect 284767 155085 284801 155113
rect 284829 155085 284864 155113
rect 284704 155051 284864 155085
rect 284704 155023 284739 155051
rect 284767 155023 284801 155051
rect 284829 155023 284864 155051
rect 284704 154989 284864 155023
rect 284704 154961 284739 154989
rect 284767 154961 284801 154989
rect 284829 154961 284864 154989
rect 284704 154944 284864 154961
rect 281049 149147 281097 149175
rect 281125 149147 281159 149175
rect 281187 149147 281221 149175
rect 281249 149147 281283 149175
rect 281311 149147 281359 149175
rect 281049 149113 281359 149147
rect 281049 149085 281097 149113
rect 281125 149085 281159 149113
rect 281187 149085 281221 149113
rect 281249 149085 281283 149113
rect 281311 149085 281359 149113
rect 281049 149051 281359 149085
rect 281049 149023 281097 149051
rect 281125 149023 281159 149051
rect 281187 149023 281221 149051
rect 281249 149023 281283 149051
rect 281311 149023 281359 149051
rect 281049 148989 281359 149023
rect 281049 148961 281097 148989
rect 281125 148961 281159 148989
rect 281187 148961 281221 148989
rect 281249 148961 281283 148989
rect 281311 148961 281359 148989
rect 281049 140175 281359 148961
rect 287686 151410 287714 151415
rect 284704 146175 284864 146192
rect 284704 146147 284739 146175
rect 284767 146147 284801 146175
rect 284829 146147 284864 146175
rect 284704 146113 284864 146147
rect 284704 146085 284739 146113
rect 284767 146085 284801 146113
rect 284829 146085 284864 146113
rect 284704 146051 284864 146085
rect 284704 146023 284739 146051
rect 284767 146023 284801 146051
rect 284829 146023 284864 146051
rect 284704 145989 284864 146023
rect 284704 145961 284739 145989
rect 284767 145961 284801 145989
rect 284829 145961 284864 145989
rect 284704 145944 284864 145961
rect 281049 140147 281097 140175
rect 281125 140147 281159 140175
rect 281187 140147 281221 140175
rect 281249 140147 281283 140175
rect 281311 140147 281359 140175
rect 281049 140113 281359 140147
rect 281049 140085 281097 140113
rect 281125 140085 281159 140113
rect 281187 140085 281221 140113
rect 281249 140085 281283 140113
rect 281311 140085 281359 140113
rect 281049 140051 281359 140085
rect 281049 140023 281097 140051
rect 281125 140023 281159 140051
rect 281187 140023 281221 140051
rect 281249 140023 281283 140051
rect 281311 140023 281359 140051
rect 281049 139989 281359 140023
rect 281049 139961 281097 139989
rect 281125 139961 281159 139989
rect 281187 139961 281221 139989
rect 281249 139961 281283 139989
rect 281311 139961 281359 139989
rect 281049 131175 281359 139961
rect 284704 137175 284864 137192
rect 284704 137147 284739 137175
rect 284767 137147 284801 137175
rect 284829 137147 284864 137175
rect 284704 137113 284864 137147
rect 284704 137085 284739 137113
rect 284767 137085 284801 137113
rect 284829 137085 284864 137113
rect 284704 137051 284864 137085
rect 284704 137023 284739 137051
rect 284767 137023 284801 137051
rect 284829 137023 284864 137051
rect 284704 136989 284864 137023
rect 284704 136961 284739 136989
rect 284767 136961 284801 136989
rect 284829 136961 284864 136989
rect 284704 136944 284864 136961
rect 287686 135730 287714 151382
rect 287742 148946 287770 165942
rect 294549 164175 294859 172961
rect 294549 164147 294597 164175
rect 294625 164147 294659 164175
rect 294687 164147 294721 164175
rect 294749 164147 294783 164175
rect 294811 164147 294859 164175
rect 294549 164113 294859 164147
rect 294549 164085 294597 164113
rect 294625 164085 294659 164113
rect 294687 164085 294721 164113
rect 294749 164085 294783 164113
rect 294811 164085 294859 164113
rect 294549 164051 294859 164085
rect 294549 164023 294597 164051
rect 294625 164023 294659 164051
rect 294687 164023 294721 164051
rect 294749 164023 294783 164051
rect 294811 164023 294859 164051
rect 294549 163989 294859 164023
rect 294549 163961 294597 163989
rect 294625 163961 294659 163989
rect 294687 163961 294721 163989
rect 294749 163961 294783 163989
rect 294811 163961 294859 163989
rect 287742 148913 287770 148918
rect 287798 158690 287826 158695
rect 287686 135697 287714 135702
rect 287742 144130 287770 144135
rect 281049 131147 281097 131175
rect 281125 131147 281159 131175
rect 281187 131147 281221 131175
rect 281249 131147 281283 131175
rect 281311 131147 281359 131175
rect 281049 131113 281359 131147
rect 281049 131085 281097 131113
rect 281125 131085 281159 131113
rect 281187 131085 281221 131113
rect 281249 131085 281283 131113
rect 281311 131085 281359 131113
rect 281049 131051 281359 131085
rect 281049 131023 281097 131051
rect 281125 131023 281159 131051
rect 281187 131023 281221 131051
rect 281249 131023 281283 131051
rect 281311 131023 281359 131051
rect 281049 130989 281359 131023
rect 281049 130961 281097 130989
rect 281125 130961 281159 130989
rect 281187 130961 281221 130989
rect 281249 130961 281283 130989
rect 281311 130961 281359 130989
rect 281049 122175 281359 130961
rect 287686 129570 287714 129575
rect 284704 128175 284864 128192
rect 284704 128147 284739 128175
rect 284767 128147 284801 128175
rect 284829 128147 284864 128175
rect 284704 128113 284864 128147
rect 284704 128085 284739 128113
rect 284767 128085 284801 128113
rect 284829 128085 284864 128113
rect 284704 128051 284864 128085
rect 284704 128023 284739 128051
rect 284767 128023 284801 128051
rect 284829 128023 284864 128051
rect 284704 127989 284864 128023
rect 284704 127961 284739 127989
rect 284767 127961 284801 127989
rect 284829 127961 284864 127989
rect 284704 127944 284864 127961
rect 281049 122147 281097 122175
rect 281125 122147 281159 122175
rect 281187 122147 281221 122175
rect 281249 122147 281283 122175
rect 281311 122147 281359 122175
rect 281049 122113 281359 122147
rect 281049 122085 281097 122113
rect 281125 122085 281159 122113
rect 281187 122085 281221 122113
rect 281249 122085 281283 122113
rect 281311 122085 281359 122113
rect 281049 122051 281359 122085
rect 281049 122023 281097 122051
rect 281125 122023 281159 122051
rect 281187 122023 281221 122051
rect 281249 122023 281283 122051
rect 281311 122023 281359 122051
rect 281049 121989 281359 122023
rect 281049 121961 281097 121989
rect 281125 121961 281159 121989
rect 281187 121961 281221 121989
rect 281249 121961 281283 121989
rect 281311 121961 281359 121989
rect 281049 113175 281359 121961
rect 284704 119175 284864 119192
rect 284704 119147 284739 119175
rect 284767 119147 284801 119175
rect 284829 119147 284864 119175
rect 284704 119113 284864 119147
rect 284704 119085 284739 119113
rect 284767 119085 284801 119113
rect 284829 119085 284864 119113
rect 284704 119051 284864 119085
rect 284704 119023 284739 119051
rect 284767 119023 284801 119051
rect 284829 119023 284864 119051
rect 284704 118989 284864 119023
rect 284704 118961 284739 118989
rect 284767 118961 284801 118989
rect 284829 118961 284864 118989
rect 284704 118944 284864 118961
rect 287686 115962 287714 129542
rect 287742 129122 287770 144102
rect 287798 142338 287826 158662
rect 287798 142305 287826 142310
rect 294549 155175 294859 163961
rect 294549 155147 294597 155175
rect 294625 155147 294659 155175
rect 294687 155147 294721 155175
rect 294749 155147 294783 155175
rect 294811 155147 294859 155175
rect 294549 155113 294859 155147
rect 294549 155085 294597 155113
rect 294625 155085 294659 155113
rect 294687 155085 294721 155113
rect 294749 155085 294783 155113
rect 294811 155085 294859 155113
rect 294549 155051 294859 155085
rect 294549 155023 294597 155051
rect 294625 155023 294659 155051
rect 294687 155023 294721 155051
rect 294749 155023 294783 155051
rect 294811 155023 294859 155051
rect 294549 154989 294859 155023
rect 294549 154961 294597 154989
rect 294625 154961 294659 154989
rect 294687 154961 294721 154989
rect 294749 154961 294783 154989
rect 294811 154961 294859 154989
rect 294549 146175 294859 154961
rect 294549 146147 294597 146175
rect 294625 146147 294659 146175
rect 294687 146147 294721 146175
rect 294749 146147 294783 146175
rect 294811 146147 294859 146175
rect 294549 146113 294859 146147
rect 294549 146085 294597 146113
rect 294625 146085 294659 146113
rect 294687 146085 294721 146113
rect 294749 146085 294783 146113
rect 294811 146085 294859 146113
rect 294549 146051 294859 146085
rect 294549 146023 294597 146051
rect 294625 146023 294659 146051
rect 294687 146023 294721 146051
rect 294749 146023 294783 146051
rect 294811 146023 294859 146051
rect 294549 145989 294859 146023
rect 294549 145961 294597 145989
rect 294625 145961 294659 145989
rect 294687 145961 294721 145989
rect 294749 145961 294783 145989
rect 294811 145961 294859 145989
rect 294549 137175 294859 145961
rect 294549 137147 294597 137175
rect 294625 137147 294659 137175
rect 294687 137147 294721 137175
rect 294749 137147 294783 137175
rect 294811 137147 294859 137175
rect 294549 137113 294859 137147
rect 294549 137085 294597 137113
rect 294625 137085 294659 137113
rect 294687 137085 294721 137113
rect 294749 137085 294783 137113
rect 294811 137085 294859 137113
rect 294549 137051 294859 137085
rect 294549 137023 294597 137051
rect 294625 137023 294659 137051
rect 294687 137023 294721 137051
rect 294749 137023 294783 137051
rect 294811 137023 294859 137051
rect 294549 136989 294859 137023
rect 294549 136961 294597 136989
rect 294625 136961 294659 136989
rect 294687 136961 294721 136989
rect 294749 136961 294783 136989
rect 294811 136961 294859 136989
rect 287742 129089 287770 129094
rect 287798 136850 287826 136855
rect 287798 122514 287826 136822
rect 287798 122481 287826 122486
rect 294549 128175 294859 136961
rect 294549 128147 294597 128175
rect 294625 128147 294659 128175
rect 294687 128147 294721 128175
rect 294749 128147 294783 128175
rect 294811 128147 294859 128175
rect 294549 128113 294859 128147
rect 294549 128085 294597 128113
rect 294625 128085 294659 128113
rect 294687 128085 294721 128113
rect 294749 128085 294783 128113
rect 294811 128085 294859 128113
rect 294549 128051 294859 128085
rect 294549 128023 294597 128051
rect 294625 128023 294659 128051
rect 294687 128023 294721 128051
rect 294749 128023 294783 128051
rect 294811 128023 294859 128051
rect 294549 127989 294859 128023
rect 294549 127961 294597 127989
rect 294625 127961 294659 127989
rect 294687 127961 294721 127989
rect 294749 127961 294783 127989
rect 294811 127961 294859 127989
rect 287686 115929 287714 115934
rect 287910 122290 287938 122295
rect 281049 113147 281097 113175
rect 281125 113147 281159 113175
rect 281187 113147 281221 113175
rect 281249 113147 281283 113175
rect 281311 113147 281359 113175
rect 281049 113113 281359 113147
rect 281049 113085 281097 113113
rect 281125 113085 281159 113113
rect 281187 113085 281221 113113
rect 281249 113085 281283 113113
rect 281311 113085 281359 113113
rect 281049 113051 281359 113085
rect 281049 113023 281097 113051
rect 281125 113023 281159 113051
rect 281187 113023 281221 113051
rect 281249 113023 281283 113051
rect 281311 113023 281359 113051
rect 281049 112989 281359 113023
rect 281049 112961 281097 112989
rect 281125 112961 281159 112989
rect 281187 112961 281221 112989
rect 281249 112961 281283 112989
rect 281311 112961 281359 112989
rect 281049 104175 281359 112961
rect 287742 115010 287770 115015
rect 284704 110175 284864 110192
rect 284704 110147 284739 110175
rect 284767 110147 284801 110175
rect 284829 110147 284864 110175
rect 284704 110113 284864 110147
rect 284704 110085 284739 110113
rect 284767 110085 284801 110113
rect 284829 110085 284864 110113
rect 284704 110051 284864 110085
rect 284704 110023 284739 110051
rect 284767 110023 284801 110051
rect 284829 110023 284864 110051
rect 284704 109989 284864 110023
rect 284704 109961 284739 109989
rect 284767 109961 284801 109989
rect 284829 109961 284864 109989
rect 284704 109944 284864 109961
rect 281049 104147 281097 104175
rect 281125 104147 281159 104175
rect 281187 104147 281221 104175
rect 281249 104147 281283 104175
rect 281311 104147 281359 104175
rect 281049 104113 281359 104147
rect 281049 104085 281097 104113
rect 281125 104085 281159 104113
rect 281187 104085 281221 104113
rect 281249 104085 281283 104113
rect 281311 104085 281359 104113
rect 281049 104051 281359 104085
rect 281049 104023 281097 104051
rect 281125 104023 281159 104051
rect 281187 104023 281221 104051
rect 281249 104023 281283 104051
rect 281311 104023 281359 104051
rect 281049 103989 281359 104023
rect 281049 103961 281097 103989
rect 281125 103961 281159 103989
rect 281187 103961 281221 103989
rect 281249 103961 281283 103989
rect 281311 103961 281359 103989
rect 281049 95175 281359 103961
rect 287686 107730 287714 107735
rect 284704 101175 284864 101192
rect 284704 101147 284739 101175
rect 284767 101147 284801 101175
rect 284829 101147 284864 101175
rect 284704 101113 284864 101147
rect 284704 101085 284739 101113
rect 284767 101085 284801 101113
rect 284829 101085 284864 101113
rect 284704 101051 284864 101085
rect 284704 101023 284739 101051
rect 284767 101023 284801 101051
rect 284829 101023 284864 101051
rect 284704 100989 284864 101023
rect 284704 100961 284739 100989
rect 284767 100961 284801 100989
rect 284829 100961 284864 100989
rect 284704 100944 284864 100961
rect 287686 96082 287714 107702
rect 287742 102690 287770 114982
rect 287910 109298 287938 122262
rect 287910 109265 287938 109270
rect 294549 119175 294859 127961
rect 294549 119147 294597 119175
rect 294625 119147 294659 119175
rect 294687 119147 294721 119175
rect 294749 119147 294783 119175
rect 294811 119147 294859 119175
rect 294549 119113 294859 119147
rect 294549 119085 294597 119113
rect 294625 119085 294659 119113
rect 294687 119085 294721 119113
rect 294749 119085 294783 119113
rect 294811 119085 294859 119113
rect 294549 119051 294859 119085
rect 294549 119023 294597 119051
rect 294625 119023 294659 119051
rect 294687 119023 294721 119051
rect 294749 119023 294783 119051
rect 294811 119023 294859 119051
rect 294549 118989 294859 119023
rect 294549 118961 294597 118989
rect 294625 118961 294659 118989
rect 294687 118961 294721 118989
rect 294749 118961 294783 118989
rect 294811 118961 294859 118989
rect 294549 110175 294859 118961
rect 294549 110147 294597 110175
rect 294625 110147 294659 110175
rect 294687 110147 294721 110175
rect 294749 110147 294783 110175
rect 294811 110147 294859 110175
rect 294549 110113 294859 110147
rect 294549 110085 294597 110113
rect 294625 110085 294659 110113
rect 294687 110085 294721 110113
rect 294749 110085 294783 110113
rect 294811 110085 294859 110113
rect 294549 110051 294859 110085
rect 294549 110023 294597 110051
rect 294625 110023 294659 110051
rect 294687 110023 294721 110051
rect 294749 110023 294783 110051
rect 294811 110023 294859 110051
rect 294549 109989 294859 110023
rect 294549 109961 294597 109989
rect 294625 109961 294659 109989
rect 294687 109961 294721 109989
rect 294749 109961 294783 109989
rect 294811 109961 294859 109989
rect 287742 102657 287770 102662
rect 294549 101175 294859 109961
rect 294549 101147 294597 101175
rect 294625 101147 294659 101175
rect 294687 101147 294721 101175
rect 294749 101147 294783 101175
rect 294811 101147 294859 101175
rect 294549 101113 294859 101147
rect 294549 101085 294597 101113
rect 294625 101085 294659 101113
rect 294687 101085 294721 101113
rect 294749 101085 294783 101113
rect 294811 101085 294859 101113
rect 294549 101051 294859 101085
rect 294549 101023 294597 101051
rect 294625 101023 294659 101051
rect 294687 101023 294721 101051
rect 294749 101023 294783 101051
rect 294811 101023 294859 101051
rect 294549 100989 294859 101023
rect 294549 100961 294597 100989
rect 294625 100961 294659 100989
rect 294687 100961 294721 100989
rect 294749 100961 294783 100989
rect 294811 100961 294859 100989
rect 287686 96049 287714 96054
rect 287742 100450 287770 100455
rect 281049 95147 281097 95175
rect 281125 95147 281159 95175
rect 281187 95147 281221 95175
rect 281249 95147 281283 95175
rect 281311 95147 281359 95175
rect 281049 95113 281359 95147
rect 281049 95085 281097 95113
rect 281125 95085 281159 95113
rect 281187 95085 281221 95113
rect 281249 95085 281283 95113
rect 281311 95085 281359 95113
rect 281049 95051 281359 95085
rect 281049 95023 281097 95051
rect 281125 95023 281159 95051
rect 281187 95023 281221 95051
rect 281249 95023 281283 95051
rect 281311 95023 281359 95051
rect 281049 94989 281359 95023
rect 281049 94961 281097 94989
rect 281125 94961 281159 94989
rect 281187 94961 281221 94989
rect 281249 94961 281283 94989
rect 281311 94961 281359 94989
rect 281049 86175 281359 94961
rect 284704 92175 284864 92192
rect 284704 92147 284739 92175
rect 284767 92147 284801 92175
rect 284829 92147 284864 92175
rect 284704 92113 284864 92147
rect 284704 92085 284739 92113
rect 284767 92085 284801 92113
rect 284829 92085 284864 92113
rect 284704 92051 284864 92085
rect 284704 92023 284739 92051
rect 284767 92023 284801 92051
rect 284829 92023 284864 92051
rect 284704 91989 284864 92023
rect 284704 91961 284739 91989
rect 284767 91961 284801 91989
rect 284829 91961 284864 91989
rect 284704 91944 284864 91961
rect 287742 89474 287770 100422
rect 287742 89441 287770 89446
rect 287798 93170 287826 93175
rect 281049 86147 281097 86175
rect 281125 86147 281159 86175
rect 281187 86147 281221 86175
rect 281249 86147 281283 86175
rect 281311 86147 281359 86175
rect 281049 86113 281359 86147
rect 281049 86085 281097 86113
rect 281125 86085 281159 86113
rect 281187 86085 281221 86113
rect 281249 86085 281283 86113
rect 281311 86085 281359 86113
rect 281049 86051 281359 86085
rect 281049 86023 281097 86051
rect 281125 86023 281159 86051
rect 281187 86023 281221 86051
rect 281249 86023 281283 86051
rect 281311 86023 281359 86051
rect 281049 85989 281359 86023
rect 281049 85961 281097 85989
rect 281125 85961 281159 85989
rect 281187 85961 281221 85989
rect 281249 85961 281283 85989
rect 281311 85961 281359 85989
rect 281049 77175 281359 85961
rect 287686 85890 287714 85895
rect 284704 83175 284864 83192
rect 284704 83147 284739 83175
rect 284767 83147 284801 83175
rect 284829 83147 284864 83175
rect 284704 83113 284864 83147
rect 284704 83085 284739 83113
rect 284767 83085 284801 83113
rect 284829 83085 284864 83113
rect 284704 83051 284864 83085
rect 284704 83023 284739 83051
rect 284767 83023 284801 83051
rect 284829 83023 284864 83051
rect 284704 82989 284864 83023
rect 284704 82961 284739 82989
rect 284767 82961 284801 82989
rect 284829 82961 284864 82989
rect 284704 82944 284864 82961
rect 281049 77147 281097 77175
rect 281125 77147 281159 77175
rect 281187 77147 281221 77175
rect 281249 77147 281283 77175
rect 281311 77147 281359 77175
rect 281049 77113 281359 77147
rect 281049 77085 281097 77113
rect 281125 77085 281159 77113
rect 281187 77085 281221 77113
rect 281249 77085 281283 77113
rect 281311 77085 281359 77113
rect 281049 77051 281359 77085
rect 281049 77023 281097 77051
rect 281125 77023 281159 77051
rect 281187 77023 281221 77051
rect 281249 77023 281283 77051
rect 281311 77023 281359 77051
rect 281049 76989 281359 77023
rect 281049 76961 281097 76989
rect 281125 76961 281159 76989
rect 281187 76961 281221 76989
rect 281249 76961 281283 76989
rect 281311 76961 281359 76989
rect 281049 68175 281359 76961
rect 287686 76258 287714 85862
rect 287798 82866 287826 93142
rect 287798 82833 287826 82838
rect 294549 92175 294859 100961
rect 294549 92147 294597 92175
rect 294625 92147 294659 92175
rect 294687 92147 294721 92175
rect 294749 92147 294783 92175
rect 294811 92147 294859 92175
rect 294549 92113 294859 92147
rect 294549 92085 294597 92113
rect 294625 92085 294659 92113
rect 294687 92085 294721 92113
rect 294749 92085 294783 92113
rect 294811 92085 294859 92113
rect 294549 92051 294859 92085
rect 294549 92023 294597 92051
rect 294625 92023 294659 92051
rect 294687 92023 294721 92051
rect 294749 92023 294783 92051
rect 294811 92023 294859 92051
rect 294549 91989 294859 92023
rect 294549 91961 294597 91989
rect 294625 91961 294659 91989
rect 294687 91961 294721 91989
rect 294749 91961 294783 91989
rect 294811 91961 294859 91989
rect 294549 83175 294859 91961
rect 294549 83147 294597 83175
rect 294625 83147 294659 83175
rect 294687 83147 294721 83175
rect 294749 83147 294783 83175
rect 294811 83147 294859 83175
rect 294549 83113 294859 83147
rect 294549 83085 294597 83113
rect 294625 83085 294659 83113
rect 294687 83085 294721 83113
rect 294749 83085 294783 83113
rect 294811 83085 294859 83113
rect 294549 83051 294859 83085
rect 294549 83023 294597 83051
rect 294625 83023 294659 83051
rect 294687 83023 294721 83051
rect 294749 83023 294783 83051
rect 294811 83023 294859 83051
rect 294549 82989 294859 83023
rect 294549 82961 294597 82989
rect 294625 82961 294659 82989
rect 294687 82961 294721 82989
rect 294749 82961 294783 82989
rect 294811 82961 294859 82989
rect 287686 76225 287714 76230
rect 287742 78610 287770 78615
rect 284704 74175 284864 74192
rect 284704 74147 284739 74175
rect 284767 74147 284801 74175
rect 284829 74147 284864 74175
rect 284704 74113 284864 74147
rect 284704 74085 284739 74113
rect 284767 74085 284801 74113
rect 284829 74085 284864 74113
rect 284704 74051 284864 74085
rect 284704 74023 284739 74051
rect 284767 74023 284801 74051
rect 284829 74023 284864 74051
rect 284704 73989 284864 74023
rect 284704 73961 284739 73989
rect 284767 73961 284801 73989
rect 284829 73961 284864 73989
rect 284704 73944 284864 73961
rect 287742 69650 287770 78582
rect 294549 74175 294859 82961
rect 294549 74147 294597 74175
rect 294625 74147 294659 74175
rect 294687 74147 294721 74175
rect 294749 74147 294783 74175
rect 294811 74147 294859 74175
rect 294549 74113 294859 74147
rect 294549 74085 294597 74113
rect 294625 74085 294659 74113
rect 294687 74085 294721 74113
rect 294749 74085 294783 74113
rect 294811 74085 294859 74113
rect 294549 74051 294859 74085
rect 294549 74023 294597 74051
rect 294625 74023 294659 74051
rect 294687 74023 294721 74051
rect 294749 74023 294783 74051
rect 294811 74023 294859 74051
rect 294549 73989 294859 74023
rect 294549 73961 294597 73989
rect 294625 73961 294659 73989
rect 294687 73961 294721 73989
rect 294749 73961 294783 73989
rect 294811 73961 294859 73989
rect 287742 69617 287770 69622
rect 287798 71330 287826 71335
rect 281049 68147 281097 68175
rect 281125 68147 281159 68175
rect 281187 68147 281221 68175
rect 281249 68147 281283 68175
rect 281311 68147 281359 68175
rect 281049 68113 281359 68147
rect 281049 68085 281097 68113
rect 281125 68085 281159 68113
rect 281187 68085 281221 68113
rect 281249 68085 281283 68113
rect 281311 68085 281359 68113
rect 281049 68051 281359 68085
rect 281049 68023 281097 68051
rect 281125 68023 281159 68051
rect 281187 68023 281221 68051
rect 281249 68023 281283 68051
rect 281311 68023 281359 68051
rect 281049 67989 281359 68023
rect 281049 67961 281097 67989
rect 281125 67961 281159 67989
rect 281187 67961 281221 67989
rect 281249 67961 281283 67989
rect 281311 67961 281359 67989
rect 281049 59175 281359 67961
rect 284704 65175 284864 65192
rect 284704 65147 284739 65175
rect 284767 65147 284801 65175
rect 284829 65147 284864 65175
rect 284704 65113 284864 65147
rect 284704 65085 284739 65113
rect 284767 65085 284801 65113
rect 284829 65085 284864 65113
rect 284704 65051 284864 65085
rect 284704 65023 284739 65051
rect 284767 65023 284801 65051
rect 284829 65023 284864 65051
rect 284704 64989 284864 65023
rect 284704 64961 284739 64989
rect 284767 64961 284801 64989
rect 284829 64961 284864 64989
rect 284704 64944 284864 64961
rect 281049 59147 281097 59175
rect 281125 59147 281159 59175
rect 281187 59147 281221 59175
rect 281249 59147 281283 59175
rect 281311 59147 281359 59175
rect 281049 59113 281359 59147
rect 281049 59085 281097 59113
rect 281125 59085 281159 59113
rect 281187 59085 281221 59113
rect 281249 59085 281283 59113
rect 281311 59085 281359 59113
rect 281049 59051 281359 59085
rect 281049 59023 281097 59051
rect 281125 59023 281159 59051
rect 281187 59023 281221 59051
rect 281249 59023 281283 59051
rect 281311 59023 281359 59051
rect 281049 58989 281359 59023
rect 281049 58961 281097 58989
rect 281125 58961 281159 58989
rect 281187 58961 281221 58989
rect 281249 58961 281283 58989
rect 281311 58961 281359 58989
rect 281049 50175 281359 58961
rect 287686 64050 287714 64055
rect 287686 56434 287714 64022
rect 287798 63042 287826 71302
rect 287798 63009 287826 63014
rect 294549 65175 294859 73961
rect 294549 65147 294597 65175
rect 294625 65147 294659 65175
rect 294687 65147 294721 65175
rect 294749 65147 294783 65175
rect 294811 65147 294859 65175
rect 294549 65113 294859 65147
rect 294549 65085 294597 65113
rect 294625 65085 294659 65113
rect 294687 65085 294721 65113
rect 294749 65085 294783 65113
rect 294811 65085 294859 65113
rect 294549 65051 294859 65085
rect 294549 65023 294597 65051
rect 294625 65023 294659 65051
rect 294687 65023 294721 65051
rect 294749 65023 294783 65051
rect 294811 65023 294859 65051
rect 294549 64989 294859 65023
rect 294549 64961 294597 64989
rect 294625 64961 294659 64989
rect 294687 64961 294721 64989
rect 294749 64961 294783 64989
rect 294811 64961 294859 64989
rect 287686 56401 287714 56406
rect 284704 56175 284864 56192
rect 284704 56147 284739 56175
rect 284767 56147 284801 56175
rect 284829 56147 284864 56175
rect 284704 56113 284864 56147
rect 284704 56085 284739 56113
rect 284767 56085 284801 56113
rect 284829 56085 284864 56113
rect 284704 56051 284864 56085
rect 284704 56023 284739 56051
rect 284767 56023 284801 56051
rect 284829 56023 284864 56051
rect 284704 55989 284864 56023
rect 284704 55961 284739 55989
rect 284767 55961 284801 55989
rect 284829 55961 284864 55989
rect 284704 55944 284864 55961
rect 294549 56175 294859 64961
rect 296409 299086 296719 299134
rect 296409 299058 296457 299086
rect 296485 299058 296519 299086
rect 296547 299058 296581 299086
rect 296609 299058 296643 299086
rect 296671 299058 296719 299086
rect 296409 299024 296719 299058
rect 296409 298996 296457 299024
rect 296485 298996 296519 299024
rect 296547 298996 296581 299024
rect 296609 298996 296643 299024
rect 296671 298996 296719 299024
rect 296409 298962 296719 298996
rect 296409 298934 296457 298962
rect 296485 298934 296519 298962
rect 296547 298934 296581 298962
rect 296609 298934 296643 298962
rect 296671 298934 296719 298962
rect 296409 298900 296719 298934
rect 296409 298872 296457 298900
rect 296485 298872 296519 298900
rect 296547 298872 296581 298900
rect 296609 298872 296643 298900
rect 296671 298872 296719 298900
rect 296409 293175 296719 298872
rect 298680 299086 298990 299134
rect 298680 299058 298728 299086
rect 298756 299058 298790 299086
rect 298818 299058 298852 299086
rect 298880 299058 298914 299086
rect 298942 299058 298990 299086
rect 298680 299024 298990 299058
rect 298680 298996 298728 299024
rect 298756 298996 298790 299024
rect 298818 298996 298852 299024
rect 298880 298996 298914 299024
rect 298942 298996 298990 299024
rect 298680 298962 298990 298996
rect 298680 298934 298728 298962
rect 298756 298934 298790 298962
rect 298818 298934 298852 298962
rect 298880 298934 298914 298962
rect 298942 298934 298990 298962
rect 298680 298900 298990 298934
rect 298680 298872 298728 298900
rect 298756 298872 298790 298900
rect 298818 298872 298852 298900
rect 298880 298872 298914 298900
rect 298942 298872 298990 298900
rect 296409 293147 296457 293175
rect 296485 293147 296519 293175
rect 296547 293147 296581 293175
rect 296609 293147 296643 293175
rect 296671 293147 296719 293175
rect 296409 293113 296719 293147
rect 296409 293085 296457 293113
rect 296485 293085 296519 293113
rect 296547 293085 296581 293113
rect 296609 293085 296643 293113
rect 296671 293085 296719 293113
rect 296409 293051 296719 293085
rect 296409 293023 296457 293051
rect 296485 293023 296519 293051
rect 296547 293023 296581 293051
rect 296609 293023 296643 293051
rect 296671 293023 296719 293051
rect 296409 292989 296719 293023
rect 296409 292961 296457 292989
rect 296485 292961 296519 292989
rect 296547 292961 296581 292989
rect 296609 292961 296643 292989
rect 296671 292961 296719 292989
rect 296409 284175 296719 292961
rect 296409 284147 296457 284175
rect 296485 284147 296519 284175
rect 296547 284147 296581 284175
rect 296609 284147 296643 284175
rect 296671 284147 296719 284175
rect 296409 284113 296719 284147
rect 296409 284085 296457 284113
rect 296485 284085 296519 284113
rect 296547 284085 296581 284113
rect 296609 284085 296643 284113
rect 296671 284085 296719 284113
rect 296409 284051 296719 284085
rect 296409 284023 296457 284051
rect 296485 284023 296519 284051
rect 296547 284023 296581 284051
rect 296609 284023 296643 284051
rect 296671 284023 296719 284051
rect 296409 283989 296719 284023
rect 296409 283961 296457 283989
rect 296485 283961 296519 283989
rect 296547 283961 296581 283989
rect 296609 283961 296643 283989
rect 296671 283961 296719 283989
rect 296409 275175 296719 283961
rect 296409 275147 296457 275175
rect 296485 275147 296519 275175
rect 296547 275147 296581 275175
rect 296609 275147 296643 275175
rect 296671 275147 296719 275175
rect 296409 275113 296719 275147
rect 296409 275085 296457 275113
rect 296485 275085 296519 275113
rect 296547 275085 296581 275113
rect 296609 275085 296643 275113
rect 296671 275085 296719 275113
rect 296409 275051 296719 275085
rect 296409 275023 296457 275051
rect 296485 275023 296519 275051
rect 296547 275023 296581 275051
rect 296609 275023 296643 275051
rect 296671 275023 296719 275051
rect 296409 274989 296719 275023
rect 296409 274961 296457 274989
rect 296485 274961 296519 274989
rect 296547 274961 296581 274989
rect 296609 274961 296643 274989
rect 296671 274961 296719 274989
rect 296409 266175 296719 274961
rect 296409 266147 296457 266175
rect 296485 266147 296519 266175
rect 296547 266147 296581 266175
rect 296609 266147 296643 266175
rect 296671 266147 296719 266175
rect 296409 266113 296719 266147
rect 296409 266085 296457 266113
rect 296485 266085 296519 266113
rect 296547 266085 296581 266113
rect 296609 266085 296643 266113
rect 296671 266085 296719 266113
rect 296409 266051 296719 266085
rect 296409 266023 296457 266051
rect 296485 266023 296519 266051
rect 296547 266023 296581 266051
rect 296609 266023 296643 266051
rect 296671 266023 296719 266051
rect 296409 265989 296719 266023
rect 296409 265961 296457 265989
rect 296485 265961 296519 265989
rect 296547 265961 296581 265989
rect 296609 265961 296643 265989
rect 296671 265961 296719 265989
rect 296409 257175 296719 265961
rect 296409 257147 296457 257175
rect 296485 257147 296519 257175
rect 296547 257147 296581 257175
rect 296609 257147 296643 257175
rect 296671 257147 296719 257175
rect 296409 257113 296719 257147
rect 296409 257085 296457 257113
rect 296485 257085 296519 257113
rect 296547 257085 296581 257113
rect 296609 257085 296643 257113
rect 296671 257085 296719 257113
rect 296409 257051 296719 257085
rect 296409 257023 296457 257051
rect 296485 257023 296519 257051
rect 296547 257023 296581 257051
rect 296609 257023 296643 257051
rect 296671 257023 296719 257051
rect 296409 256989 296719 257023
rect 296409 256961 296457 256989
rect 296485 256961 296519 256989
rect 296547 256961 296581 256989
rect 296609 256961 296643 256989
rect 296671 256961 296719 256989
rect 296409 248175 296719 256961
rect 296409 248147 296457 248175
rect 296485 248147 296519 248175
rect 296547 248147 296581 248175
rect 296609 248147 296643 248175
rect 296671 248147 296719 248175
rect 296409 248113 296719 248147
rect 296409 248085 296457 248113
rect 296485 248085 296519 248113
rect 296547 248085 296581 248113
rect 296609 248085 296643 248113
rect 296671 248085 296719 248113
rect 296409 248051 296719 248085
rect 296409 248023 296457 248051
rect 296485 248023 296519 248051
rect 296547 248023 296581 248051
rect 296609 248023 296643 248051
rect 296671 248023 296719 248051
rect 296409 247989 296719 248023
rect 296409 247961 296457 247989
rect 296485 247961 296519 247989
rect 296547 247961 296581 247989
rect 296609 247961 296643 247989
rect 296671 247961 296719 247989
rect 296409 239175 296719 247961
rect 296409 239147 296457 239175
rect 296485 239147 296519 239175
rect 296547 239147 296581 239175
rect 296609 239147 296643 239175
rect 296671 239147 296719 239175
rect 296409 239113 296719 239147
rect 296409 239085 296457 239113
rect 296485 239085 296519 239113
rect 296547 239085 296581 239113
rect 296609 239085 296643 239113
rect 296671 239085 296719 239113
rect 296409 239051 296719 239085
rect 296409 239023 296457 239051
rect 296485 239023 296519 239051
rect 296547 239023 296581 239051
rect 296609 239023 296643 239051
rect 296671 239023 296719 239051
rect 296409 238989 296719 239023
rect 296409 238961 296457 238989
rect 296485 238961 296519 238989
rect 296547 238961 296581 238989
rect 296609 238961 296643 238989
rect 296671 238961 296719 238989
rect 296409 230175 296719 238961
rect 296409 230147 296457 230175
rect 296485 230147 296519 230175
rect 296547 230147 296581 230175
rect 296609 230147 296643 230175
rect 296671 230147 296719 230175
rect 296409 230113 296719 230147
rect 296409 230085 296457 230113
rect 296485 230085 296519 230113
rect 296547 230085 296581 230113
rect 296609 230085 296643 230113
rect 296671 230085 296719 230113
rect 296409 230051 296719 230085
rect 296409 230023 296457 230051
rect 296485 230023 296519 230051
rect 296547 230023 296581 230051
rect 296609 230023 296643 230051
rect 296671 230023 296719 230051
rect 296409 229989 296719 230023
rect 296409 229961 296457 229989
rect 296485 229961 296519 229989
rect 296547 229961 296581 229989
rect 296609 229961 296643 229989
rect 296671 229961 296719 229989
rect 296409 221175 296719 229961
rect 296409 221147 296457 221175
rect 296485 221147 296519 221175
rect 296547 221147 296581 221175
rect 296609 221147 296643 221175
rect 296671 221147 296719 221175
rect 296409 221113 296719 221147
rect 296409 221085 296457 221113
rect 296485 221085 296519 221113
rect 296547 221085 296581 221113
rect 296609 221085 296643 221113
rect 296671 221085 296719 221113
rect 296409 221051 296719 221085
rect 296409 221023 296457 221051
rect 296485 221023 296519 221051
rect 296547 221023 296581 221051
rect 296609 221023 296643 221051
rect 296671 221023 296719 221051
rect 296409 220989 296719 221023
rect 296409 220961 296457 220989
rect 296485 220961 296519 220989
rect 296547 220961 296581 220989
rect 296609 220961 296643 220989
rect 296671 220961 296719 220989
rect 296409 212175 296719 220961
rect 296409 212147 296457 212175
rect 296485 212147 296519 212175
rect 296547 212147 296581 212175
rect 296609 212147 296643 212175
rect 296671 212147 296719 212175
rect 296409 212113 296719 212147
rect 296409 212085 296457 212113
rect 296485 212085 296519 212113
rect 296547 212085 296581 212113
rect 296609 212085 296643 212113
rect 296671 212085 296719 212113
rect 296409 212051 296719 212085
rect 296409 212023 296457 212051
rect 296485 212023 296519 212051
rect 296547 212023 296581 212051
rect 296609 212023 296643 212051
rect 296671 212023 296719 212051
rect 296409 211989 296719 212023
rect 296409 211961 296457 211989
rect 296485 211961 296519 211989
rect 296547 211961 296581 211989
rect 296609 211961 296643 211989
rect 296671 211961 296719 211989
rect 296409 203175 296719 211961
rect 296409 203147 296457 203175
rect 296485 203147 296519 203175
rect 296547 203147 296581 203175
rect 296609 203147 296643 203175
rect 296671 203147 296719 203175
rect 296409 203113 296719 203147
rect 296409 203085 296457 203113
rect 296485 203085 296519 203113
rect 296547 203085 296581 203113
rect 296609 203085 296643 203113
rect 296671 203085 296719 203113
rect 296409 203051 296719 203085
rect 296409 203023 296457 203051
rect 296485 203023 296519 203051
rect 296547 203023 296581 203051
rect 296609 203023 296643 203051
rect 296671 203023 296719 203051
rect 296409 202989 296719 203023
rect 296409 202961 296457 202989
rect 296485 202961 296519 202989
rect 296547 202961 296581 202989
rect 296609 202961 296643 202989
rect 296671 202961 296719 202989
rect 296409 194175 296719 202961
rect 296409 194147 296457 194175
rect 296485 194147 296519 194175
rect 296547 194147 296581 194175
rect 296609 194147 296643 194175
rect 296671 194147 296719 194175
rect 296409 194113 296719 194147
rect 296409 194085 296457 194113
rect 296485 194085 296519 194113
rect 296547 194085 296581 194113
rect 296609 194085 296643 194113
rect 296671 194085 296719 194113
rect 296409 194051 296719 194085
rect 296409 194023 296457 194051
rect 296485 194023 296519 194051
rect 296547 194023 296581 194051
rect 296609 194023 296643 194051
rect 296671 194023 296719 194051
rect 296409 193989 296719 194023
rect 296409 193961 296457 193989
rect 296485 193961 296519 193989
rect 296547 193961 296581 193989
rect 296609 193961 296643 193989
rect 296671 193961 296719 193989
rect 296409 185175 296719 193961
rect 296409 185147 296457 185175
rect 296485 185147 296519 185175
rect 296547 185147 296581 185175
rect 296609 185147 296643 185175
rect 296671 185147 296719 185175
rect 296409 185113 296719 185147
rect 296409 185085 296457 185113
rect 296485 185085 296519 185113
rect 296547 185085 296581 185113
rect 296609 185085 296643 185113
rect 296671 185085 296719 185113
rect 296409 185051 296719 185085
rect 296409 185023 296457 185051
rect 296485 185023 296519 185051
rect 296547 185023 296581 185051
rect 296609 185023 296643 185051
rect 296671 185023 296719 185051
rect 296409 184989 296719 185023
rect 296409 184961 296457 184989
rect 296485 184961 296519 184989
rect 296547 184961 296581 184989
rect 296609 184961 296643 184989
rect 296671 184961 296719 184989
rect 296409 176175 296719 184961
rect 296409 176147 296457 176175
rect 296485 176147 296519 176175
rect 296547 176147 296581 176175
rect 296609 176147 296643 176175
rect 296671 176147 296719 176175
rect 296409 176113 296719 176147
rect 296409 176085 296457 176113
rect 296485 176085 296519 176113
rect 296547 176085 296581 176113
rect 296609 176085 296643 176113
rect 296671 176085 296719 176113
rect 296409 176051 296719 176085
rect 296409 176023 296457 176051
rect 296485 176023 296519 176051
rect 296547 176023 296581 176051
rect 296609 176023 296643 176051
rect 296671 176023 296719 176051
rect 296409 175989 296719 176023
rect 296409 175961 296457 175989
rect 296485 175961 296519 175989
rect 296547 175961 296581 175989
rect 296609 175961 296643 175989
rect 296671 175961 296719 175989
rect 296409 167175 296719 175961
rect 296409 167147 296457 167175
rect 296485 167147 296519 167175
rect 296547 167147 296581 167175
rect 296609 167147 296643 167175
rect 296671 167147 296719 167175
rect 296409 167113 296719 167147
rect 296409 167085 296457 167113
rect 296485 167085 296519 167113
rect 296547 167085 296581 167113
rect 296609 167085 296643 167113
rect 296671 167085 296719 167113
rect 296409 167051 296719 167085
rect 296409 167023 296457 167051
rect 296485 167023 296519 167051
rect 296547 167023 296581 167051
rect 296609 167023 296643 167051
rect 296671 167023 296719 167051
rect 296409 166989 296719 167023
rect 296409 166961 296457 166989
rect 296485 166961 296519 166989
rect 296547 166961 296581 166989
rect 296609 166961 296643 166989
rect 296671 166961 296719 166989
rect 296409 158175 296719 166961
rect 296409 158147 296457 158175
rect 296485 158147 296519 158175
rect 296547 158147 296581 158175
rect 296609 158147 296643 158175
rect 296671 158147 296719 158175
rect 296409 158113 296719 158147
rect 296409 158085 296457 158113
rect 296485 158085 296519 158113
rect 296547 158085 296581 158113
rect 296609 158085 296643 158113
rect 296671 158085 296719 158113
rect 296409 158051 296719 158085
rect 296409 158023 296457 158051
rect 296485 158023 296519 158051
rect 296547 158023 296581 158051
rect 296609 158023 296643 158051
rect 296671 158023 296719 158051
rect 296409 157989 296719 158023
rect 296409 157961 296457 157989
rect 296485 157961 296519 157989
rect 296547 157961 296581 157989
rect 296609 157961 296643 157989
rect 296671 157961 296719 157989
rect 296409 149175 296719 157961
rect 296409 149147 296457 149175
rect 296485 149147 296519 149175
rect 296547 149147 296581 149175
rect 296609 149147 296643 149175
rect 296671 149147 296719 149175
rect 296409 149113 296719 149147
rect 296409 149085 296457 149113
rect 296485 149085 296519 149113
rect 296547 149085 296581 149113
rect 296609 149085 296643 149113
rect 296671 149085 296719 149113
rect 296409 149051 296719 149085
rect 296409 149023 296457 149051
rect 296485 149023 296519 149051
rect 296547 149023 296581 149051
rect 296609 149023 296643 149051
rect 296671 149023 296719 149051
rect 296409 148989 296719 149023
rect 296409 148961 296457 148989
rect 296485 148961 296519 148989
rect 296547 148961 296581 148989
rect 296609 148961 296643 148989
rect 296671 148961 296719 148989
rect 296409 140175 296719 148961
rect 296409 140147 296457 140175
rect 296485 140147 296519 140175
rect 296547 140147 296581 140175
rect 296609 140147 296643 140175
rect 296671 140147 296719 140175
rect 296409 140113 296719 140147
rect 296409 140085 296457 140113
rect 296485 140085 296519 140113
rect 296547 140085 296581 140113
rect 296609 140085 296643 140113
rect 296671 140085 296719 140113
rect 296409 140051 296719 140085
rect 296409 140023 296457 140051
rect 296485 140023 296519 140051
rect 296547 140023 296581 140051
rect 296609 140023 296643 140051
rect 296671 140023 296719 140051
rect 296409 139989 296719 140023
rect 296409 139961 296457 139989
rect 296485 139961 296519 139989
rect 296547 139961 296581 139989
rect 296609 139961 296643 139989
rect 296671 139961 296719 139989
rect 296409 131175 296719 139961
rect 296409 131147 296457 131175
rect 296485 131147 296519 131175
rect 296547 131147 296581 131175
rect 296609 131147 296643 131175
rect 296671 131147 296719 131175
rect 296409 131113 296719 131147
rect 296409 131085 296457 131113
rect 296485 131085 296519 131113
rect 296547 131085 296581 131113
rect 296609 131085 296643 131113
rect 296671 131085 296719 131113
rect 296409 131051 296719 131085
rect 296409 131023 296457 131051
rect 296485 131023 296519 131051
rect 296547 131023 296581 131051
rect 296609 131023 296643 131051
rect 296671 131023 296719 131051
rect 296409 130989 296719 131023
rect 296409 130961 296457 130989
rect 296485 130961 296519 130989
rect 296547 130961 296581 130989
rect 296609 130961 296643 130989
rect 296671 130961 296719 130989
rect 296409 122175 296719 130961
rect 296409 122147 296457 122175
rect 296485 122147 296519 122175
rect 296547 122147 296581 122175
rect 296609 122147 296643 122175
rect 296671 122147 296719 122175
rect 296409 122113 296719 122147
rect 296409 122085 296457 122113
rect 296485 122085 296519 122113
rect 296547 122085 296581 122113
rect 296609 122085 296643 122113
rect 296671 122085 296719 122113
rect 296409 122051 296719 122085
rect 296409 122023 296457 122051
rect 296485 122023 296519 122051
rect 296547 122023 296581 122051
rect 296609 122023 296643 122051
rect 296671 122023 296719 122051
rect 296409 121989 296719 122023
rect 296409 121961 296457 121989
rect 296485 121961 296519 121989
rect 296547 121961 296581 121989
rect 296609 121961 296643 121989
rect 296671 121961 296719 121989
rect 296409 113175 296719 121961
rect 296409 113147 296457 113175
rect 296485 113147 296519 113175
rect 296547 113147 296581 113175
rect 296609 113147 296643 113175
rect 296671 113147 296719 113175
rect 296409 113113 296719 113147
rect 296409 113085 296457 113113
rect 296485 113085 296519 113113
rect 296547 113085 296581 113113
rect 296609 113085 296643 113113
rect 296671 113085 296719 113113
rect 296409 113051 296719 113085
rect 296409 113023 296457 113051
rect 296485 113023 296519 113051
rect 296547 113023 296581 113051
rect 296609 113023 296643 113051
rect 296671 113023 296719 113051
rect 296409 112989 296719 113023
rect 296409 112961 296457 112989
rect 296485 112961 296519 112989
rect 296547 112961 296581 112989
rect 296609 112961 296643 112989
rect 296671 112961 296719 112989
rect 296409 104175 296719 112961
rect 296409 104147 296457 104175
rect 296485 104147 296519 104175
rect 296547 104147 296581 104175
rect 296609 104147 296643 104175
rect 296671 104147 296719 104175
rect 296409 104113 296719 104147
rect 296409 104085 296457 104113
rect 296485 104085 296519 104113
rect 296547 104085 296581 104113
rect 296609 104085 296643 104113
rect 296671 104085 296719 104113
rect 296409 104051 296719 104085
rect 296409 104023 296457 104051
rect 296485 104023 296519 104051
rect 296547 104023 296581 104051
rect 296609 104023 296643 104051
rect 296671 104023 296719 104051
rect 296409 103989 296719 104023
rect 296409 103961 296457 103989
rect 296485 103961 296519 103989
rect 296547 103961 296581 103989
rect 296609 103961 296643 103989
rect 296671 103961 296719 103989
rect 296409 95175 296719 103961
rect 296409 95147 296457 95175
rect 296485 95147 296519 95175
rect 296547 95147 296581 95175
rect 296609 95147 296643 95175
rect 296671 95147 296719 95175
rect 296409 95113 296719 95147
rect 296409 95085 296457 95113
rect 296485 95085 296519 95113
rect 296547 95085 296581 95113
rect 296609 95085 296643 95113
rect 296671 95085 296719 95113
rect 296409 95051 296719 95085
rect 296409 95023 296457 95051
rect 296485 95023 296519 95051
rect 296547 95023 296581 95051
rect 296609 95023 296643 95051
rect 296671 95023 296719 95051
rect 296409 94989 296719 95023
rect 296409 94961 296457 94989
rect 296485 94961 296519 94989
rect 296547 94961 296581 94989
rect 296609 94961 296643 94989
rect 296671 94961 296719 94989
rect 296409 86175 296719 94961
rect 296409 86147 296457 86175
rect 296485 86147 296519 86175
rect 296547 86147 296581 86175
rect 296609 86147 296643 86175
rect 296671 86147 296719 86175
rect 296409 86113 296719 86147
rect 296409 86085 296457 86113
rect 296485 86085 296519 86113
rect 296547 86085 296581 86113
rect 296609 86085 296643 86113
rect 296671 86085 296719 86113
rect 296409 86051 296719 86085
rect 296409 86023 296457 86051
rect 296485 86023 296519 86051
rect 296547 86023 296581 86051
rect 296609 86023 296643 86051
rect 296671 86023 296719 86051
rect 296409 85989 296719 86023
rect 296409 85961 296457 85989
rect 296485 85961 296519 85989
rect 296547 85961 296581 85989
rect 296609 85961 296643 85989
rect 296671 85961 296719 85989
rect 296409 77175 296719 85961
rect 296409 77147 296457 77175
rect 296485 77147 296519 77175
rect 296547 77147 296581 77175
rect 296609 77147 296643 77175
rect 296671 77147 296719 77175
rect 296409 77113 296719 77147
rect 296409 77085 296457 77113
rect 296485 77085 296519 77113
rect 296547 77085 296581 77113
rect 296609 77085 296643 77113
rect 296671 77085 296719 77113
rect 296409 77051 296719 77085
rect 296409 77023 296457 77051
rect 296485 77023 296519 77051
rect 296547 77023 296581 77051
rect 296609 77023 296643 77051
rect 296671 77023 296719 77051
rect 296409 76989 296719 77023
rect 296409 76961 296457 76989
rect 296485 76961 296519 76989
rect 296547 76961 296581 76989
rect 296609 76961 296643 76989
rect 296671 76961 296719 76989
rect 296409 68175 296719 76961
rect 296409 68147 296457 68175
rect 296485 68147 296519 68175
rect 296547 68147 296581 68175
rect 296609 68147 296643 68175
rect 296671 68147 296719 68175
rect 296409 68113 296719 68147
rect 296409 68085 296457 68113
rect 296485 68085 296519 68113
rect 296547 68085 296581 68113
rect 296609 68085 296643 68113
rect 296671 68085 296719 68113
rect 296409 68051 296719 68085
rect 296409 68023 296457 68051
rect 296485 68023 296519 68051
rect 296547 68023 296581 68051
rect 296609 68023 296643 68051
rect 296671 68023 296719 68051
rect 296409 67989 296719 68023
rect 296409 67961 296457 67989
rect 296485 67961 296519 67989
rect 296547 67961 296581 67989
rect 296609 67961 296643 67989
rect 296671 67961 296719 67989
rect 296409 59175 296719 67961
rect 296409 59147 296457 59175
rect 296485 59147 296519 59175
rect 296547 59147 296581 59175
rect 296609 59147 296643 59175
rect 296671 59147 296719 59175
rect 296409 59113 296719 59147
rect 296409 59085 296457 59113
rect 296485 59085 296519 59113
rect 296547 59085 296581 59113
rect 296609 59085 296643 59113
rect 296671 59085 296719 59113
rect 296409 59051 296719 59085
rect 296409 59023 296457 59051
rect 296485 59023 296519 59051
rect 296547 59023 296581 59051
rect 296609 59023 296643 59051
rect 296671 59023 296719 59051
rect 296409 58989 296719 59023
rect 296409 58961 296457 58989
rect 296485 58961 296519 58989
rect 296547 58961 296581 58989
rect 296609 58961 296643 58989
rect 296671 58961 296719 58989
rect 294549 56147 294597 56175
rect 294625 56147 294659 56175
rect 294687 56147 294721 56175
rect 294749 56147 294783 56175
rect 294811 56147 294859 56175
rect 294549 56113 294859 56147
rect 294549 56085 294597 56113
rect 294625 56085 294659 56113
rect 294687 56085 294721 56113
rect 294749 56085 294783 56113
rect 294811 56085 294859 56113
rect 294549 56051 294859 56085
rect 294549 56023 294597 56051
rect 294625 56023 294659 56051
rect 294687 56023 294721 56051
rect 294749 56023 294783 56051
rect 294811 56023 294859 56051
rect 294549 55989 294859 56023
rect 294549 55961 294597 55989
rect 294625 55961 294659 55989
rect 294687 55961 294721 55989
rect 294749 55961 294783 55989
rect 294811 55961 294859 55989
rect 281049 50147 281097 50175
rect 281125 50147 281159 50175
rect 281187 50147 281221 50175
rect 281249 50147 281283 50175
rect 281311 50147 281359 50175
rect 281049 50113 281359 50147
rect 281049 50085 281097 50113
rect 281125 50085 281159 50113
rect 281187 50085 281221 50113
rect 281249 50085 281283 50113
rect 281311 50085 281359 50113
rect 281049 50051 281359 50085
rect 281049 50023 281097 50051
rect 281125 50023 281159 50051
rect 281187 50023 281221 50051
rect 281249 50023 281283 50051
rect 281311 50023 281359 50051
rect 281049 49989 281359 50023
rect 281049 49961 281097 49989
rect 281125 49961 281159 49989
rect 281187 49961 281221 49989
rect 281249 49961 281283 49989
rect 281311 49961 281359 49989
rect 281049 41175 281359 49961
rect 293566 49490 293594 49495
rect 284704 47175 284864 47192
rect 284704 47147 284739 47175
rect 284767 47147 284801 47175
rect 284829 47147 284864 47175
rect 284704 47113 284864 47147
rect 284704 47085 284739 47113
rect 284767 47085 284801 47113
rect 284829 47085 284864 47113
rect 284704 47051 284864 47085
rect 284704 47023 284739 47051
rect 284767 47023 284801 47051
rect 284829 47023 284864 47051
rect 284704 46989 284864 47023
rect 284704 46961 284739 46989
rect 284767 46961 284801 46989
rect 284829 46961 284864 46989
rect 284704 46944 284864 46961
rect 293566 43218 293594 49462
rect 293566 43185 293594 43190
rect 294549 47175 294859 55961
rect 295246 56770 295274 56775
rect 295246 49938 295274 56742
rect 295246 49905 295274 49910
rect 296409 50175 296719 58961
rect 296409 50147 296457 50175
rect 296485 50147 296519 50175
rect 296547 50147 296581 50175
rect 296609 50147 296643 50175
rect 296671 50147 296719 50175
rect 296409 50113 296719 50147
rect 296409 50085 296457 50113
rect 296485 50085 296519 50113
rect 296547 50085 296581 50113
rect 296609 50085 296643 50113
rect 296671 50085 296719 50113
rect 296409 50051 296719 50085
rect 296409 50023 296457 50051
rect 296485 50023 296519 50051
rect 296547 50023 296581 50051
rect 296609 50023 296643 50051
rect 296671 50023 296719 50051
rect 296409 49989 296719 50023
rect 296409 49961 296457 49989
rect 296485 49961 296519 49989
rect 296547 49961 296581 49989
rect 296609 49961 296643 49989
rect 296671 49961 296719 49989
rect 294549 47147 294597 47175
rect 294625 47147 294659 47175
rect 294687 47147 294721 47175
rect 294749 47147 294783 47175
rect 294811 47147 294859 47175
rect 294549 47113 294859 47147
rect 294549 47085 294597 47113
rect 294625 47085 294659 47113
rect 294687 47085 294721 47113
rect 294749 47085 294783 47113
rect 294811 47085 294859 47113
rect 294549 47051 294859 47085
rect 294549 47023 294597 47051
rect 294625 47023 294659 47051
rect 294687 47023 294721 47051
rect 294749 47023 294783 47051
rect 294811 47023 294859 47051
rect 294549 46989 294859 47023
rect 294549 46961 294597 46989
rect 294625 46961 294659 46989
rect 294687 46961 294721 46989
rect 294749 46961 294783 46989
rect 294811 46961 294859 46989
rect 281049 41147 281097 41175
rect 281125 41147 281159 41175
rect 281187 41147 281221 41175
rect 281249 41147 281283 41175
rect 281311 41147 281359 41175
rect 281049 41113 281359 41147
rect 281049 41085 281097 41113
rect 281125 41085 281159 41113
rect 281187 41085 281221 41113
rect 281249 41085 281283 41113
rect 281311 41085 281359 41113
rect 281049 41051 281359 41085
rect 281049 41023 281097 41051
rect 281125 41023 281159 41051
rect 281187 41023 281221 41051
rect 281249 41023 281283 41051
rect 281311 41023 281359 41051
rect 281049 40989 281359 41023
rect 281049 40961 281097 40989
rect 281125 40961 281159 40989
rect 281187 40961 281221 40989
rect 281249 40961 281283 40989
rect 281311 40961 281359 40989
rect 281049 32175 281359 40961
rect 293566 42210 293594 42215
rect 284704 38175 284864 38192
rect 284704 38147 284739 38175
rect 284767 38147 284801 38175
rect 284829 38147 284864 38175
rect 284704 38113 284864 38147
rect 284704 38085 284739 38113
rect 284767 38085 284801 38113
rect 284829 38085 284864 38113
rect 284704 38051 284864 38085
rect 284704 38023 284739 38051
rect 284767 38023 284801 38051
rect 284829 38023 284864 38051
rect 284704 37989 284864 38023
rect 284704 37961 284739 37989
rect 284767 37961 284801 37989
rect 284829 37961 284864 37989
rect 284704 37944 284864 37961
rect 293566 36610 293594 42182
rect 293566 36577 293594 36582
rect 294549 38175 294859 46961
rect 294549 38147 294597 38175
rect 294625 38147 294659 38175
rect 294687 38147 294721 38175
rect 294749 38147 294783 38175
rect 294811 38147 294859 38175
rect 294549 38113 294859 38147
rect 294549 38085 294597 38113
rect 294625 38085 294659 38113
rect 294687 38085 294721 38113
rect 294749 38085 294783 38113
rect 294811 38085 294859 38113
rect 294549 38051 294859 38085
rect 294549 38023 294597 38051
rect 294625 38023 294659 38051
rect 294687 38023 294721 38051
rect 294749 38023 294783 38051
rect 294811 38023 294859 38051
rect 294549 37989 294859 38023
rect 294549 37961 294597 37989
rect 294625 37961 294659 37989
rect 294687 37961 294721 37989
rect 294749 37961 294783 37989
rect 294811 37961 294859 37989
rect 281049 32147 281097 32175
rect 281125 32147 281159 32175
rect 281187 32147 281221 32175
rect 281249 32147 281283 32175
rect 281311 32147 281359 32175
rect 281049 32113 281359 32147
rect 281049 32085 281097 32113
rect 281125 32085 281159 32113
rect 281187 32085 281221 32113
rect 281249 32085 281283 32113
rect 281311 32085 281359 32113
rect 281049 32051 281359 32085
rect 281049 32023 281097 32051
rect 281125 32023 281159 32051
rect 281187 32023 281221 32051
rect 281249 32023 281283 32051
rect 281311 32023 281359 32051
rect 281049 31989 281359 32023
rect 281049 31961 281097 31989
rect 281125 31961 281159 31989
rect 281187 31961 281221 31989
rect 281249 31961 281283 31989
rect 281311 31961 281359 31989
rect 281049 23175 281359 31961
rect 293174 34930 293202 34935
rect 293174 30002 293202 34902
rect 293174 29969 293202 29974
rect 284704 29175 284864 29192
rect 284704 29147 284739 29175
rect 284767 29147 284801 29175
rect 284829 29147 284864 29175
rect 284704 29113 284864 29147
rect 284704 29085 284739 29113
rect 284767 29085 284801 29113
rect 284829 29085 284864 29113
rect 284704 29051 284864 29085
rect 284704 29023 284739 29051
rect 284767 29023 284801 29051
rect 284829 29023 284864 29051
rect 284704 28989 284864 29023
rect 284704 28961 284739 28989
rect 284767 28961 284801 28989
rect 284829 28961 284864 28989
rect 284704 28944 284864 28961
rect 294549 29175 294859 37961
rect 294549 29147 294597 29175
rect 294625 29147 294659 29175
rect 294687 29147 294721 29175
rect 294749 29147 294783 29175
rect 294811 29147 294859 29175
rect 294549 29113 294859 29147
rect 294549 29085 294597 29113
rect 294625 29085 294659 29113
rect 294687 29085 294721 29113
rect 294749 29085 294783 29113
rect 294811 29085 294859 29113
rect 294549 29051 294859 29085
rect 294549 29023 294597 29051
rect 294625 29023 294659 29051
rect 294687 29023 294721 29051
rect 294749 29023 294783 29051
rect 294811 29023 294859 29051
rect 294549 28989 294859 29023
rect 294549 28961 294597 28989
rect 294625 28961 294659 28989
rect 294687 28961 294721 28989
rect 294749 28961 294783 28989
rect 294811 28961 294859 28989
rect 293566 27650 293594 27655
rect 293566 23394 293594 27622
rect 293566 23361 293594 23366
rect 281049 23147 281097 23175
rect 281125 23147 281159 23175
rect 281187 23147 281221 23175
rect 281249 23147 281283 23175
rect 281311 23147 281359 23175
rect 281049 23113 281359 23147
rect 281049 23085 281097 23113
rect 281125 23085 281159 23113
rect 281187 23085 281221 23113
rect 281249 23085 281283 23113
rect 281311 23085 281359 23113
rect 281049 23051 281359 23085
rect 281049 23023 281097 23051
rect 281125 23023 281159 23051
rect 281187 23023 281221 23051
rect 281249 23023 281283 23051
rect 281311 23023 281359 23051
rect 281049 22989 281359 23023
rect 281049 22961 281097 22989
rect 281125 22961 281159 22989
rect 281187 22961 281221 22989
rect 281249 22961 281283 22989
rect 281311 22961 281359 22989
rect 281049 14175 281359 22961
rect 293566 20370 293594 20375
rect 284704 20175 284864 20192
rect 284704 20147 284739 20175
rect 284767 20147 284801 20175
rect 284829 20147 284864 20175
rect 284704 20113 284864 20147
rect 284704 20085 284739 20113
rect 284767 20085 284801 20113
rect 284829 20085 284864 20113
rect 284704 20051 284864 20085
rect 284704 20023 284739 20051
rect 284767 20023 284801 20051
rect 284829 20023 284864 20051
rect 284704 19989 284864 20023
rect 284704 19961 284739 19989
rect 284767 19961 284801 19989
rect 284829 19961 284864 19989
rect 284704 19944 284864 19961
rect 293566 16842 293594 20342
rect 293566 16809 293594 16814
rect 294549 20175 294859 28961
rect 294549 20147 294597 20175
rect 294625 20147 294659 20175
rect 294687 20147 294721 20175
rect 294749 20147 294783 20175
rect 294811 20147 294859 20175
rect 294549 20113 294859 20147
rect 294549 20085 294597 20113
rect 294625 20085 294659 20113
rect 294687 20085 294721 20113
rect 294749 20085 294783 20113
rect 294811 20085 294859 20113
rect 294549 20051 294859 20085
rect 294549 20023 294597 20051
rect 294625 20023 294659 20051
rect 294687 20023 294721 20051
rect 294749 20023 294783 20051
rect 294811 20023 294859 20051
rect 294549 19989 294859 20023
rect 294549 19961 294597 19989
rect 294625 19961 294659 19989
rect 294687 19961 294721 19989
rect 294749 19961 294783 19989
rect 294811 19961 294859 19989
rect 281049 14147 281097 14175
rect 281125 14147 281159 14175
rect 281187 14147 281221 14175
rect 281249 14147 281283 14175
rect 281311 14147 281359 14175
rect 281049 14113 281359 14147
rect 281049 14085 281097 14113
rect 281125 14085 281159 14113
rect 281187 14085 281221 14113
rect 281249 14085 281283 14113
rect 281311 14085 281359 14113
rect 281049 14051 281359 14085
rect 281049 14023 281097 14051
rect 281125 14023 281159 14051
rect 281187 14023 281221 14051
rect 281249 14023 281283 14051
rect 281311 14023 281359 14051
rect 281049 13989 281359 14023
rect 281049 13961 281097 13989
rect 281125 13961 281159 13989
rect 281187 13961 281221 13989
rect 281249 13961 281283 13989
rect 281311 13961 281359 13989
rect 281049 5175 281359 13961
rect 293566 13090 293594 13095
rect 284704 11175 284864 11192
rect 284704 11147 284739 11175
rect 284767 11147 284801 11175
rect 284829 11147 284864 11175
rect 284704 11113 284864 11147
rect 284704 11085 284739 11113
rect 284767 11085 284801 11113
rect 284829 11085 284864 11113
rect 284704 11051 284864 11085
rect 284704 11023 284739 11051
rect 284767 11023 284801 11051
rect 284829 11023 284864 11051
rect 284704 10989 284864 11023
rect 284704 10961 284739 10989
rect 284767 10961 284801 10989
rect 284829 10961 284864 10989
rect 284704 10944 284864 10961
rect 293566 10178 293594 13062
rect 293566 10145 293594 10150
rect 294549 11175 294859 19961
rect 294549 11147 294597 11175
rect 294625 11147 294659 11175
rect 294687 11147 294721 11175
rect 294749 11147 294783 11175
rect 294811 11147 294859 11175
rect 294549 11113 294859 11147
rect 294549 11085 294597 11113
rect 294625 11085 294659 11113
rect 294687 11085 294721 11113
rect 294749 11085 294783 11113
rect 294811 11085 294859 11113
rect 294549 11051 294859 11085
rect 294549 11023 294597 11051
rect 294625 11023 294659 11051
rect 294687 11023 294721 11051
rect 294749 11023 294783 11051
rect 294811 11023 294859 11051
rect 294549 10989 294859 11023
rect 294549 10961 294597 10989
rect 294625 10961 294659 10989
rect 294687 10961 294721 10989
rect 294749 10961 294783 10989
rect 294811 10961 294859 10989
rect 281049 5147 281097 5175
rect 281125 5147 281159 5175
rect 281187 5147 281221 5175
rect 281249 5147 281283 5175
rect 281311 5147 281359 5175
rect 281049 5113 281359 5147
rect 281049 5085 281097 5113
rect 281125 5085 281159 5113
rect 281187 5085 281221 5113
rect 281249 5085 281283 5113
rect 281311 5085 281359 5113
rect 281049 5051 281359 5085
rect 281049 5023 281097 5051
rect 281125 5023 281159 5051
rect 281187 5023 281221 5051
rect 281249 5023 281283 5051
rect 281311 5023 281359 5051
rect 281049 4989 281359 5023
rect 281049 4961 281097 4989
rect 281125 4961 281159 4989
rect 281187 4961 281221 4989
rect 281249 4961 281283 4989
rect 281311 4961 281359 4989
rect 281049 -560 281359 4961
rect 281049 -588 281097 -560
rect 281125 -588 281159 -560
rect 281187 -588 281221 -560
rect 281249 -588 281283 -560
rect 281311 -588 281359 -560
rect 281049 -622 281359 -588
rect 281049 -650 281097 -622
rect 281125 -650 281159 -622
rect 281187 -650 281221 -622
rect 281249 -650 281283 -622
rect 281311 -650 281359 -622
rect 281049 -684 281359 -650
rect 281049 -712 281097 -684
rect 281125 -712 281159 -684
rect 281187 -712 281221 -684
rect 281249 -712 281283 -684
rect 281311 -712 281359 -684
rect 281049 -746 281359 -712
rect 281049 -774 281097 -746
rect 281125 -774 281159 -746
rect 281187 -774 281221 -746
rect 281249 -774 281283 -746
rect 281311 -774 281359 -746
rect 281049 -822 281359 -774
rect 294549 2175 294859 10961
rect 296409 41175 296719 49961
rect 296409 41147 296457 41175
rect 296485 41147 296519 41175
rect 296547 41147 296581 41175
rect 296609 41147 296643 41175
rect 296671 41147 296719 41175
rect 296409 41113 296719 41147
rect 296409 41085 296457 41113
rect 296485 41085 296519 41113
rect 296547 41085 296581 41113
rect 296609 41085 296643 41113
rect 296671 41085 296719 41113
rect 296409 41051 296719 41085
rect 296409 41023 296457 41051
rect 296485 41023 296519 41051
rect 296547 41023 296581 41051
rect 296609 41023 296643 41051
rect 296671 41023 296719 41051
rect 296409 40989 296719 41023
rect 296409 40961 296457 40989
rect 296485 40961 296519 40989
rect 296547 40961 296581 40989
rect 296609 40961 296643 40989
rect 296671 40961 296719 40989
rect 296409 32175 296719 40961
rect 296409 32147 296457 32175
rect 296485 32147 296519 32175
rect 296547 32147 296581 32175
rect 296609 32147 296643 32175
rect 296671 32147 296719 32175
rect 296409 32113 296719 32147
rect 296409 32085 296457 32113
rect 296485 32085 296519 32113
rect 296547 32085 296581 32113
rect 296609 32085 296643 32113
rect 296671 32085 296719 32113
rect 296409 32051 296719 32085
rect 296409 32023 296457 32051
rect 296485 32023 296519 32051
rect 296547 32023 296581 32051
rect 296609 32023 296643 32051
rect 296671 32023 296719 32051
rect 296409 31989 296719 32023
rect 296409 31961 296457 31989
rect 296485 31961 296519 31989
rect 296547 31961 296581 31989
rect 296609 31961 296643 31989
rect 296671 31961 296719 31989
rect 296409 23175 296719 31961
rect 296409 23147 296457 23175
rect 296485 23147 296519 23175
rect 296547 23147 296581 23175
rect 296609 23147 296643 23175
rect 296671 23147 296719 23175
rect 296409 23113 296719 23147
rect 296409 23085 296457 23113
rect 296485 23085 296519 23113
rect 296547 23085 296581 23113
rect 296609 23085 296643 23113
rect 296671 23085 296719 23113
rect 296409 23051 296719 23085
rect 296409 23023 296457 23051
rect 296485 23023 296519 23051
rect 296547 23023 296581 23051
rect 296609 23023 296643 23051
rect 296671 23023 296719 23051
rect 296409 22989 296719 23023
rect 296409 22961 296457 22989
rect 296485 22961 296519 22989
rect 296547 22961 296581 22989
rect 296609 22961 296643 22989
rect 296671 22961 296719 22989
rect 296409 14175 296719 22961
rect 296409 14147 296457 14175
rect 296485 14147 296519 14175
rect 296547 14147 296581 14175
rect 296609 14147 296643 14175
rect 296671 14147 296719 14175
rect 296409 14113 296719 14147
rect 296409 14085 296457 14113
rect 296485 14085 296519 14113
rect 296547 14085 296581 14113
rect 296609 14085 296643 14113
rect 296671 14085 296719 14113
rect 296409 14051 296719 14085
rect 296409 14023 296457 14051
rect 296485 14023 296519 14051
rect 296547 14023 296581 14051
rect 296609 14023 296643 14051
rect 296671 14023 296719 14051
rect 296409 13989 296719 14023
rect 296409 13961 296457 13989
rect 296485 13961 296519 13989
rect 296547 13961 296581 13989
rect 296609 13961 296643 13989
rect 296671 13961 296719 13989
rect 295638 5810 295666 5815
rect 295638 3682 295666 5782
rect 295638 3649 295666 3654
rect 296409 5175 296719 13961
rect 296409 5147 296457 5175
rect 296485 5147 296519 5175
rect 296547 5147 296581 5175
rect 296609 5147 296643 5175
rect 296671 5147 296719 5175
rect 296409 5113 296719 5147
rect 296409 5085 296457 5113
rect 296485 5085 296519 5113
rect 296547 5085 296581 5113
rect 296609 5085 296643 5113
rect 296671 5085 296719 5113
rect 296409 5051 296719 5085
rect 296409 5023 296457 5051
rect 296485 5023 296519 5051
rect 296547 5023 296581 5051
rect 296609 5023 296643 5051
rect 296671 5023 296719 5051
rect 296409 4989 296719 5023
rect 296409 4961 296457 4989
rect 296485 4961 296519 4989
rect 296547 4961 296581 4989
rect 296609 4961 296643 4989
rect 296671 4961 296719 4989
rect 294549 2147 294597 2175
rect 294625 2147 294659 2175
rect 294687 2147 294721 2175
rect 294749 2147 294783 2175
rect 294811 2147 294859 2175
rect 294549 2113 294859 2147
rect 294549 2085 294597 2113
rect 294625 2085 294659 2113
rect 294687 2085 294721 2113
rect 294749 2085 294783 2113
rect 294811 2085 294859 2113
rect 294549 2051 294859 2085
rect 294549 2023 294597 2051
rect 294625 2023 294659 2051
rect 294687 2023 294721 2051
rect 294749 2023 294783 2051
rect 294811 2023 294859 2051
rect 294549 1989 294859 2023
rect 294549 1961 294597 1989
rect 294625 1961 294659 1989
rect 294687 1961 294721 1989
rect 294749 1961 294783 1989
rect 294811 1961 294859 1989
rect 294549 -80 294859 1961
rect 294549 -108 294597 -80
rect 294625 -108 294659 -80
rect 294687 -108 294721 -80
rect 294749 -108 294783 -80
rect 294811 -108 294859 -80
rect 294549 -142 294859 -108
rect 294549 -170 294597 -142
rect 294625 -170 294659 -142
rect 294687 -170 294721 -142
rect 294749 -170 294783 -142
rect 294811 -170 294859 -142
rect 294549 -204 294859 -170
rect 294549 -232 294597 -204
rect 294625 -232 294659 -204
rect 294687 -232 294721 -204
rect 294749 -232 294783 -204
rect 294811 -232 294859 -204
rect 294549 -266 294859 -232
rect 294549 -294 294597 -266
rect 294625 -294 294659 -266
rect 294687 -294 294721 -266
rect 294749 -294 294783 -266
rect 294811 -294 294859 -266
rect 294549 -822 294859 -294
rect 296409 -560 296719 4961
rect 298200 298606 298510 298654
rect 298200 298578 298248 298606
rect 298276 298578 298310 298606
rect 298338 298578 298372 298606
rect 298400 298578 298434 298606
rect 298462 298578 298510 298606
rect 298200 298544 298510 298578
rect 298200 298516 298248 298544
rect 298276 298516 298310 298544
rect 298338 298516 298372 298544
rect 298400 298516 298434 298544
rect 298462 298516 298510 298544
rect 298200 298482 298510 298516
rect 298200 298454 298248 298482
rect 298276 298454 298310 298482
rect 298338 298454 298372 298482
rect 298400 298454 298434 298482
rect 298462 298454 298510 298482
rect 298200 298420 298510 298454
rect 298200 298392 298248 298420
rect 298276 298392 298310 298420
rect 298338 298392 298372 298420
rect 298400 298392 298434 298420
rect 298462 298392 298510 298420
rect 298200 290175 298510 298392
rect 298200 290147 298248 290175
rect 298276 290147 298310 290175
rect 298338 290147 298372 290175
rect 298400 290147 298434 290175
rect 298462 290147 298510 290175
rect 298200 290113 298510 290147
rect 298200 290085 298248 290113
rect 298276 290085 298310 290113
rect 298338 290085 298372 290113
rect 298400 290085 298434 290113
rect 298462 290085 298510 290113
rect 298200 290051 298510 290085
rect 298200 290023 298248 290051
rect 298276 290023 298310 290051
rect 298338 290023 298372 290051
rect 298400 290023 298434 290051
rect 298462 290023 298510 290051
rect 298200 289989 298510 290023
rect 298200 289961 298248 289989
rect 298276 289961 298310 289989
rect 298338 289961 298372 289989
rect 298400 289961 298434 289989
rect 298462 289961 298510 289989
rect 298200 281175 298510 289961
rect 298200 281147 298248 281175
rect 298276 281147 298310 281175
rect 298338 281147 298372 281175
rect 298400 281147 298434 281175
rect 298462 281147 298510 281175
rect 298200 281113 298510 281147
rect 298200 281085 298248 281113
rect 298276 281085 298310 281113
rect 298338 281085 298372 281113
rect 298400 281085 298434 281113
rect 298462 281085 298510 281113
rect 298200 281051 298510 281085
rect 298200 281023 298248 281051
rect 298276 281023 298310 281051
rect 298338 281023 298372 281051
rect 298400 281023 298434 281051
rect 298462 281023 298510 281051
rect 298200 280989 298510 281023
rect 298200 280961 298248 280989
rect 298276 280961 298310 280989
rect 298338 280961 298372 280989
rect 298400 280961 298434 280989
rect 298462 280961 298510 280989
rect 298200 272175 298510 280961
rect 298200 272147 298248 272175
rect 298276 272147 298310 272175
rect 298338 272147 298372 272175
rect 298400 272147 298434 272175
rect 298462 272147 298510 272175
rect 298200 272113 298510 272147
rect 298200 272085 298248 272113
rect 298276 272085 298310 272113
rect 298338 272085 298372 272113
rect 298400 272085 298434 272113
rect 298462 272085 298510 272113
rect 298200 272051 298510 272085
rect 298200 272023 298248 272051
rect 298276 272023 298310 272051
rect 298338 272023 298372 272051
rect 298400 272023 298434 272051
rect 298462 272023 298510 272051
rect 298200 271989 298510 272023
rect 298200 271961 298248 271989
rect 298276 271961 298310 271989
rect 298338 271961 298372 271989
rect 298400 271961 298434 271989
rect 298462 271961 298510 271989
rect 298200 263175 298510 271961
rect 298200 263147 298248 263175
rect 298276 263147 298310 263175
rect 298338 263147 298372 263175
rect 298400 263147 298434 263175
rect 298462 263147 298510 263175
rect 298200 263113 298510 263147
rect 298200 263085 298248 263113
rect 298276 263085 298310 263113
rect 298338 263085 298372 263113
rect 298400 263085 298434 263113
rect 298462 263085 298510 263113
rect 298200 263051 298510 263085
rect 298200 263023 298248 263051
rect 298276 263023 298310 263051
rect 298338 263023 298372 263051
rect 298400 263023 298434 263051
rect 298462 263023 298510 263051
rect 298200 262989 298510 263023
rect 298200 262961 298248 262989
rect 298276 262961 298310 262989
rect 298338 262961 298372 262989
rect 298400 262961 298434 262989
rect 298462 262961 298510 262989
rect 298200 254175 298510 262961
rect 298200 254147 298248 254175
rect 298276 254147 298310 254175
rect 298338 254147 298372 254175
rect 298400 254147 298434 254175
rect 298462 254147 298510 254175
rect 298200 254113 298510 254147
rect 298200 254085 298248 254113
rect 298276 254085 298310 254113
rect 298338 254085 298372 254113
rect 298400 254085 298434 254113
rect 298462 254085 298510 254113
rect 298200 254051 298510 254085
rect 298200 254023 298248 254051
rect 298276 254023 298310 254051
rect 298338 254023 298372 254051
rect 298400 254023 298434 254051
rect 298462 254023 298510 254051
rect 298200 253989 298510 254023
rect 298200 253961 298248 253989
rect 298276 253961 298310 253989
rect 298338 253961 298372 253989
rect 298400 253961 298434 253989
rect 298462 253961 298510 253989
rect 298200 245175 298510 253961
rect 298200 245147 298248 245175
rect 298276 245147 298310 245175
rect 298338 245147 298372 245175
rect 298400 245147 298434 245175
rect 298462 245147 298510 245175
rect 298200 245113 298510 245147
rect 298200 245085 298248 245113
rect 298276 245085 298310 245113
rect 298338 245085 298372 245113
rect 298400 245085 298434 245113
rect 298462 245085 298510 245113
rect 298200 245051 298510 245085
rect 298200 245023 298248 245051
rect 298276 245023 298310 245051
rect 298338 245023 298372 245051
rect 298400 245023 298434 245051
rect 298462 245023 298510 245051
rect 298200 244989 298510 245023
rect 298200 244961 298248 244989
rect 298276 244961 298310 244989
rect 298338 244961 298372 244989
rect 298400 244961 298434 244989
rect 298462 244961 298510 244989
rect 298200 236175 298510 244961
rect 298200 236147 298248 236175
rect 298276 236147 298310 236175
rect 298338 236147 298372 236175
rect 298400 236147 298434 236175
rect 298462 236147 298510 236175
rect 298200 236113 298510 236147
rect 298200 236085 298248 236113
rect 298276 236085 298310 236113
rect 298338 236085 298372 236113
rect 298400 236085 298434 236113
rect 298462 236085 298510 236113
rect 298200 236051 298510 236085
rect 298200 236023 298248 236051
rect 298276 236023 298310 236051
rect 298338 236023 298372 236051
rect 298400 236023 298434 236051
rect 298462 236023 298510 236051
rect 298200 235989 298510 236023
rect 298200 235961 298248 235989
rect 298276 235961 298310 235989
rect 298338 235961 298372 235989
rect 298400 235961 298434 235989
rect 298462 235961 298510 235989
rect 298200 227175 298510 235961
rect 298200 227147 298248 227175
rect 298276 227147 298310 227175
rect 298338 227147 298372 227175
rect 298400 227147 298434 227175
rect 298462 227147 298510 227175
rect 298200 227113 298510 227147
rect 298200 227085 298248 227113
rect 298276 227085 298310 227113
rect 298338 227085 298372 227113
rect 298400 227085 298434 227113
rect 298462 227085 298510 227113
rect 298200 227051 298510 227085
rect 298200 227023 298248 227051
rect 298276 227023 298310 227051
rect 298338 227023 298372 227051
rect 298400 227023 298434 227051
rect 298462 227023 298510 227051
rect 298200 226989 298510 227023
rect 298200 226961 298248 226989
rect 298276 226961 298310 226989
rect 298338 226961 298372 226989
rect 298400 226961 298434 226989
rect 298462 226961 298510 226989
rect 298200 218175 298510 226961
rect 298200 218147 298248 218175
rect 298276 218147 298310 218175
rect 298338 218147 298372 218175
rect 298400 218147 298434 218175
rect 298462 218147 298510 218175
rect 298200 218113 298510 218147
rect 298200 218085 298248 218113
rect 298276 218085 298310 218113
rect 298338 218085 298372 218113
rect 298400 218085 298434 218113
rect 298462 218085 298510 218113
rect 298200 218051 298510 218085
rect 298200 218023 298248 218051
rect 298276 218023 298310 218051
rect 298338 218023 298372 218051
rect 298400 218023 298434 218051
rect 298462 218023 298510 218051
rect 298200 217989 298510 218023
rect 298200 217961 298248 217989
rect 298276 217961 298310 217989
rect 298338 217961 298372 217989
rect 298400 217961 298434 217989
rect 298462 217961 298510 217989
rect 298200 209175 298510 217961
rect 298200 209147 298248 209175
rect 298276 209147 298310 209175
rect 298338 209147 298372 209175
rect 298400 209147 298434 209175
rect 298462 209147 298510 209175
rect 298200 209113 298510 209147
rect 298200 209085 298248 209113
rect 298276 209085 298310 209113
rect 298338 209085 298372 209113
rect 298400 209085 298434 209113
rect 298462 209085 298510 209113
rect 298200 209051 298510 209085
rect 298200 209023 298248 209051
rect 298276 209023 298310 209051
rect 298338 209023 298372 209051
rect 298400 209023 298434 209051
rect 298462 209023 298510 209051
rect 298200 208989 298510 209023
rect 298200 208961 298248 208989
rect 298276 208961 298310 208989
rect 298338 208961 298372 208989
rect 298400 208961 298434 208989
rect 298462 208961 298510 208989
rect 298200 200175 298510 208961
rect 298200 200147 298248 200175
rect 298276 200147 298310 200175
rect 298338 200147 298372 200175
rect 298400 200147 298434 200175
rect 298462 200147 298510 200175
rect 298200 200113 298510 200147
rect 298200 200085 298248 200113
rect 298276 200085 298310 200113
rect 298338 200085 298372 200113
rect 298400 200085 298434 200113
rect 298462 200085 298510 200113
rect 298200 200051 298510 200085
rect 298200 200023 298248 200051
rect 298276 200023 298310 200051
rect 298338 200023 298372 200051
rect 298400 200023 298434 200051
rect 298462 200023 298510 200051
rect 298200 199989 298510 200023
rect 298200 199961 298248 199989
rect 298276 199961 298310 199989
rect 298338 199961 298372 199989
rect 298400 199961 298434 199989
rect 298462 199961 298510 199989
rect 298200 191175 298510 199961
rect 298200 191147 298248 191175
rect 298276 191147 298310 191175
rect 298338 191147 298372 191175
rect 298400 191147 298434 191175
rect 298462 191147 298510 191175
rect 298200 191113 298510 191147
rect 298200 191085 298248 191113
rect 298276 191085 298310 191113
rect 298338 191085 298372 191113
rect 298400 191085 298434 191113
rect 298462 191085 298510 191113
rect 298200 191051 298510 191085
rect 298200 191023 298248 191051
rect 298276 191023 298310 191051
rect 298338 191023 298372 191051
rect 298400 191023 298434 191051
rect 298462 191023 298510 191051
rect 298200 190989 298510 191023
rect 298200 190961 298248 190989
rect 298276 190961 298310 190989
rect 298338 190961 298372 190989
rect 298400 190961 298434 190989
rect 298462 190961 298510 190989
rect 298200 182175 298510 190961
rect 298200 182147 298248 182175
rect 298276 182147 298310 182175
rect 298338 182147 298372 182175
rect 298400 182147 298434 182175
rect 298462 182147 298510 182175
rect 298200 182113 298510 182147
rect 298200 182085 298248 182113
rect 298276 182085 298310 182113
rect 298338 182085 298372 182113
rect 298400 182085 298434 182113
rect 298462 182085 298510 182113
rect 298200 182051 298510 182085
rect 298200 182023 298248 182051
rect 298276 182023 298310 182051
rect 298338 182023 298372 182051
rect 298400 182023 298434 182051
rect 298462 182023 298510 182051
rect 298200 181989 298510 182023
rect 298200 181961 298248 181989
rect 298276 181961 298310 181989
rect 298338 181961 298372 181989
rect 298400 181961 298434 181989
rect 298462 181961 298510 181989
rect 298200 173175 298510 181961
rect 298200 173147 298248 173175
rect 298276 173147 298310 173175
rect 298338 173147 298372 173175
rect 298400 173147 298434 173175
rect 298462 173147 298510 173175
rect 298200 173113 298510 173147
rect 298200 173085 298248 173113
rect 298276 173085 298310 173113
rect 298338 173085 298372 173113
rect 298400 173085 298434 173113
rect 298462 173085 298510 173113
rect 298200 173051 298510 173085
rect 298200 173023 298248 173051
rect 298276 173023 298310 173051
rect 298338 173023 298372 173051
rect 298400 173023 298434 173051
rect 298462 173023 298510 173051
rect 298200 172989 298510 173023
rect 298200 172961 298248 172989
rect 298276 172961 298310 172989
rect 298338 172961 298372 172989
rect 298400 172961 298434 172989
rect 298462 172961 298510 172989
rect 298200 164175 298510 172961
rect 298200 164147 298248 164175
rect 298276 164147 298310 164175
rect 298338 164147 298372 164175
rect 298400 164147 298434 164175
rect 298462 164147 298510 164175
rect 298200 164113 298510 164147
rect 298200 164085 298248 164113
rect 298276 164085 298310 164113
rect 298338 164085 298372 164113
rect 298400 164085 298434 164113
rect 298462 164085 298510 164113
rect 298200 164051 298510 164085
rect 298200 164023 298248 164051
rect 298276 164023 298310 164051
rect 298338 164023 298372 164051
rect 298400 164023 298434 164051
rect 298462 164023 298510 164051
rect 298200 163989 298510 164023
rect 298200 163961 298248 163989
rect 298276 163961 298310 163989
rect 298338 163961 298372 163989
rect 298400 163961 298434 163989
rect 298462 163961 298510 163989
rect 298200 155175 298510 163961
rect 298200 155147 298248 155175
rect 298276 155147 298310 155175
rect 298338 155147 298372 155175
rect 298400 155147 298434 155175
rect 298462 155147 298510 155175
rect 298200 155113 298510 155147
rect 298200 155085 298248 155113
rect 298276 155085 298310 155113
rect 298338 155085 298372 155113
rect 298400 155085 298434 155113
rect 298462 155085 298510 155113
rect 298200 155051 298510 155085
rect 298200 155023 298248 155051
rect 298276 155023 298310 155051
rect 298338 155023 298372 155051
rect 298400 155023 298434 155051
rect 298462 155023 298510 155051
rect 298200 154989 298510 155023
rect 298200 154961 298248 154989
rect 298276 154961 298310 154989
rect 298338 154961 298372 154989
rect 298400 154961 298434 154989
rect 298462 154961 298510 154989
rect 298200 146175 298510 154961
rect 298200 146147 298248 146175
rect 298276 146147 298310 146175
rect 298338 146147 298372 146175
rect 298400 146147 298434 146175
rect 298462 146147 298510 146175
rect 298200 146113 298510 146147
rect 298200 146085 298248 146113
rect 298276 146085 298310 146113
rect 298338 146085 298372 146113
rect 298400 146085 298434 146113
rect 298462 146085 298510 146113
rect 298200 146051 298510 146085
rect 298200 146023 298248 146051
rect 298276 146023 298310 146051
rect 298338 146023 298372 146051
rect 298400 146023 298434 146051
rect 298462 146023 298510 146051
rect 298200 145989 298510 146023
rect 298200 145961 298248 145989
rect 298276 145961 298310 145989
rect 298338 145961 298372 145989
rect 298400 145961 298434 145989
rect 298462 145961 298510 145989
rect 298200 137175 298510 145961
rect 298200 137147 298248 137175
rect 298276 137147 298310 137175
rect 298338 137147 298372 137175
rect 298400 137147 298434 137175
rect 298462 137147 298510 137175
rect 298200 137113 298510 137147
rect 298200 137085 298248 137113
rect 298276 137085 298310 137113
rect 298338 137085 298372 137113
rect 298400 137085 298434 137113
rect 298462 137085 298510 137113
rect 298200 137051 298510 137085
rect 298200 137023 298248 137051
rect 298276 137023 298310 137051
rect 298338 137023 298372 137051
rect 298400 137023 298434 137051
rect 298462 137023 298510 137051
rect 298200 136989 298510 137023
rect 298200 136961 298248 136989
rect 298276 136961 298310 136989
rect 298338 136961 298372 136989
rect 298400 136961 298434 136989
rect 298462 136961 298510 136989
rect 298200 128175 298510 136961
rect 298200 128147 298248 128175
rect 298276 128147 298310 128175
rect 298338 128147 298372 128175
rect 298400 128147 298434 128175
rect 298462 128147 298510 128175
rect 298200 128113 298510 128147
rect 298200 128085 298248 128113
rect 298276 128085 298310 128113
rect 298338 128085 298372 128113
rect 298400 128085 298434 128113
rect 298462 128085 298510 128113
rect 298200 128051 298510 128085
rect 298200 128023 298248 128051
rect 298276 128023 298310 128051
rect 298338 128023 298372 128051
rect 298400 128023 298434 128051
rect 298462 128023 298510 128051
rect 298200 127989 298510 128023
rect 298200 127961 298248 127989
rect 298276 127961 298310 127989
rect 298338 127961 298372 127989
rect 298400 127961 298434 127989
rect 298462 127961 298510 127989
rect 298200 119175 298510 127961
rect 298200 119147 298248 119175
rect 298276 119147 298310 119175
rect 298338 119147 298372 119175
rect 298400 119147 298434 119175
rect 298462 119147 298510 119175
rect 298200 119113 298510 119147
rect 298200 119085 298248 119113
rect 298276 119085 298310 119113
rect 298338 119085 298372 119113
rect 298400 119085 298434 119113
rect 298462 119085 298510 119113
rect 298200 119051 298510 119085
rect 298200 119023 298248 119051
rect 298276 119023 298310 119051
rect 298338 119023 298372 119051
rect 298400 119023 298434 119051
rect 298462 119023 298510 119051
rect 298200 118989 298510 119023
rect 298200 118961 298248 118989
rect 298276 118961 298310 118989
rect 298338 118961 298372 118989
rect 298400 118961 298434 118989
rect 298462 118961 298510 118989
rect 298200 110175 298510 118961
rect 298200 110147 298248 110175
rect 298276 110147 298310 110175
rect 298338 110147 298372 110175
rect 298400 110147 298434 110175
rect 298462 110147 298510 110175
rect 298200 110113 298510 110147
rect 298200 110085 298248 110113
rect 298276 110085 298310 110113
rect 298338 110085 298372 110113
rect 298400 110085 298434 110113
rect 298462 110085 298510 110113
rect 298200 110051 298510 110085
rect 298200 110023 298248 110051
rect 298276 110023 298310 110051
rect 298338 110023 298372 110051
rect 298400 110023 298434 110051
rect 298462 110023 298510 110051
rect 298200 109989 298510 110023
rect 298200 109961 298248 109989
rect 298276 109961 298310 109989
rect 298338 109961 298372 109989
rect 298400 109961 298434 109989
rect 298462 109961 298510 109989
rect 298200 101175 298510 109961
rect 298200 101147 298248 101175
rect 298276 101147 298310 101175
rect 298338 101147 298372 101175
rect 298400 101147 298434 101175
rect 298462 101147 298510 101175
rect 298200 101113 298510 101147
rect 298200 101085 298248 101113
rect 298276 101085 298310 101113
rect 298338 101085 298372 101113
rect 298400 101085 298434 101113
rect 298462 101085 298510 101113
rect 298200 101051 298510 101085
rect 298200 101023 298248 101051
rect 298276 101023 298310 101051
rect 298338 101023 298372 101051
rect 298400 101023 298434 101051
rect 298462 101023 298510 101051
rect 298200 100989 298510 101023
rect 298200 100961 298248 100989
rect 298276 100961 298310 100989
rect 298338 100961 298372 100989
rect 298400 100961 298434 100989
rect 298462 100961 298510 100989
rect 298200 92175 298510 100961
rect 298200 92147 298248 92175
rect 298276 92147 298310 92175
rect 298338 92147 298372 92175
rect 298400 92147 298434 92175
rect 298462 92147 298510 92175
rect 298200 92113 298510 92147
rect 298200 92085 298248 92113
rect 298276 92085 298310 92113
rect 298338 92085 298372 92113
rect 298400 92085 298434 92113
rect 298462 92085 298510 92113
rect 298200 92051 298510 92085
rect 298200 92023 298248 92051
rect 298276 92023 298310 92051
rect 298338 92023 298372 92051
rect 298400 92023 298434 92051
rect 298462 92023 298510 92051
rect 298200 91989 298510 92023
rect 298200 91961 298248 91989
rect 298276 91961 298310 91989
rect 298338 91961 298372 91989
rect 298400 91961 298434 91989
rect 298462 91961 298510 91989
rect 298200 83175 298510 91961
rect 298200 83147 298248 83175
rect 298276 83147 298310 83175
rect 298338 83147 298372 83175
rect 298400 83147 298434 83175
rect 298462 83147 298510 83175
rect 298200 83113 298510 83147
rect 298200 83085 298248 83113
rect 298276 83085 298310 83113
rect 298338 83085 298372 83113
rect 298400 83085 298434 83113
rect 298462 83085 298510 83113
rect 298200 83051 298510 83085
rect 298200 83023 298248 83051
rect 298276 83023 298310 83051
rect 298338 83023 298372 83051
rect 298400 83023 298434 83051
rect 298462 83023 298510 83051
rect 298200 82989 298510 83023
rect 298200 82961 298248 82989
rect 298276 82961 298310 82989
rect 298338 82961 298372 82989
rect 298400 82961 298434 82989
rect 298462 82961 298510 82989
rect 298200 74175 298510 82961
rect 298200 74147 298248 74175
rect 298276 74147 298310 74175
rect 298338 74147 298372 74175
rect 298400 74147 298434 74175
rect 298462 74147 298510 74175
rect 298200 74113 298510 74147
rect 298200 74085 298248 74113
rect 298276 74085 298310 74113
rect 298338 74085 298372 74113
rect 298400 74085 298434 74113
rect 298462 74085 298510 74113
rect 298200 74051 298510 74085
rect 298200 74023 298248 74051
rect 298276 74023 298310 74051
rect 298338 74023 298372 74051
rect 298400 74023 298434 74051
rect 298462 74023 298510 74051
rect 298200 73989 298510 74023
rect 298200 73961 298248 73989
rect 298276 73961 298310 73989
rect 298338 73961 298372 73989
rect 298400 73961 298434 73989
rect 298462 73961 298510 73989
rect 298200 65175 298510 73961
rect 298200 65147 298248 65175
rect 298276 65147 298310 65175
rect 298338 65147 298372 65175
rect 298400 65147 298434 65175
rect 298462 65147 298510 65175
rect 298200 65113 298510 65147
rect 298200 65085 298248 65113
rect 298276 65085 298310 65113
rect 298338 65085 298372 65113
rect 298400 65085 298434 65113
rect 298462 65085 298510 65113
rect 298200 65051 298510 65085
rect 298200 65023 298248 65051
rect 298276 65023 298310 65051
rect 298338 65023 298372 65051
rect 298400 65023 298434 65051
rect 298462 65023 298510 65051
rect 298200 64989 298510 65023
rect 298200 64961 298248 64989
rect 298276 64961 298310 64989
rect 298338 64961 298372 64989
rect 298400 64961 298434 64989
rect 298462 64961 298510 64989
rect 298200 56175 298510 64961
rect 298200 56147 298248 56175
rect 298276 56147 298310 56175
rect 298338 56147 298372 56175
rect 298400 56147 298434 56175
rect 298462 56147 298510 56175
rect 298200 56113 298510 56147
rect 298200 56085 298248 56113
rect 298276 56085 298310 56113
rect 298338 56085 298372 56113
rect 298400 56085 298434 56113
rect 298462 56085 298510 56113
rect 298200 56051 298510 56085
rect 298200 56023 298248 56051
rect 298276 56023 298310 56051
rect 298338 56023 298372 56051
rect 298400 56023 298434 56051
rect 298462 56023 298510 56051
rect 298200 55989 298510 56023
rect 298200 55961 298248 55989
rect 298276 55961 298310 55989
rect 298338 55961 298372 55989
rect 298400 55961 298434 55989
rect 298462 55961 298510 55989
rect 298200 47175 298510 55961
rect 298200 47147 298248 47175
rect 298276 47147 298310 47175
rect 298338 47147 298372 47175
rect 298400 47147 298434 47175
rect 298462 47147 298510 47175
rect 298200 47113 298510 47147
rect 298200 47085 298248 47113
rect 298276 47085 298310 47113
rect 298338 47085 298372 47113
rect 298400 47085 298434 47113
rect 298462 47085 298510 47113
rect 298200 47051 298510 47085
rect 298200 47023 298248 47051
rect 298276 47023 298310 47051
rect 298338 47023 298372 47051
rect 298400 47023 298434 47051
rect 298462 47023 298510 47051
rect 298200 46989 298510 47023
rect 298200 46961 298248 46989
rect 298276 46961 298310 46989
rect 298338 46961 298372 46989
rect 298400 46961 298434 46989
rect 298462 46961 298510 46989
rect 298200 38175 298510 46961
rect 298200 38147 298248 38175
rect 298276 38147 298310 38175
rect 298338 38147 298372 38175
rect 298400 38147 298434 38175
rect 298462 38147 298510 38175
rect 298200 38113 298510 38147
rect 298200 38085 298248 38113
rect 298276 38085 298310 38113
rect 298338 38085 298372 38113
rect 298400 38085 298434 38113
rect 298462 38085 298510 38113
rect 298200 38051 298510 38085
rect 298200 38023 298248 38051
rect 298276 38023 298310 38051
rect 298338 38023 298372 38051
rect 298400 38023 298434 38051
rect 298462 38023 298510 38051
rect 298200 37989 298510 38023
rect 298200 37961 298248 37989
rect 298276 37961 298310 37989
rect 298338 37961 298372 37989
rect 298400 37961 298434 37989
rect 298462 37961 298510 37989
rect 298200 29175 298510 37961
rect 298200 29147 298248 29175
rect 298276 29147 298310 29175
rect 298338 29147 298372 29175
rect 298400 29147 298434 29175
rect 298462 29147 298510 29175
rect 298200 29113 298510 29147
rect 298200 29085 298248 29113
rect 298276 29085 298310 29113
rect 298338 29085 298372 29113
rect 298400 29085 298434 29113
rect 298462 29085 298510 29113
rect 298200 29051 298510 29085
rect 298200 29023 298248 29051
rect 298276 29023 298310 29051
rect 298338 29023 298372 29051
rect 298400 29023 298434 29051
rect 298462 29023 298510 29051
rect 298200 28989 298510 29023
rect 298200 28961 298248 28989
rect 298276 28961 298310 28989
rect 298338 28961 298372 28989
rect 298400 28961 298434 28989
rect 298462 28961 298510 28989
rect 298200 20175 298510 28961
rect 298200 20147 298248 20175
rect 298276 20147 298310 20175
rect 298338 20147 298372 20175
rect 298400 20147 298434 20175
rect 298462 20147 298510 20175
rect 298200 20113 298510 20147
rect 298200 20085 298248 20113
rect 298276 20085 298310 20113
rect 298338 20085 298372 20113
rect 298400 20085 298434 20113
rect 298462 20085 298510 20113
rect 298200 20051 298510 20085
rect 298200 20023 298248 20051
rect 298276 20023 298310 20051
rect 298338 20023 298372 20051
rect 298400 20023 298434 20051
rect 298462 20023 298510 20051
rect 298200 19989 298510 20023
rect 298200 19961 298248 19989
rect 298276 19961 298310 19989
rect 298338 19961 298372 19989
rect 298400 19961 298434 19989
rect 298462 19961 298510 19989
rect 298200 11175 298510 19961
rect 298200 11147 298248 11175
rect 298276 11147 298310 11175
rect 298338 11147 298372 11175
rect 298400 11147 298434 11175
rect 298462 11147 298510 11175
rect 298200 11113 298510 11147
rect 298200 11085 298248 11113
rect 298276 11085 298310 11113
rect 298338 11085 298372 11113
rect 298400 11085 298434 11113
rect 298462 11085 298510 11113
rect 298200 11051 298510 11085
rect 298200 11023 298248 11051
rect 298276 11023 298310 11051
rect 298338 11023 298372 11051
rect 298400 11023 298434 11051
rect 298462 11023 298510 11051
rect 298200 10989 298510 11023
rect 298200 10961 298248 10989
rect 298276 10961 298310 10989
rect 298338 10961 298372 10989
rect 298400 10961 298434 10989
rect 298462 10961 298510 10989
rect 298200 2175 298510 10961
rect 298200 2147 298248 2175
rect 298276 2147 298310 2175
rect 298338 2147 298372 2175
rect 298400 2147 298434 2175
rect 298462 2147 298510 2175
rect 298200 2113 298510 2147
rect 298200 2085 298248 2113
rect 298276 2085 298310 2113
rect 298338 2085 298372 2113
rect 298400 2085 298434 2113
rect 298462 2085 298510 2113
rect 298200 2051 298510 2085
rect 298200 2023 298248 2051
rect 298276 2023 298310 2051
rect 298338 2023 298372 2051
rect 298400 2023 298434 2051
rect 298462 2023 298510 2051
rect 298200 1989 298510 2023
rect 298200 1961 298248 1989
rect 298276 1961 298310 1989
rect 298338 1961 298372 1989
rect 298400 1961 298434 1989
rect 298462 1961 298510 1989
rect 298200 -80 298510 1961
rect 298200 -108 298248 -80
rect 298276 -108 298310 -80
rect 298338 -108 298372 -80
rect 298400 -108 298434 -80
rect 298462 -108 298510 -80
rect 298200 -142 298510 -108
rect 298200 -170 298248 -142
rect 298276 -170 298310 -142
rect 298338 -170 298372 -142
rect 298400 -170 298434 -142
rect 298462 -170 298510 -142
rect 298200 -204 298510 -170
rect 298200 -232 298248 -204
rect 298276 -232 298310 -204
rect 298338 -232 298372 -204
rect 298400 -232 298434 -204
rect 298462 -232 298510 -204
rect 298200 -266 298510 -232
rect 298200 -294 298248 -266
rect 298276 -294 298310 -266
rect 298338 -294 298372 -266
rect 298400 -294 298434 -266
rect 298462 -294 298510 -266
rect 298200 -342 298510 -294
rect 298680 293175 298990 298872
rect 298680 293147 298728 293175
rect 298756 293147 298790 293175
rect 298818 293147 298852 293175
rect 298880 293147 298914 293175
rect 298942 293147 298990 293175
rect 298680 293113 298990 293147
rect 298680 293085 298728 293113
rect 298756 293085 298790 293113
rect 298818 293085 298852 293113
rect 298880 293085 298914 293113
rect 298942 293085 298990 293113
rect 298680 293051 298990 293085
rect 298680 293023 298728 293051
rect 298756 293023 298790 293051
rect 298818 293023 298852 293051
rect 298880 293023 298914 293051
rect 298942 293023 298990 293051
rect 298680 292989 298990 293023
rect 298680 292961 298728 292989
rect 298756 292961 298790 292989
rect 298818 292961 298852 292989
rect 298880 292961 298914 292989
rect 298942 292961 298990 292989
rect 298680 284175 298990 292961
rect 298680 284147 298728 284175
rect 298756 284147 298790 284175
rect 298818 284147 298852 284175
rect 298880 284147 298914 284175
rect 298942 284147 298990 284175
rect 298680 284113 298990 284147
rect 298680 284085 298728 284113
rect 298756 284085 298790 284113
rect 298818 284085 298852 284113
rect 298880 284085 298914 284113
rect 298942 284085 298990 284113
rect 298680 284051 298990 284085
rect 298680 284023 298728 284051
rect 298756 284023 298790 284051
rect 298818 284023 298852 284051
rect 298880 284023 298914 284051
rect 298942 284023 298990 284051
rect 298680 283989 298990 284023
rect 298680 283961 298728 283989
rect 298756 283961 298790 283989
rect 298818 283961 298852 283989
rect 298880 283961 298914 283989
rect 298942 283961 298990 283989
rect 298680 275175 298990 283961
rect 298680 275147 298728 275175
rect 298756 275147 298790 275175
rect 298818 275147 298852 275175
rect 298880 275147 298914 275175
rect 298942 275147 298990 275175
rect 298680 275113 298990 275147
rect 298680 275085 298728 275113
rect 298756 275085 298790 275113
rect 298818 275085 298852 275113
rect 298880 275085 298914 275113
rect 298942 275085 298990 275113
rect 298680 275051 298990 275085
rect 298680 275023 298728 275051
rect 298756 275023 298790 275051
rect 298818 275023 298852 275051
rect 298880 275023 298914 275051
rect 298942 275023 298990 275051
rect 298680 274989 298990 275023
rect 298680 274961 298728 274989
rect 298756 274961 298790 274989
rect 298818 274961 298852 274989
rect 298880 274961 298914 274989
rect 298942 274961 298990 274989
rect 298680 266175 298990 274961
rect 298680 266147 298728 266175
rect 298756 266147 298790 266175
rect 298818 266147 298852 266175
rect 298880 266147 298914 266175
rect 298942 266147 298990 266175
rect 298680 266113 298990 266147
rect 298680 266085 298728 266113
rect 298756 266085 298790 266113
rect 298818 266085 298852 266113
rect 298880 266085 298914 266113
rect 298942 266085 298990 266113
rect 298680 266051 298990 266085
rect 298680 266023 298728 266051
rect 298756 266023 298790 266051
rect 298818 266023 298852 266051
rect 298880 266023 298914 266051
rect 298942 266023 298990 266051
rect 298680 265989 298990 266023
rect 298680 265961 298728 265989
rect 298756 265961 298790 265989
rect 298818 265961 298852 265989
rect 298880 265961 298914 265989
rect 298942 265961 298990 265989
rect 298680 257175 298990 265961
rect 298680 257147 298728 257175
rect 298756 257147 298790 257175
rect 298818 257147 298852 257175
rect 298880 257147 298914 257175
rect 298942 257147 298990 257175
rect 298680 257113 298990 257147
rect 298680 257085 298728 257113
rect 298756 257085 298790 257113
rect 298818 257085 298852 257113
rect 298880 257085 298914 257113
rect 298942 257085 298990 257113
rect 298680 257051 298990 257085
rect 298680 257023 298728 257051
rect 298756 257023 298790 257051
rect 298818 257023 298852 257051
rect 298880 257023 298914 257051
rect 298942 257023 298990 257051
rect 298680 256989 298990 257023
rect 298680 256961 298728 256989
rect 298756 256961 298790 256989
rect 298818 256961 298852 256989
rect 298880 256961 298914 256989
rect 298942 256961 298990 256989
rect 298680 248175 298990 256961
rect 298680 248147 298728 248175
rect 298756 248147 298790 248175
rect 298818 248147 298852 248175
rect 298880 248147 298914 248175
rect 298942 248147 298990 248175
rect 298680 248113 298990 248147
rect 298680 248085 298728 248113
rect 298756 248085 298790 248113
rect 298818 248085 298852 248113
rect 298880 248085 298914 248113
rect 298942 248085 298990 248113
rect 298680 248051 298990 248085
rect 298680 248023 298728 248051
rect 298756 248023 298790 248051
rect 298818 248023 298852 248051
rect 298880 248023 298914 248051
rect 298942 248023 298990 248051
rect 298680 247989 298990 248023
rect 298680 247961 298728 247989
rect 298756 247961 298790 247989
rect 298818 247961 298852 247989
rect 298880 247961 298914 247989
rect 298942 247961 298990 247989
rect 298680 239175 298990 247961
rect 298680 239147 298728 239175
rect 298756 239147 298790 239175
rect 298818 239147 298852 239175
rect 298880 239147 298914 239175
rect 298942 239147 298990 239175
rect 298680 239113 298990 239147
rect 298680 239085 298728 239113
rect 298756 239085 298790 239113
rect 298818 239085 298852 239113
rect 298880 239085 298914 239113
rect 298942 239085 298990 239113
rect 298680 239051 298990 239085
rect 298680 239023 298728 239051
rect 298756 239023 298790 239051
rect 298818 239023 298852 239051
rect 298880 239023 298914 239051
rect 298942 239023 298990 239051
rect 298680 238989 298990 239023
rect 298680 238961 298728 238989
rect 298756 238961 298790 238989
rect 298818 238961 298852 238989
rect 298880 238961 298914 238989
rect 298942 238961 298990 238989
rect 298680 230175 298990 238961
rect 298680 230147 298728 230175
rect 298756 230147 298790 230175
rect 298818 230147 298852 230175
rect 298880 230147 298914 230175
rect 298942 230147 298990 230175
rect 298680 230113 298990 230147
rect 298680 230085 298728 230113
rect 298756 230085 298790 230113
rect 298818 230085 298852 230113
rect 298880 230085 298914 230113
rect 298942 230085 298990 230113
rect 298680 230051 298990 230085
rect 298680 230023 298728 230051
rect 298756 230023 298790 230051
rect 298818 230023 298852 230051
rect 298880 230023 298914 230051
rect 298942 230023 298990 230051
rect 298680 229989 298990 230023
rect 298680 229961 298728 229989
rect 298756 229961 298790 229989
rect 298818 229961 298852 229989
rect 298880 229961 298914 229989
rect 298942 229961 298990 229989
rect 298680 221175 298990 229961
rect 298680 221147 298728 221175
rect 298756 221147 298790 221175
rect 298818 221147 298852 221175
rect 298880 221147 298914 221175
rect 298942 221147 298990 221175
rect 298680 221113 298990 221147
rect 298680 221085 298728 221113
rect 298756 221085 298790 221113
rect 298818 221085 298852 221113
rect 298880 221085 298914 221113
rect 298942 221085 298990 221113
rect 298680 221051 298990 221085
rect 298680 221023 298728 221051
rect 298756 221023 298790 221051
rect 298818 221023 298852 221051
rect 298880 221023 298914 221051
rect 298942 221023 298990 221051
rect 298680 220989 298990 221023
rect 298680 220961 298728 220989
rect 298756 220961 298790 220989
rect 298818 220961 298852 220989
rect 298880 220961 298914 220989
rect 298942 220961 298990 220989
rect 298680 212175 298990 220961
rect 298680 212147 298728 212175
rect 298756 212147 298790 212175
rect 298818 212147 298852 212175
rect 298880 212147 298914 212175
rect 298942 212147 298990 212175
rect 298680 212113 298990 212147
rect 298680 212085 298728 212113
rect 298756 212085 298790 212113
rect 298818 212085 298852 212113
rect 298880 212085 298914 212113
rect 298942 212085 298990 212113
rect 298680 212051 298990 212085
rect 298680 212023 298728 212051
rect 298756 212023 298790 212051
rect 298818 212023 298852 212051
rect 298880 212023 298914 212051
rect 298942 212023 298990 212051
rect 298680 211989 298990 212023
rect 298680 211961 298728 211989
rect 298756 211961 298790 211989
rect 298818 211961 298852 211989
rect 298880 211961 298914 211989
rect 298942 211961 298990 211989
rect 298680 203175 298990 211961
rect 298680 203147 298728 203175
rect 298756 203147 298790 203175
rect 298818 203147 298852 203175
rect 298880 203147 298914 203175
rect 298942 203147 298990 203175
rect 298680 203113 298990 203147
rect 298680 203085 298728 203113
rect 298756 203085 298790 203113
rect 298818 203085 298852 203113
rect 298880 203085 298914 203113
rect 298942 203085 298990 203113
rect 298680 203051 298990 203085
rect 298680 203023 298728 203051
rect 298756 203023 298790 203051
rect 298818 203023 298852 203051
rect 298880 203023 298914 203051
rect 298942 203023 298990 203051
rect 298680 202989 298990 203023
rect 298680 202961 298728 202989
rect 298756 202961 298790 202989
rect 298818 202961 298852 202989
rect 298880 202961 298914 202989
rect 298942 202961 298990 202989
rect 298680 194175 298990 202961
rect 298680 194147 298728 194175
rect 298756 194147 298790 194175
rect 298818 194147 298852 194175
rect 298880 194147 298914 194175
rect 298942 194147 298990 194175
rect 298680 194113 298990 194147
rect 298680 194085 298728 194113
rect 298756 194085 298790 194113
rect 298818 194085 298852 194113
rect 298880 194085 298914 194113
rect 298942 194085 298990 194113
rect 298680 194051 298990 194085
rect 298680 194023 298728 194051
rect 298756 194023 298790 194051
rect 298818 194023 298852 194051
rect 298880 194023 298914 194051
rect 298942 194023 298990 194051
rect 298680 193989 298990 194023
rect 298680 193961 298728 193989
rect 298756 193961 298790 193989
rect 298818 193961 298852 193989
rect 298880 193961 298914 193989
rect 298942 193961 298990 193989
rect 298680 185175 298990 193961
rect 298680 185147 298728 185175
rect 298756 185147 298790 185175
rect 298818 185147 298852 185175
rect 298880 185147 298914 185175
rect 298942 185147 298990 185175
rect 298680 185113 298990 185147
rect 298680 185085 298728 185113
rect 298756 185085 298790 185113
rect 298818 185085 298852 185113
rect 298880 185085 298914 185113
rect 298942 185085 298990 185113
rect 298680 185051 298990 185085
rect 298680 185023 298728 185051
rect 298756 185023 298790 185051
rect 298818 185023 298852 185051
rect 298880 185023 298914 185051
rect 298942 185023 298990 185051
rect 298680 184989 298990 185023
rect 298680 184961 298728 184989
rect 298756 184961 298790 184989
rect 298818 184961 298852 184989
rect 298880 184961 298914 184989
rect 298942 184961 298990 184989
rect 298680 176175 298990 184961
rect 298680 176147 298728 176175
rect 298756 176147 298790 176175
rect 298818 176147 298852 176175
rect 298880 176147 298914 176175
rect 298942 176147 298990 176175
rect 298680 176113 298990 176147
rect 298680 176085 298728 176113
rect 298756 176085 298790 176113
rect 298818 176085 298852 176113
rect 298880 176085 298914 176113
rect 298942 176085 298990 176113
rect 298680 176051 298990 176085
rect 298680 176023 298728 176051
rect 298756 176023 298790 176051
rect 298818 176023 298852 176051
rect 298880 176023 298914 176051
rect 298942 176023 298990 176051
rect 298680 175989 298990 176023
rect 298680 175961 298728 175989
rect 298756 175961 298790 175989
rect 298818 175961 298852 175989
rect 298880 175961 298914 175989
rect 298942 175961 298990 175989
rect 298680 167175 298990 175961
rect 298680 167147 298728 167175
rect 298756 167147 298790 167175
rect 298818 167147 298852 167175
rect 298880 167147 298914 167175
rect 298942 167147 298990 167175
rect 298680 167113 298990 167147
rect 298680 167085 298728 167113
rect 298756 167085 298790 167113
rect 298818 167085 298852 167113
rect 298880 167085 298914 167113
rect 298942 167085 298990 167113
rect 298680 167051 298990 167085
rect 298680 167023 298728 167051
rect 298756 167023 298790 167051
rect 298818 167023 298852 167051
rect 298880 167023 298914 167051
rect 298942 167023 298990 167051
rect 298680 166989 298990 167023
rect 298680 166961 298728 166989
rect 298756 166961 298790 166989
rect 298818 166961 298852 166989
rect 298880 166961 298914 166989
rect 298942 166961 298990 166989
rect 298680 158175 298990 166961
rect 298680 158147 298728 158175
rect 298756 158147 298790 158175
rect 298818 158147 298852 158175
rect 298880 158147 298914 158175
rect 298942 158147 298990 158175
rect 298680 158113 298990 158147
rect 298680 158085 298728 158113
rect 298756 158085 298790 158113
rect 298818 158085 298852 158113
rect 298880 158085 298914 158113
rect 298942 158085 298990 158113
rect 298680 158051 298990 158085
rect 298680 158023 298728 158051
rect 298756 158023 298790 158051
rect 298818 158023 298852 158051
rect 298880 158023 298914 158051
rect 298942 158023 298990 158051
rect 298680 157989 298990 158023
rect 298680 157961 298728 157989
rect 298756 157961 298790 157989
rect 298818 157961 298852 157989
rect 298880 157961 298914 157989
rect 298942 157961 298990 157989
rect 298680 149175 298990 157961
rect 298680 149147 298728 149175
rect 298756 149147 298790 149175
rect 298818 149147 298852 149175
rect 298880 149147 298914 149175
rect 298942 149147 298990 149175
rect 298680 149113 298990 149147
rect 298680 149085 298728 149113
rect 298756 149085 298790 149113
rect 298818 149085 298852 149113
rect 298880 149085 298914 149113
rect 298942 149085 298990 149113
rect 298680 149051 298990 149085
rect 298680 149023 298728 149051
rect 298756 149023 298790 149051
rect 298818 149023 298852 149051
rect 298880 149023 298914 149051
rect 298942 149023 298990 149051
rect 298680 148989 298990 149023
rect 298680 148961 298728 148989
rect 298756 148961 298790 148989
rect 298818 148961 298852 148989
rect 298880 148961 298914 148989
rect 298942 148961 298990 148989
rect 298680 140175 298990 148961
rect 298680 140147 298728 140175
rect 298756 140147 298790 140175
rect 298818 140147 298852 140175
rect 298880 140147 298914 140175
rect 298942 140147 298990 140175
rect 298680 140113 298990 140147
rect 298680 140085 298728 140113
rect 298756 140085 298790 140113
rect 298818 140085 298852 140113
rect 298880 140085 298914 140113
rect 298942 140085 298990 140113
rect 298680 140051 298990 140085
rect 298680 140023 298728 140051
rect 298756 140023 298790 140051
rect 298818 140023 298852 140051
rect 298880 140023 298914 140051
rect 298942 140023 298990 140051
rect 298680 139989 298990 140023
rect 298680 139961 298728 139989
rect 298756 139961 298790 139989
rect 298818 139961 298852 139989
rect 298880 139961 298914 139989
rect 298942 139961 298990 139989
rect 298680 131175 298990 139961
rect 298680 131147 298728 131175
rect 298756 131147 298790 131175
rect 298818 131147 298852 131175
rect 298880 131147 298914 131175
rect 298942 131147 298990 131175
rect 298680 131113 298990 131147
rect 298680 131085 298728 131113
rect 298756 131085 298790 131113
rect 298818 131085 298852 131113
rect 298880 131085 298914 131113
rect 298942 131085 298990 131113
rect 298680 131051 298990 131085
rect 298680 131023 298728 131051
rect 298756 131023 298790 131051
rect 298818 131023 298852 131051
rect 298880 131023 298914 131051
rect 298942 131023 298990 131051
rect 298680 130989 298990 131023
rect 298680 130961 298728 130989
rect 298756 130961 298790 130989
rect 298818 130961 298852 130989
rect 298880 130961 298914 130989
rect 298942 130961 298990 130989
rect 298680 122175 298990 130961
rect 298680 122147 298728 122175
rect 298756 122147 298790 122175
rect 298818 122147 298852 122175
rect 298880 122147 298914 122175
rect 298942 122147 298990 122175
rect 298680 122113 298990 122147
rect 298680 122085 298728 122113
rect 298756 122085 298790 122113
rect 298818 122085 298852 122113
rect 298880 122085 298914 122113
rect 298942 122085 298990 122113
rect 298680 122051 298990 122085
rect 298680 122023 298728 122051
rect 298756 122023 298790 122051
rect 298818 122023 298852 122051
rect 298880 122023 298914 122051
rect 298942 122023 298990 122051
rect 298680 121989 298990 122023
rect 298680 121961 298728 121989
rect 298756 121961 298790 121989
rect 298818 121961 298852 121989
rect 298880 121961 298914 121989
rect 298942 121961 298990 121989
rect 298680 113175 298990 121961
rect 298680 113147 298728 113175
rect 298756 113147 298790 113175
rect 298818 113147 298852 113175
rect 298880 113147 298914 113175
rect 298942 113147 298990 113175
rect 298680 113113 298990 113147
rect 298680 113085 298728 113113
rect 298756 113085 298790 113113
rect 298818 113085 298852 113113
rect 298880 113085 298914 113113
rect 298942 113085 298990 113113
rect 298680 113051 298990 113085
rect 298680 113023 298728 113051
rect 298756 113023 298790 113051
rect 298818 113023 298852 113051
rect 298880 113023 298914 113051
rect 298942 113023 298990 113051
rect 298680 112989 298990 113023
rect 298680 112961 298728 112989
rect 298756 112961 298790 112989
rect 298818 112961 298852 112989
rect 298880 112961 298914 112989
rect 298942 112961 298990 112989
rect 298680 104175 298990 112961
rect 298680 104147 298728 104175
rect 298756 104147 298790 104175
rect 298818 104147 298852 104175
rect 298880 104147 298914 104175
rect 298942 104147 298990 104175
rect 298680 104113 298990 104147
rect 298680 104085 298728 104113
rect 298756 104085 298790 104113
rect 298818 104085 298852 104113
rect 298880 104085 298914 104113
rect 298942 104085 298990 104113
rect 298680 104051 298990 104085
rect 298680 104023 298728 104051
rect 298756 104023 298790 104051
rect 298818 104023 298852 104051
rect 298880 104023 298914 104051
rect 298942 104023 298990 104051
rect 298680 103989 298990 104023
rect 298680 103961 298728 103989
rect 298756 103961 298790 103989
rect 298818 103961 298852 103989
rect 298880 103961 298914 103989
rect 298942 103961 298990 103989
rect 298680 95175 298990 103961
rect 298680 95147 298728 95175
rect 298756 95147 298790 95175
rect 298818 95147 298852 95175
rect 298880 95147 298914 95175
rect 298942 95147 298990 95175
rect 298680 95113 298990 95147
rect 298680 95085 298728 95113
rect 298756 95085 298790 95113
rect 298818 95085 298852 95113
rect 298880 95085 298914 95113
rect 298942 95085 298990 95113
rect 298680 95051 298990 95085
rect 298680 95023 298728 95051
rect 298756 95023 298790 95051
rect 298818 95023 298852 95051
rect 298880 95023 298914 95051
rect 298942 95023 298990 95051
rect 298680 94989 298990 95023
rect 298680 94961 298728 94989
rect 298756 94961 298790 94989
rect 298818 94961 298852 94989
rect 298880 94961 298914 94989
rect 298942 94961 298990 94989
rect 298680 86175 298990 94961
rect 298680 86147 298728 86175
rect 298756 86147 298790 86175
rect 298818 86147 298852 86175
rect 298880 86147 298914 86175
rect 298942 86147 298990 86175
rect 298680 86113 298990 86147
rect 298680 86085 298728 86113
rect 298756 86085 298790 86113
rect 298818 86085 298852 86113
rect 298880 86085 298914 86113
rect 298942 86085 298990 86113
rect 298680 86051 298990 86085
rect 298680 86023 298728 86051
rect 298756 86023 298790 86051
rect 298818 86023 298852 86051
rect 298880 86023 298914 86051
rect 298942 86023 298990 86051
rect 298680 85989 298990 86023
rect 298680 85961 298728 85989
rect 298756 85961 298790 85989
rect 298818 85961 298852 85989
rect 298880 85961 298914 85989
rect 298942 85961 298990 85989
rect 298680 77175 298990 85961
rect 298680 77147 298728 77175
rect 298756 77147 298790 77175
rect 298818 77147 298852 77175
rect 298880 77147 298914 77175
rect 298942 77147 298990 77175
rect 298680 77113 298990 77147
rect 298680 77085 298728 77113
rect 298756 77085 298790 77113
rect 298818 77085 298852 77113
rect 298880 77085 298914 77113
rect 298942 77085 298990 77113
rect 298680 77051 298990 77085
rect 298680 77023 298728 77051
rect 298756 77023 298790 77051
rect 298818 77023 298852 77051
rect 298880 77023 298914 77051
rect 298942 77023 298990 77051
rect 298680 76989 298990 77023
rect 298680 76961 298728 76989
rect 298756 76961 298790 76989
rect 298818 76961 298852 76989
rect 298880 76961 298914 76989
rect 298942 76961 298990 76989
rect 298680 68175 298990 76961
rect 298680 68147 298728 68175
rect 298756 68147 298790 68175
rect 298818 68147 298852 68175
rect 298880 68147 298914 68175
rect 298942 68147 298990 68175
rect 298680 68113 298990 68147
rect 298680 68085 298728 68113
rect 298756 68085 298790 68113
rect 298818 68085 298852 68113
rect 298880 68085 298914 68113
rect 298942 68085 298990 68113
rect 298680 68051 298990 68085
rect 298680 68023 298728 68051
rect 298756 68023 298790 68051
rect 298818 68023 298852 68051
rect 298880 68023 298914 68051
rect 298942 68023 298990 68051
rect 298680 67989 298990 68023
rect 298680 67961 298728 67989
rect 298756 67961 298790 67989
rect 298818 67961 298852 67989
rect 298880 67961 298914 67989
rect 298942 67961 298990 67989
rect 298680 59175 298990 67961
rect 298680 59147 298728 59175
rect 298756 59147 298790 59175
rect 298818 59147 298852 59175
rect 298880 59147 298914 59175
rect 298942 59147 298990 59175
rect 298680 59113 298990 59147
rect 298680 59085 298728 59113
rect 298756 59085 298790 59113
rect 298818 59085 298852 59113
rect 298880 59085 298914 59113
rect 298942 59085 298990 59113
rect 298680 59051 298990 59085
rect 298680 59023 298728 59051
rect 298756 59023 298790 59051
rect 298818 59023 298852 59051
rect 298880 59023 298914 59051
rect 298942 59023 298990 59051
rect 298680 58989 298990 59023
rect 298680 58961 298728 58989
rect 298756 58961 298790 58989
rect 298818 58961 298852 58989
rect 298880 58961 298914 58989
rect 298942 58961 298990 58989
rect 298680 50175 298990 58961
rect 298680 50147 298728 50175
rect 298756 50147 298790 50175
rect 298818 50147 298852 50175
rect 298880 50147 298914 50175
rect 298942 50147 298990 50175
rect 298680 50113 298990 50147
rect 298680 50085 298728 50113
rect 298756 50085 298790 50113
rect 298818 50085 298852 50113
rect 298880 50085 298914 50113
rect 298942 50085 298990 50113
rect 298680 50051 298990 50085
rect 298680 50023 298728 50051
rect 298756 50023 298790 50051
rect 298818 50023 298852 50051
rect 298880 50023 298914 50051
rect 298942 50023 298990 50051
rect 298680 49989 298990 50023
rect 298680 49961 298728 49989
rect 298756 49961 298790 49989
rect 298818 49961 298852 49989
rect 298880 49961 298914 49989
rect 298942 49961 298990 49989
rect 298680 41175 298990 49961
rect 298680 41147 298728 41175
rect 298756 41147 298790 41175
rect 298818 41147 298852 41175
rect 298880 41147 298914 41175
rect 298942 41147 298990 41175
rect 298680 41113 298990 41147
rect 298680 41085 298728 41113
rect 298756 41085 298790 41113
rect 298818 41085 298852 41113
rect 298880 41085 298914 41113
rect 298942 41085 298990 41113
rect 298680 41051 298990 41085
rect 298680 41023 298728 41051
rect 298756 41023 298790 41051
rect 298818 41023 298852 41051
rect 298880 41023 298914 41051
rect 298942 41023 298990 41051
rect 298680 40989 298990 41023
rect 298680 40961 298728 40989
rect 298756 40961 298790 40989
rect 298818 40961 298852 40989
rect 298880 40961 298914 40989
rect 298942 40961 298990 40989
rect 298680 32175 298990 40961
rect 298680 32147 298728 32175
rect 298756 32147 298790 32175
rect 298818 32147 298852 32175
rect 298880 32147 298914 32175
rect 298942 32147 298990 32175
rect 298680 32113 298990 32147
rect 298680 32085 298728 32113
rect 298756 32085 298790 32113
rect 298818 32085 298852 32113
rect 298880 32085 298914 32113
rect 298942 32085 298990 32113
rect 298680 32051 298990 32085
rect 298680 32023 298728 32051
rect 298756 32023 298790 32051
rect 298818 32023 298852 32051
rect 298880 32023 298914 32051
rect 298942 32023 298990 32051
rect 298680 31989 298990 32023
rect 298680 31961 298728 31989
rect 298756 31961 298790 31989
rect 298818 31961 298852 31989
rect 298880 31961 298914 31989
rect 298942 31961 298990 31989
rect 298680 23175 298990 31961
rect 298680 23147 298728 23175
rect 298756 23147 298790 23175
rect 298818 23147 298852 23175
rect 298880 23147 298914 23175
rect 298942 23147 298990 23175
rect 298680 23113 298990 23147
rect 298680 23085 298728 23113
rect 298756 23085 298790 23113
rect 298818 23085 298852 23113
rect 298880 23085 298914 23113
rect 298942 23085 298990 23113
rect 298680 23051 298990 23085
rect 298680 23023 298728 23051
rect 298756 23023 298790 23051
rect 298818 23023 298852 23051
rect 298880 23023 298914 23051
rect 298942 23023 298990 23051
rect 298680 22989 298990 23023
rect 298680 22961 298728 22989
rect 298756 22961 298790 22989
rect 298818 22961 298852 22989
rect 298880 22961 298914 22989
rect 298942 22961 298990 22989
rect 298680 14175 298990 22961
rect 298680 14147 298728 14175
rect 298756 14147 298790 14175
rect 298818 14147 298852 14175
rect 298880 14147 298914 14175
rect 298942 14147 298990 14175
rect 298680 14113 298990 14147
rect 298680 14085 298728 14113
rect 298756 14085 298790 14113
rect 298818 14085 298852 14113
rect 298880 14085 298914 14113
rect 298942 14085 298990 14113
rect 298680 14051 298990 14085
rect 298680 14023 298728 14051
rect 298756 14023 298790 14051
rect 298818 14023 298852 14051
rect 298880 14023 298914 14051
rect 298942 14023 298990 14051
rect 298680 13989 298990 14023
rect 298680 13961 298728 13989
rect 298756 13961 298790 13989
rect 298818 13961 298852 13989
rect 298880 13961 298914 13989
rect 298942 13961 298990 13989
rect 298680 5175 298990 13961
rect 298680 5147 298728 5175
rect 298756 5147 298790 5175
rect 298818 5147 298852 5175
rect 298880 5147 298914 5175
rect 298942 5147 298990 5175
rect 298680 5113 298990 5147
rect 298680 5085 298728 5113
rect 298756 5085 298790 5113
rect 298818 5085 298852 5113
rect 298880 5085 298914 5113
rect 298942 5085 298990 5113
rect 298680 5051 298990 5085
rect 298680 5023 298728 5051
rect 298756 5023 298790 5051
rect 298818 5023 298852 5051
rect 298880 5023 298914 5051
rect 298942 5023 298990 5051
rect 298680 4989 298990 5023
rect 298680 4961 298728 4989
rect 298756 4961 298790 4989
rect 298818 4961 298852 4989
rect 298880 4961 298914 4989
rect 298942 4961 298990 4989
rect 296409 -588 296457 -560
rect 296485 -588 296519 -560
rect 296547 -588 296581 -560
rect 296609 -588 296643 -560
rect 296671 -588 296719 -560
rect 296409 -622 296719 -588
rect 296409 -650 296457 -622
rect 296485 -650 296519 -622
rect 296547 -650 296581 -622
rect 296609 -650 296643 -622
rect 296671 -650 296719 -622
rect 296409 -684 296719 -650
rect 296409 -712 296457 -684
rect 296485 -712 296519 -684
rect 296547 -712 296581 -684
rect 296609 -712 296643 -684
rect 296671 -712 296719 -684
rect 296409 -746 296719 -712
rect 296409 -774 296457 -746
rect 296485 -774 296519 -746
rect 296547 -774 296581 -746
rect 296609 -774 296643 -746
rect 296671 -774 296719 -746
rect 296409 -822 296719 -774
rect 298680 -560 298990 4961
rect 298680 -588 298728 -560
rect 298756 -588 298790 -560
rect 298818 -588 298852 -560
rect 298880 -588 298914 -560
rect 298942 -588 298990 -560
rect 298680 -622 298990 -588
rect 298680 -650 298728 -622
rect 298756 -650 298790 -622
rect 298818 -650 298852 -622
rect 298880 -650 298914 -622
rect 298942 -650 298990 -622
rect 298680 -684 298990 -650
rect 298680 -712 298728 -684
rect 298756 -712 298790 -684
rect 298818 -712 298852 -684
rect 298880 -712 298914 -684
rect 298942 -712 298990 -684
rect 298680 -746 298990 -712
rect 298680 -774 298728 -746
rect 298756 -774 298790 -746
rect 298818 -774 298852 -746
rect 298880 -774 298914 -746
rect 298942 -774 298990 -746
rect 298680 -822 298990 -774
<< via4 >>
rect -910 299058 -882 299086
rect -848 299058 -820 299086
rect -786 299058 -758 299086
rect -724 299058 -696 299086
rect -910 298996 -882 299024
rect -848 298996 -820 299024
rect -786 298996 -758 299024
rect -724 298996 -696 299024
rect -910 298934 -882 298962
rect -848 298934 -820 298962
rect -786 298934 -758 298962
rect -724 298934 -696 298962
rect -910 298872 -882 298900
rect -848 298872 -820 298900
rect -786 298872 -758 298900
rect -724 298872 -696 298900
rect -910 293147 -882 293175
rect -848 293147 -820 293175
rect -786 293147 -758 293175
rect -724 293147 -696 293175
rect -910 293085 -882 293113
rect -848 293085 -820 293113
rect -786 293085 -758 293113
rect -724 293085 -696 293113
rect -910 293023 -882 293051
rect -848 293023 -820 293051
rect -786 293023 -758 293051
rect -724 293023 -696 293051
rect -910 292961 -882 292989
rect -848 292961 -820 292989
rect -786 292961 -758 292989
rect -724 292961 -696 292989
rect -910 284147 -882 284175
rect -848 284147 -820 284175
rect -786 284147 -758 284175
rect -724 284147 -696 284175
rect -910 284085 -882 284113
rect -848 284085 -820 284113
rect -786 284085 -758 284113
rect -724 284085 -696 284113
rect -910 284023 -882 284051
rect -848 284023 -820 284051
rect -786 284023 -758 284051
rect -724 284023 -696 284051
rect -910 283961 -882 283989
rect -848 283961 -820 283989
rect -786 283961 -758 283989
rect -724 283961 -696 283989
rect -910 275147 -882 275175
rect -848 275147 -820 275175
rect -786 275147 -758 275175
rect -724 275147 -696 275175
rect -910 275085 -882 275113
rect -848 275085 -820 275113
rect -786 275085 -758 275113
rect -724 275085 -696 275113
rect -910 275023 -882 275051
rect -848 275023 -820 275051
rect -786 275023 -758 275051
rect -724 275023 -696 275051
rect -910 274961 -882 274989
rect -848 274961 -820 274989
rect -786 274961 -758 274989
rect -724 274961 -696 274989
rect -910 266147 -882 266175
rect -848 266147 -820 266175
rect -786 266147 -758 266175
rect -724 266147 -696 266175
rect -910 266085 -882 266113
rect -848 266085 -820 266113
rect -786 266085 -758 266113
rect -724 266085 -696 266113
rect -910 266023 -882 266051
rect -848 266023 -820 266051
rect -786 266023 -758 266051
rect -724 266023 -696 266051
rect -910 265961 -882 265989
rect -848 265961 -820 265989
rect -786 265961 -758 265989
rect -724 265961 -696 265989
rect -910 257147 -882 257175
rect -848 257147 -820 257175
rect -786 257147 -758 257175
rect -724 257147 -696 257175
rect -910 257085 -882 257113
rect -848 257085 -820 257113
rect -786 257085 -758 257113
rect -724 257085 -696 257113
rect -910 257023 -882 257051
rect -848 257023 -820 257051
rect -786 257023 -758 257051
rect -724 257023 -696 257051
rect -910 256961 -882 256989
rect -848 256961 -820 256989
rect -786 256961 -758 256989
rect -724 256961 -696 256989
rect -910 248147 -882 248175
rect -848 248147 -820 248175
rect -786 248147 -758 248175
rect -724 248147 -696 248175
rect -910 248085 -882 248113
rect -848 248085 -820 248113
rect -786 248085 -758 248113
rect -724 248085 -696 248113
rect -910 248023 -882 248051
rect -848 248023 -820 248051
rect -786 248023 -758 248051
rect -724 248023 -696 248051
rect -910 247961 -882 247989
rect -848 247961 -820 247989
rect -786 247961 -758 247989
rect -724 247961 -696 247989
rect -910 239147 -882 239175
rect -848 239147 -820 239175
rect -786 239147 -758 239175
rect -724 239147 -696 239175
rect -910 239085 -882 239113
rect -848 239085 -820 239113
rect -786 239085 -758 239113
rect -724 239085 -696 239113
rect -910 239023 -882 239051
rect -848 239023 -820 239051
rect -786 239023 -758 239051
rect -724 239023 -696 239051
rect -910 238961 -882 238989
rect -848 238961 -820 238989
rect -786 238961 -758 238989
rect -724 238961 -696 238989
rect -910 230147 -882 230175
rect -848 230147 -820 230175
rect -786 230147 -758 230175
rect -724 230147 -696 230175
rect -910 230085 -882 230113
rect -848 230085 -820 230113
rect -786 230085 -758 230113
rect -724 230085 -696 230113
rect -910 230023 -882 230051
rect -848 230023 -820 230051
rect -786 230023 -758 230051
rect -724 230023 -696 230051
rect -910 229961 -882 229989
rect -848 229961 -820 229989
rect -786 229961 -758 229989
rect -724 229961 -696 229989
rect -910 221147 -882 221175
rect -848 221147 -820 221175
rect -786 221147 -758 221175
rect -724 221147 -696 221175
rect -910 221085 -882 221113
rect -848 221085 -820 221113
rect -786 221085 -758 221113
rect -724 221085 -696 221113
rect -910 221023 -882 221051
rect -848 221023 -820 221051
rect -786 221023 -758 221051
rect -724 221023 -696 221051
rect -910 220961 -882 220989
rect -848 220961 -820 220989
rect -786 220961 -758 220989
rect -724 220961 -696 220989
rect -910 212147 -882 212175
rect -848 212147 -820 212175
rect -786 212147 -758 212175
rect -724 212147 -696 212175
rect -910 212085 -882 212113
rect -848 212085 -820 212113
rect -786 212085 -758 212113
rect -724 212085 -696 212113
rect -910 212023 -882 212051
rect -848 212023 -820 212051
rect -786 212023 -758 212051
rect -724 212023 -696 212051
rect -910 211961 -882 211989
rect -848 211961 -820 211989
rect -786 211961 -758 211989
rect -724 211961 -696 211989
rect -910 203147 -882 203175
rect -848 203147 -820 203175
rect -786 203147 -758 203175
rect -724 203147 -696 203175
rect -910 203085 -882 203113
rect -848 203085 -820 203113
rect -786 203085 -758 203113
rect -724 203085 -696 203113
rect -910 203023 -882 203051
rect -848 203023 -820 203051
rect -786 203023 -758 203051
rect -724 203023 -696 203051
rect -910 202961 -882 202989
rect -848 202961 -820 202989
rect -786 202961 -758 202989
rect -724 202961 -696 202989
rect -910 194147 -882 194175
rect -848 194147 -820 194175
rect -786 194147 -758 194175
rect -724 194147 -696 194175
rect -910 194085 -882 194113
rect -848 194085 -820 194113
rect -786 194085 -758 194113
rect -724 194085 -696 194113
rect -910 194023 -882 194051
rect -848 194023 -820 194051
rect -786 194023 -758 194051
rect -724 194023 -696 194051
rect -910 193961 -882 193989
rect -848 193961 -820 193989
rect -786 193961 -758 193989
rect -724 193961 -696 193989
rect -910 185147 -882 185175
rect -848 185147 -820 185175
rect -786 185147 -758 185175
rect -724 185147 -696 185175
rect -910 185085 -882 185113
rect -848 185085 -820 185113
rect -786 185085 -758 185113
rect -724 185085 -696 185113
rect -910 185023 -882 185051
rect -848 185023 -820 185051
rect -786 185023 -758 185051
rect -724 185023 -696 185051
rect -910 184961 -882 184989
rect -848 184961 -820 184989
rect -786 184961 -758 184989
rect -724 184961 -696 184989
rect -910 176147 -882 176175
rect -848 176147 -820 176175
rect -786 176147 -758 176175
rect -724 176147 -696 176175
rect -910 176085 -882 176113
rect -848 176085 -820 176113
rect -786 176085 -758 176113
rect -724 176085 -696 176113
rect -910 176023 -882 176051
rect -848 176023 -820 176051
rect -786 176023 -758 176051
rect -724 176023 -696 176051
rect -910 175961 -882 175989
rect -848 175961 -820 175989
rect -786 175961 -758 175989
rect -724 175961 -696 175989
rect -910 167147 -882 167175
rect -848 167147 -820 167175
rect -786 167147 -758 167175
rect -724 167147 -696 167175
rect -910 167085 -882 167113
rect -848 167085 -820 167113
rect -786 167085 -758 167113
rect -724 167085 -696 167113
rect -910 167023 -882 167051
rect -848 167023 -820 167051
rect -786 167023 -758 167051
rect -724 167023 -696 167051
rect -910 166961 -882 166989
rect -848 166961 -820 166989
rect -786 166961 -758 166989
rect -724 166961 -696 166989
rect -910 158147 -882 158175
rect -848 158147 -820 158175
rect -786 158147 -758 158175
rect -724 158147 -696 158175
rect -910 158085 -882 158113
rect -848 158085 -820 158113
rect -786 158085 -758 158113
rect -724 158085 -696 158113
rect -910 158023 -882 158051
rect -848 158023 -820 158051
rect -786 158023 -758 158051
rect -724 158023 -696 158051
rect -910 157961 -882 157989
rect -848 157961 -820 157989
rect -786 157961 -758 157989
rect -724 157961 -696 157989
rect -910 149147 -882 149175
rect -848 149147 -820 149175
rect -786 149147 -758 149175
rect -724 149147 -696 149175
rect -910 149085 -882 149113
rect -848 149085 -820 149113
rect -786 149085 -758 149113
rect -724 149085 -696 149113
rect -910 149023 -882 149051
rect -848 149023 -820 149051
rect -786 149023 -758 149051
rect -724 149023 -696 149051
rect -910 148961 -882 148989
rect -848 148961 -820 148989
rect -786 148961 -758 148989
rect -724 148961 -696 148989
rect -910 140147 -882 140175
rect -848 140147 -820 140175
rect -786 140147 -758 140175
rect -724 140147 -696 140175
rect -910 140085 -882 140113
rect -848 140085 -820 140113
rect -786 140085 -758 140113
rect -724 140085 -696 140113
rect -910 140023 -882 140051
rect -848 140023 -820 140051
rect -786 140023 -758 140051
rect -724 140023 -696 140051
rect -910 139961 -882 139989
rect -848 139961 -820 139989
rect -786 139961 -758 139989
rect -724 139961 -696 139989
rect -910 131147 -882 131175
rect -848 131147 -820 131175
rect -786 131147 -758 131175
rect -724 131147 -696 131175
rect -910 131085 -882 131113
rect -848 131085 -820 131113
rect -786 131085 -758 131113
rect -724 131085 -696 131113
rect -910 131023 -882 131051
rect -848 131023 -820 131051
rect -786 131023 -758 131051
rect -724 131023 -696 131051
rect -910 130961 -882 130989
rect -848 130961 -820 130989
rect -786 130961 -758 130989
rect -724 130961 -696 130989
rect -910 122147 -882 122175
rect -848 122147 -820 122175
rect -786 122147 -758 122175
rect -724 122147 -696 122175
rect -910 122085 -882 122113
rect -848 122085 -820 122113
rect -786 122085 -758 122113
rect -724 122085 -696 122113
rect -910 122023 -882 122051
rect -848 122023 -820 122051
rect -786 122023 -758 122051
rect -724 122023 -696 122051
rect -910 121961 -882 121989
rect -848 121961 -820 121989
rect -786 121961 -758 121989
rect -724 121961 -696 121989
rect -910 113147 -882 113175
rect -848 113147 -820 113175
rect -786 113147 -758 113175
rect -724 113147 -696 113175
rect -910 113085 -882 113113
rect -848 113085 -820 113113
rect -786 113085 -758 113113
rect -724 113085 -696 113113
rect -910 113023 -882 113051
rect -848 113023 -820 113051
rect -786 113023 -758 113051
rect -724 113023 -696 113051
rect -910 112961 -882 112989
rect -848 112961 -820 112989
rect -786 112961 -758 112989
rect -724 112961 -696 112989
rect -910 104147 -882 104175
rect -848 104147 -820 104175
rect -786 104147 -758 104175
rect -724 104147 -696 104175
rect -910 104085 -882 104113
rect -848 104085 -820 104113
rect -786 104085 -758 104113
rect -724 104085 -696 104113
rect -910 104023 -882 104051
rect -848 104023 -820 104051
rect -786 104023 -758 104051
rect -724 104023 -696 104051
rect -910 103961 -882 103989
rect -848 103961 -820 103989
rect -786 103961 -758 103989
rect -724 103961 -696 103989
rect -910 95147 -882 95175
rect -848 95147 -820 95175
rect -786 95147 -758 95175
rect -724 95147 -696 95175
rect -910 95085 -882 95113
rect -848 95085 -820 95113
rect -786 95085 -758 95113
rect -724 95085 -696 95113
rect -910 95023 -882 95051
rect -848 95023 -820 95051
rect -786 95023 -758 95051
rect -724 95023 -696 95051
rect -910 94961 -882 94989
rect -848 94961 -820 94989
rect -786 94961 -758 94989
rect -724 94961 -696 94989
rect -910 86147 -882 86175
rect -848 86147 -820 86175
rect -786 86147 -758 86175
rect -724 86147 -696 86175
rect -910 86085 -882 86113
rect -848 86085 -820 86113
rect -786 86085 -758 86113
rect -724 86085 -696 86113
rect -910 86023 -882 86051
rect -848 86023 -820 86051
rect -786 86023 -758 86051
rect -724 86023 -696 86051
rect -910 85961 -882 85989
rect -848 85961 -820 85989
rect -786 85961 -758 85989
rect -724 85961 -696 85989
rect -910 77147 -882 77175
rect -848 77147 -820 77175
rect -786 77147 -758 77175
rect -724 77147 -696 77175
rect -910 77085 -882 77113
rect -848 77085 -820 77113
rect -786 77085 -758 77113
rect -724 77085 -696 77113
rect -910 77023 -882 77051
rect -848 77023 -820 77051
rect -786 77023 -758 77051
rect -724 77023 -696 77051
rect -910 76961 -882 76989
rect -848 76961 -820 76989
rect -786 76961 -758 76989
rect -724 76961 -696 76989
rect -910 68147 -882 68175
rect -848 68147 -820 68175
rect -786 68147 -758 68175
rect -724 68147 -696 68175
rect -910 68085 -882 68113
rect -848 68085 -820 68113
rect -786 68085 -758 68113
rect -724 68085 -696 68113
rect -910 68023 -882 68051
rect -848 68023 -820 68051
rect -786 68023 -758 68051
rect -724 68023 -696 68051
rect -910 67961 -882 67989
rect -848 67961 -820 67989
rect -786 67961 -758 67989
rect -724 67961 -696 67989
rect -910 59147 -882 59175
rect -848 59147 -820 59175
rect -786 59147 -758 59175
rect -724 59147 -696 59175
rect -910 59085 -882 59113
rect -848 59085 -820 59113
rect -786 59085 -758 59113
rect -724 59085 -696 59113
rect -910 59023 -882 59051
rect -848 59023 -820 59051
rect -786 59023 -758 59051
rect -724 59023 -696 59051
rect -910 58961 -882 58989
rect -848 58961 -820 58989
rect -786 58961 -758 58989
rect -724 58961 -696 58989
rect -910 50147 -882 50175
rect -848 50147 -820 50175
rect -786 50147 -758 50175
rect -724 50147 -696 50175
rect -910 50085 -882 50113
rect -848 50085 -820 50113
rect -786 50085 -758 50113
rect -724 50085 -696 50113
rect -910 50023 -882 50051
rect -848 50023 -820 50051
rect -786 50023 -758 50051
rect -724 50023 -696 50051
rect -910 49961 -882 49989
rect -848 49961 -820 49989
rect -786 49961 -758 49989
rect -724 49961 -696 49989
rect -910 41147 -882 41175
rect -848 41147 -820 41175
rect -786 41147 -758 41175
rect -724 41147 -696 41175
rect -910 41085 -882 41113
rect -848 41085 -820 41113
rect -786 41085 -758 41113
rect -724 41085 -696 41113
rect -910 41023 -882 41051
rect -848 41023 -820 41051
rect -786 41023 -758 41051
rect -724 41023 -696 41051
rect -910 40961 -882 40989
rect -848 40961 -820 40989
rect -786 40961 -758 40989
rect -724 40961 -696 40989
rect -910 32147 -882 32175
rect -848 32147 -820 32175
rect -786 32147 -758 32175
rect -724 32147 -696 32175
rect -910 32085 -882 32113
rect -848 32085 -820 32113
rect -786 32085 -758 32113
rect -724 32085 -696 32113
rect -910 32023 -882 32051
rect -848 32023 -820 32051
rect -786 32023 -758 32051
rect -724 32023 -696 32051
rect -910 31961 -882 31989
rect -848 31961 -820 31989
rect -786 31961 -758 31989
rect -724 31961 -696 31989
rect -910 23147 -882 23175
rect -848 23147 -820 23175
rect -786 23147 -758 23175
rect -724 23147 -696 23175
rect -910 23085 -882 23113
rect -848 23085 -820 23113
rect -786 23085 -758 23113
rect -724 23085 -696 23113
rect -910 23023 -882 23051
rect -848 23023 -820 23051
rect -786 23023 -758 23051
rect -724 23023 -696 23051
rect -910 22961 -882 22989
rect -848 22961 -820 22989
rect -786 22961 -758 22989
rect -724 22961 -696 22989
rect -910 14147 -882 14175
rect -848 14147 -820 14175
rect -786 14147 -758 14175
rect -724 14147 -696 14175
rect -910 14085 -882 14113
rect -848 14085 -820 14113
rect -786 14085 -758 14113
rect -724 14085 -696 14113
rect -910 14023 -882 14051
rect -848 14023 -820 14051
rect -786 14023 -758 14051
rect -724 14023 -696 14051
rect -910 13961 -882 13989
rect -848 13961 -820 13989
rect -786 13961 -758 13989
rect -724 13961 -696 13989
rect -910 5147 -882 5175
rect -848 5147 -820 5175
rect -786 5147 -758 5175
rect -724 5147 -696 5175
rect -910 5085 -882 5113
rect -848 5085 -820 5113
rect -786 5085 -758 5113
rect -724 5085 -696 5113
rect -910 5023 -882 5051
rect -848 5023 -820 5051
rect -786 5023 -758 5051
rect -724 5023 -696 5051
rect -910 4961 -882 4989
rect -848 4961 -820 4989
rect -786 4961 -758 4989
rect -724 4961 -696 4989
rect -430 298578 -402 298606
rect -368 298578 -340 298606
rect -306 298578 -278 298606
rect -244 298578 -216 298606
rect -430 298516 -402 298544
rect -368 298516 -340 298544
rect -306 298516 -278 298544
rect -244 298516 -216 298544
rect -430 298454 -402 298482
rect -368 298454 -340 298482
rect -306 298454 -278 298482
rect -244 298454 -216 298482
rect -430 298392 -402 298420
rect -368 298392 -340 298420
rect -306 298392 -278 298420
rect -244 298392 -216 298420
rect -430 290147 -402 290175
rect -368 290147 -340 290175
rect -306 290147 -278 290175
rect -244 290147 -216 290175
rect -430 290085 -402 290113
rect -368 290085 -340 290113
rect -306 290085 -278 290113
rect -244 290085 -216 290113
rect -430 290023 -402 290051
rect -368 290023 -340 290051
rect -306 290023 -278 290051
rect -244 290023 -216 290051
rect -430 289961 -402 289989
rect -368 289961 -340 289989
rect -306 289961 -278 289989
rect -244 289961 -216 289989
rect -430 281147 -402 281175
rect -368 281147 -340 281175
rect -306 281147 -278 281175
rect -244 281147 -216 281175
rect -430 281085 -402 281113
rect -368 281085 -340 281113
rect -306 281085 -278 281113
rect -244 281085 -216 281113
rect -430 281023 -402 281051
rect -368 281023 -340 281051
rect -306 281023 -278 281051
rect -244 281023 -216 281051
rect -430 280961 -402 280989
rect -368 280961 -340 280989
rect -306 280961 -278 280989
rect -244 280961 -216 280989
rect -430 272147 -402 272175
rect -368 272147 -340 272175
rect -306 272147 -278 272175
rect -244 272147 -216 272175
rect -430 272085 -402 272113
rect -368 272085 -340 272113
rect -306 272085 -278 272113
rect -244 272085 -216 272113
rect -430 272023 -402 272051
rect -368 272023 -340 272051
rect -306 272023 -278 272051
rect -244 272023 -216 272051
rect -430 271961 -402 271989
rect -368 271961 -340 271989
rect -306 271961 -278 271989
rect -244 271961 -216 271989
rect -430 263147 -402 263175
rect -368 263147 -340 263175
rect -306 263147 -278 263175
rect -244 263147 -216 263175
rect -430 263085 -402 263113
rect -368 263085 -340 263113
rect -306 263085 -278 263113
rect -244 263085 -216 263113
rect -430 263023 -402 263051
rect -368 263023 -340 263051
rect -306 263023 -278 263051
rect -244 263023 -216 263051
rect -430 262961 -402 262989
rect -368 262961 -340 262989
rect -306 262961 -278 262989
rect -244 262961 -216 262989
rect -430 254147 -402 254175
rect -368 254147 -340 254175
rect -306 254147 -278 254175
rect -244 254147 -216 254175
rect -430 254085 -402 254113
rect -368 254085 -340 254113
rect -306 254085 -278 254113
rect -244 254085 -216 254113
rect -430 254023 -402 254051
rect -368 254023 -340 254051
rect -306 254023 -278 254051
rect -244 254023 -216 254051
rect -430 253961 -402 253989
rect -368 253961 -340 253989
rect -306 253961 -278 253989
rect -244 253961 -216 253989
rect -430 245147 -402 245175
rect -368 245147 -340 245175
rect -306 245147 -278 245175
rect -244 245147 -216 245175
rect -430 245085 -402 245113
rect -368 245085 -340 245113
rect -306 245085 -278 245113
rect -244 245085 -216 245113
rect -430 245023 -402 245051
rect -368 245023 -340 245051
rect -306 245023 -278 245051
rect -244 245023 -216 245051
rect -430 244961 -402 244989
rect -368 244961 -340 244989
rect -306 244961 -278 244989
rect -244 244961 -216 244989
rect -430 236147 -402 236175
rect -368 236147 -340 236175
rect -306 236147 -278 236175
rect -244 236147 -216 236175
rect -430 236085 -402 236113
rect -368 236085 -340 236113
rect -306 236085 -278 236113
rect -244 236085 -216 236113
rect -430 236023 -402 236051
rect -368 236023 -340 236051
rect -306 236023 -278 236051
rect -244 236023 -216 236051
rect -430 235961 -402 235989
rect -368 235961 -340 235989
rect -306 235961 -278 235989
rect -244 235961 -216 235989
rect -430 227147 -402 227175
rect -368 227147 -340 227175
rect -306 227147 -278 227175
rect -244 227147 -216 227175
rect -430 227085 -402 227113
rect -368 227085 -340 227113
rect -306 227085 -278 227113
rect -244 227085 -216 227113
rect -430 227023 -402 227051
rect -368 227023 -340 227051
rect -306 227023 -278 227051
rect -244 227023 -216 227051
rect -430 226961 -402 226989
rect -368 226961 -340 226989
rect -306 226961 -278 226989
rect -244 226961 -216 226989
rect -430 218147 -402 218175
rect -368 218147 -340 218175
rect -306 218147 -278 218175
rect -244 218147 -216 218175
rect -430 218085 -402 218113
rect -368 218085 -340 218113
rect -306 218085 -278 218113
rect -244 218085 -216 218113
rect -430 218023 -402 218051
rect -368 218023 -340 218051
rect -306 218023 -278 218051
rect -244 218023 -216 218051
rect -430 217961 -402 217989
rect -368 217961 -340 217989
rect -306 217961 -278 217989
rect -244 217961 -216 217989
rect -430 209147 -402 209175
rect -368 209147 -340 209175
rect -306 209147 -278 209175
rect -244 209147 -216 209175
rect -430 209085 -402 209113
rect -368 209085 -340 209113
rect -306 209085 -278 209113
rect -244 209085 -216 209113
rect -430 209023 -402 209051
rect -368 209023 -340 209051
rect -306 209023 -278 209051
rect -244 209023 -216 209051
rect -430 208961 -402 208989
rect -368 208961 -340 208989
rect -306 208961 -278 208989
rect -244 208961 -216 208989
rect -430 200147 -402 200175
rect -368 200147 -340 200175
rect -306 200147 -278 200175
rect -244 200147 -216 200175
rect -430 200085 -402 200113
rect -368 200085 -340 200113
rect -306 200085 -278 200113
rect -244 200085 -216 200113
rect -430 200023 -402 200051
rect -368 200023 -340 200051
rect -306 200023 -278 200051
rect -244 200023 -216 200051
rect -430 199961 -402 199989
rect -368 199961 -340 199989
rect -306 199961 -278 199989
rect -244 199961 -216 199989
rect -430 191147 -402 191175
rect -368 191147 -340 191175
rect -306 191147 -278 191175
rect -244 191147 -216 191175
rect -430 191085 -402 191113
rect -368 191085 -340 191113
rect -306 191085 -278 191113
rect -244 191085 -216 191113
rect -430 191023 -402 191051
rect -368 191023 -340 191051
rect -306 191023 -278 191051
rect -244 191023 -216 191051
rect -430 190961 -402 190989
rect -368 190961 -340 190989
rect -306 190961 -278 190989
rect -244 190961 -216 190989
rect -430 182147 -402 182175
rect -368 182147 -340 182175
rect -306 182147 -278 182175
rect -244 182147 -216 182175
rect -430 182085 -402 182113
rect -368 182085 -340 182113
rect -306 182085 -278 182113
rect -244 182085 -216 182113
rect -430 182023 -402 182051
rect -368 182023 -340 182051
rect -306 182023 -278 182051
rect -244 182023 -216 182051
rect -430 181961 -402 181989
rect -368 181961 -340 181989
rect -306 181961 -278 181989
rect -244 181961 -216 181989
rect -430 173147 -402 173175
rect -368 173147 -340 173175
rect -306 173147 -278 173175
rect -244 173147 -216 173175
rect -430 173085 -402 173113
rect -368 173085 -340 173113
rect -306 173085 -278 173113
rect -244 173085 -216 173113
rect -430 173023 -402 173051
rect -368 173023 -340 173051
rect -306 173023 -278 173051
rect -244 173023 -216 173051
rect -430 172961 -402 172989
rect -368 172961 -340 172989
rect -306 172961 -278 172989
rect -244 172961 -216 172989
rect -430 164147 -402 164175
rect -368 164147 -340 164175
rect -306 164147 -278 164175
rect -244 164147 -216 164175
rect -430 164085 -402 164113
rect -368 164085 -340 164113
rect -306 164085 -278 164113
rect -244 164085 -216 164113
rect -430 164023 -402 164051
rect -368 164023 -340 164051
rect -306 164023 -278 164051
rect -244 164023 -216 164051
rect -430 163961 -402 163989
rect -368 163961 -340 163989
rect -306 163961 -278 163989
rect -244 163961 -216 163989
rect -430 155147 -402 155175
rect -368 155147 -340 155175
rect -306 155147 -278 155175
rect -244 155147 -216 155175
rect -430 155085 -402 155113
rect -368 155085 -340 155113
rect -306 155085 -278 155113
rect -244 155085 -216 155113
rect -430 155023 -402 155051
rect -368 155023 -340 155051
rect -306 155023 -278 155051
rect -244 155023 -216 155051
rect -430 154961 -402 154989
rect -368 154961 -340 154989
rect -306 154961 -278 154989
rect -244 154961 -216 154989
rect -430 146147 -402 146175
rect -368 146147 -340 146175
rect -306 146147 -278 146175
rect -244 146147 -216 146175
rect -430 146085 -402 146113
rect -368 146085 -340 146113
rect -306 146085 -278 146113
rect -244 146085 -216 146113
rect -430 146023 -402 146051
rect -368 146023 -340 146051
rect -306 146023 -278 146051
rect -244 146023 -216 146051
rect -430 145961 -402 145989
rect -368 145961 -340 145989
rect -306 145961 -278 145989
rect -244 145961 -216 145989
rect -430 137147 -402 137175
rect -368 137147 -340 137175
rect -306 137147 -278 137175
rect -244 137147 -216 137175
rect -430 137085 -402 137113
rect -368 137085 -340 137113
rect -306 137085 -278 137113
rect -244 137085 -216 137113
rect -430 137023 -402 137051
rect -368 137023 -340 137051
rect -306 137023 -278 137051
rect -244 137023 -216 137051
rect -430 136961 -402 136989
rect -368 136961 -340 136989
rect -306 136961 -278 136989
rect -244 136961 -216 136989
rect -430 128147 -402 128175
rect -368 128147 -340 128175
rect -306 128147 -278 128175
rect -244 128147 -216 128175
rect -430 128085 -402 128113
rect -368 128085 -340 128113
rect -306 128085 -278 128113
rect -244 128085 -216 128113
rect -430 128023 -402 128051
rect -368 128023 -340 128051
rect -306 128023 -278 128051
rect -244 128023 -216 128051
rect -430 127961 -402 127989
rect -368 127961 -340 127989
rect -306 127961 -278 127989
rect -244 127961 -216 127989
rect -430 119147 -402 119175
rect -368 119147 -340 119175
rect -306 119147 -278 119175
rect -244 119147 -216 119175
rect -430 119085 -402 119113
rect -368 119085 -340 119113
rect -306 119085 -278 119113
rect -244 119085 -216 119113
rect -430 119023 -402 119051
rect -368 119023 -340 119051
rect -306 119023 -278 119051
rect -244 119023 -216 119051
rect -430 118961 -402 118989
rect -368 118961 -340 118989
rect -306 118961 -278 118989
rect -244 118961 -216 118989
rect 2757 298578 2785 298606
rect 2819 298578 2847 298606
rect 2881 298578 2909 298606
rect 2943 298578 2971 298606
rect 2757 298516 2785 298544
rect 2819 298516 2847 298544
rect 2881 298516 2909 298544
rect 2943 298516 2971 298544
rect 2757 298454 2785 298482
rect 2819 298454 2847 298482
rect 2881 298454 2909 298482
rect 2943 298454 2971 298482
rect 2757 298392 2785 298420
rect 2819 298392 2847 298420
rect 2881 298392 2909 298420
rect 2943 298392 2971 298420
rect 2757 290147 2785 290175
rect 2819 290147 2847 290175
rect 2881 290147 2909 290175
rect 2943 290147 2971 290175
rect 2757 290085 2785 290113
rect 2819 290085 2847 290113
rect 2881 290085 2909 290113
rect 2943 290085 2971 290113
rect 2757 290023 2785 290051
rect 2819 290023 2847 290051
rect 2881 290023 2909 290051
rect 2943 290023 2971 290051
rect 2757 289961 2785 289989
rect 2819 289961 2847 289989
rect 2881 289961 2909 289989
rect 2943 289961 2971 289989
rect 2757 281147 2785 281175
rect 2819 281147 2847 281175
rect 2881 281147 2909 281175
rect 2943 281147 2971 281175
rect 2757 281085 2785 281113
rect 2819 281085 2847 281113
rect 2881 281085 2909 281113
rect 2943 281085 2971 281113
rect 2757 281023 2785 281051
rect 2819 281023 2847 281051
rect 2881 281023 2909 281051
rect 2943 281023 2971 281051
rect 2757 280961 2785 280989
rect 2819 280961 2847 280989
rect 2881 280961 2909 280989
rect 2943 280961 2971 280989
rect 2757 272147 2785 272175
rect 2819 272147 2847 272175
rect 2881 272147 2909 272175
rect 2943 272147 2971 272175
rect 2757 272085 2785 272113
rect 2819 272085 2847 272113
rect 2881 272085 2909 272113
rect 2943 272085 2971 272113
rect 2757 272023 2785 272051
rect 2819 272023 2847 272051
rect 2881 272023 2909 272051
rect 2943 272023 2971 272051
rect 2757 271961 2785 271989
rect 2819 271961 2847 271989
rect 2881 271961 2909 271989
rect 2943 271961 2971 271989
rect 2757 263147 2785 263175
rect 2819 263147 2847 263175
rect 2881 263147 2909 263175
rect 2943 263147 2971 263175
rect 2757 263085 2785 263113
rect 2819 263085 2847 263113
rect 2881 263085 2909 263113
rect 2943 263085 2971 263113
rect 2757 263023 2785 263051
rect 2819 263023 2847 263051
rect 2881 263023 2909 263051
rect 2943 263023 2971 263051
rect 2757 262961 2785 262989
rect 2819 262961 2847 262989
rect 2881 262961 2909 262989
rect 2943 262961 2971 262989
rect 2757 254147 2785 254175
rect 2819 254147 2847 254175
rect 2881 254147 2909 254175
rect 2943 254147 2971 254175
rect 2757 254085 2785 254113
rect 2819 254085 2847 254113
rect 2881 254085 2909 254113
rect 2943 254085 2971 254113
rect 2757 254023 2785 254051
rect 2819 254023 2847 254051
rect 2881 254023 2909 254051
rect 2943 254023 2971 254051
rect 2757 253961 2785 253989
rect 2819 253961 2847 253989
rect 2881 253961 2909 253989
rect 2943 253961 2971 253989
rect 2757 245147 2785 245175
rect 2819 245147 2847 245175
rect 2881 245147 2909 245175
rect 2943 245147 2971 245175
rect 2757 245085 2785 245113
rect 2819 245085 2847 245113
rect 2881 245085 2909 245113
rect 2943 245085 2971 245113
rect 2757 245023 2785 245051
rect 2819 245023 2847 245051
rect 2881 245023 2909 245051
rect 2943 245023 2971 245051
rect 2757 244961 2785 244989
rect 2819 244961 2847 244989
rect 2881 244961 2909 244989
rect 2943 244961 2971 244989
rect 2757 236147 2785 236175
rect 2819 236147 2847 236175
rect 2881 236147 2909 236175
rect 2943 236147 2971 236175
rect 2757 236085 2785 236113
rect 2819 236085 2847 236113
rect 2881 236085 2909 236113
rect 2943 236085 2971 236113
rect 2757 236023 2785 236051
rect 2819 236023 2847 236051
rect 2881 236023 2909 236051
rect 2943 236023 2971 236051
rect 2757 235961 2785 235989
rect 2819 235961 2847 235989
rect 2881 235961 2909 235989
rect 2943 235961 2971 235989
rect 2757 227147 2785 227175
rect 2819 227147 2847 227175
rect 2881 227147 2909 227175
rect 2943 227147 2971 227175
rect 2757 227085 2785 227113
rect 2819 227085 2847 227113
rect 2881 227085 2909 227113
rect 2943 227085 2971 227113
rect 2757 227023 2785 227051
rect 2819 227023 2847 227051
rect 2881 227023 2909 227051
rect 2943 227023 2971 227051
rect 2757 226961 2785 226989
rect 2819 226961 2847 226989
rect 2881 226961 2909 226989
rect 2943 226961 2971 226989
rect 2757 218147 2785 218175
rect 2819 218147 2847 218175
rect 2881 218147 2909 218175
rect 2943 218147 2971 218175
rect 2757 218085 2785 218113
rect 2819 218085 2847 218113
rect 2881 218085 2909 218113
rect 2943 218085 2971 218113
rect 2757 218023 2785 218051
rect 2819 218023 2847 218051
rect 2881 218023 2909 218051
rect 2943 218023 2971 218051
rect 2757 217961 2785 217989
rect 2819 217961 2847 217989
rect 2881 217961 2909 217989
rect 2943 217961 2971 217989
rect 2757 209147 2785 209175
rect 2819 209147 2847 209175
rect 2881 209147 2909 209175
rect 2943 209147 2971 209175
rect 2757 209085 2785 209113
rect 2819 209085 2847 209113
rect 2881 209085 2909 209113
rect 2943 209085 2971 209113
rect 2757 209023 2785 209051
rect 2819 209023 2847 209051
rect 2881 209023 2909 209051
rect 2943 209023 2971 209051
rect 2757 208961 2785 208989
rect 2819 208961 2847 208989
rect 2881 208961 2909 208989
rect 2943 208961 2971 208989
rect 2757 200147 2785 200175
rect 2819 200147 2847 200175
rect 2881 200147 2909 200175
rect 2943 200147 2971 200175
rect 2757 200085 2785 200113
rect 2819 200085 2847 200113
rect 2881 200085 2909 200113
rect 2943 200085 2971 200113
rect 2757 200023 2785 200051
rect 2819 200023 2847 200051
rect 2881 200023 2909 200051
rect 2943 200023 2971 200051
rect 2757 199961 2785 199989
rect 2819 199961 2847 199989
rect 2881 199961 2909 199989
rect 2943 199961 2971 199989
rect 2757 191147 2785 191175
rect 2819 191147 2847 191175
rect 2881 191147 2909 191175
rect 2943 191147 2971 191175
rect 2757 191085 2785 191113
rect 2819 191085 2847 191113
rect 2881 191085 2909 191113
rect 2943 191085 2971 191113
rect 2757 191023 2785 191051
rect 2819 191023 2847 191051
rect 2881 191023 2909 191051
rect 2943 191023 2971 191051
rect 2757 190961 2785 190989
rect 2819 190961 2847 190989
rect 2881 190961 2909 190989
rect 2943 190961 2971 190989
rect 2757 182147 2785 182175
rect 2819 182147 2847 182175
rect 2881 182147 2909 182175
rect 2943 182147 2971 182175
rect 2757 182085 2785 182113
rect 2819 182085 2847 182113
rect 2881 182085 2909 182113
rect 2943 182085 2971 182113
rect 2757 182023 2785 182051
rect 2819 182023 2847 182051
rect 2881 182023 2909 182051
rect 2943 182023 2971 182051
rect 2757 181961 2785 181989
rect 2819 181961 2847 181989
rect 2881 181961 2909 181989
rect 2943 181961 2971 181989
rect 4617 299058 4645 299086
rect 4679 299058 4707 299086
rect 4741 299058 4769 299086
rect 4803 299058 4831 299086
rect 4617 298996 4645 299024
rect 4679 298996 4707 299024
rect 4741 298996 4769 299024
rect 4803 298996 4831 299024
rect 4617 298934 4645 298962
rect 4679 298934 4707 298962
rect 4741 298934 4769 298962
rect 4803 298934 4831 298962
rect 4617 298872 4645 298900
rect 4679 298872 4707 298900
rect 4741 298872 4769 298900
rect 4803 298872 4831 298900
rect 4617 293147 4645 293175
rect 4679 293147 4707 293175
rect 4741 293147 4769 293175
rect 4803 293147 4831 293175
rect 4617 293085 4645 293113
rect 4679 293085 4707 293113
rect 4741 293085 4769 293113
rect 4803 293085 4831 293113
rect 4617 293023 4645 293051
rect 4679 293023 4707 293051
rect 4741 293023 4769 293051
rect 4803 293023 4831 293051
rect 4617 292961 4645 292989
rect 4679 292961 4707 292989
rect 4741 292961 4769 292989
rect 4803 292961 4831 292989
rect 4617 284147 4645 284175
rect 4679 284147 4707 284175
rect 4741 284147 4769 284175
rect 4803 284147 4831 284175
rect 4617 284085 4645 284113
rect 4679 284085 4707 284113
rect 4741 284085 4769 284113
rect 4803 284085 4831 284113
rect 4617 284023 4645 284051
rect 4679 284023 4707 284051
rect 4741 284023 4769 284051
rect 4803 284023 4831 284051
rect 4617 283961 4645 283989
rect 4679 283961 4707 283989
rect 4741 283961 4769 283989
rect 4803 283961 4831 283989
rect 4617 275147 4645 275175
rect 4679 275147 4707 275175
rect 4741 275147 4769 275175
rect 4803 275147 4831 275175
rect 4617 275085 4645 275113
rect 4679 275085 4707 275113
rect 4741 275085 4769 275113
rect 4803 275085 4831 275113
rect 4617 275023 4645 275051
rect 4679 275023 4707 275051
rect 4741 275023 4769 275051
rect 4803 275023 4831 275051
rect 4617 274961 4645 274989
rect 4679 274961 4707 274989
rect 4741 274961 4769 274989
rect 4803 274961 4831 274989
rect 4617 266147 4645 266175
rect 4679 266147 4707 266175
rect 4741 266147 4769 266175
rect 4803 266147 4831 266175
rect 4617 266085 4645 266113
rect 4679 266085 4707 266113
rect 4741 266085 4769 266113
rect 4803 266085 4831 266113
rect 4617 266023 4645 266051
rect 4679 266023 4707 266051
rect 4741 266023 4769 266051
rect 4803 266023 4831 266051
rect 4617 265961 4645 265989
rect 4679 265961 4707 265989
rect 4741 265961 4769 265989
rect 4803 265961 4831 265989
rect 4617 257147 4645 257175
rect 4679 257147 4707 257175
rect 4741 257147 4769 257175
rect 4803 257147 4831 257175
rect 4617 257085 4645 257113
rect 4679 257085 4707 257113
rect 4741 257085 4769 257113
rect 4803 257085 4831 257113
rect 4617 257023 4645 257051
rect 4679 257023 4707 257051
rect 4741 257023 4769 257051
rect 4803 257023 4831 257051
rect 4617 256961 4645 256989
rect 4679 256961 4707 256989
rect 4741 256961 4769 256989
rect 4803 256961 4831 256989
rect 4617 248147 4645 248175
rect 4679 248147 4707 248175
rect 4741 248147 4769 248175
rect 4803 248147 4831 248175
rect 4617 248085 4645 248113
rect 4679 248085 4707 248113
rect 4741 248085 4769 248113
rect 4803 248085 4831 248113
rect 4617 248023 4645 248051
rect 4679 248023 4707 248051
rect 4741 248023 4769 248051
rect 4803 248023 4831 248051
rect 4617 247961 4645 247989
rect 4679 247961 4707 247989
rect 4741 247961 4769 247989
rect 4803 247961 4831 247989
rect 4617 239147 4645 239175
rect 4679 239147 4707 239175
rect 4741 239147 4769 239175
rect 4803 239147 4831 239175
rect 4617 239085 4645 239113
rect 4679 239085 4707 239113
rect 4741 239085 4769 239113
rect 4803 239085 4831 239113
rect 4617 239023 4645 239051
rect 4679 239023 4707 239051
rect 4741 239023 4769 239051
rect 4803 239023 4831 239051
rect 4617 238961 4645 238989
rect 4679 238961 4707 238989
rect 4741 238961 4769 238989
rect 4803 238961 4831 238989
rect 4617 230147 4645 230175
rect 4679 230147 4707 230175
rect 4741 230147 4769 230175
rect 4803 230147 4831 230175
rect 4617 230085 4645 230113
rect 4679 230085 4707 230113
rect 4741 230085 4769 230113
rect 4803 230085 4831 230113
rect 4617 230023 4645 230051
rect 4679 230023 4707 230051
rect 4741 230023 4769 230051
rect 4803 230023 4831 230051
rect 4617 229961 4645 229989
rect 4679 229961 4707 229989
rect 4741 229961 4769 229989
rect 4803 229961 4831 229989
rect 4617 221147 4645 221175
rect 4679 221147 4707 221175
rect 4741 221147 4769 221175
rect 4803 221147 4831 221175
rect 4617 221085 4645 221113
rect 4679 221085 4707 221113
rect 4741 221085 4769 221113
rect 4803 221085 4831 221113
rect 4617 221023 4645 221051
rect 4679 221023 4707 221051
rect 4741 221023 4769 221051
rect 4803 221023 4831 221051
rect 4617 220961 4645 220989
rect 4679 220961 4707 220989
rect 4741 220961 4769 220989
rect 4803 220961 4831 220989
rect 4617 212147 4645 212175
rect 4679 212147 4707 212175
rect 4741 212147 4769 212175
rect 4803 212147 4831 212175
rect 4617 212085 4645 212113
rect 4679 212085 4707 212113
rect 4741 212085 4769 212113
rect 4803 212085 4831 212113
rect 4617 212023 4645 212051
rect 4679 212023 4707 212051
rect 4741 212023 4769 212051
rect 4803 212023 4831 212051
rect 4617 211961 4645 211989
rect 4679 211961 4707 211989
rect 4741 211961 4769 211989
rect 4803 211961 4831 211989
rect 4617 203147 4645 203175
rect 4679 203147 4707 203175
rect 4741 203147 4769 203175
rect 4803 203147 4831 203175
rect 4617 203085 4645 203113
rect 4679 203085 4707 203113
rect 4741 203085 4769 203113
rect 4803 203085 4831 203113
rect 4617 203023 4645 203051
rect 4679 203023 4707 203051
rect 4741 203023 4769 203051
rect 4803 203023 4831 203051
rect 4617 202961 4645 202989
rect 4679 202961 4707 202989
rect 4741 202961 4769 202989
rect 4803 202961 4831 202989
rect 4617 194147 4645 194175
rect 4679 194147 4707 194175
rect 4741 194147 4769 194175
rect 4803 194147 4831 194175
rect 4617 194085 4645 194113
rect 4679 194085 4707 194113
rect 4741 194085 4769 194113
rect 4803 194085 4831 194113
rect 4617 194023 4645 194051
rect 4679 194023 4707 194051
rect 4741 194023 4769 194051
rect 4803 194023 4831 194051
rect 4617 193961 4645 193989
rect 4679 193961 4707 193989
rect 4741 193961 4769 193989
rect 4803 193961 4831 193989
rect 4617 185147 4645 185175
rect 4679 185147 4707 185175
rect 4741 185147 4769 185175
rect 4803 185147 4831 185175
rect 4617 185085 4645 185113
rect 4679 185085 4707 185113
rect 4741 185085 4769 185113
rect 4803 185085 4831 185113
rect 4617 185023 4645 185051
rect 4679 185023 4707 185051
rect 4741 185023 4769 185051
rect 4803 185023 4831 185051
rect 4617 184961 4645 184989
rect 4679 184961 4707 184989
rect 4741 184961 4769 184989
rect 4803 184961 4831 184989
rect 4617 176147 4645 176175
rect 4679 176147 4707 176175
rect 4741 176147 4769 176175
rect 4803 176147 4831 176175
rect 4617 176085 4645 176113
rect 4679 176085 4707 176113
rect 4741 176085 4769 176113
rect 4803 176085 4831 176113
rect 4617 176023 4645 176051
rect 4679 176023 4707 176051
rect 4741 176023 4769 176051
rect 4803 176023 4831 176051
rect 4617 175961 4645 175989
rect 4679 175961 4707 175989
rect 4741 175961 4769 175989
rect 4803 175961 4831 175989
rect 2757 173147 2785 173175
rect 2819 173147 2847 173175
rect 2881 173147 2909 173175
rect 2943 173147 2971 173175
rect 2757 173085 2785 173113
rect 2819 173085 2847 173113
rect 2881 173085 2909 173113
rect 2943 173085 2971 173113
rect 2757 173023 2785 173051
rect 2819 173023 2847 173051
rect 2881 173023 2909 173051
rect 2943 173023 2971 173051
rect 2757 172961 2785 172989
rect 2819 172961 2847 172989
rect 2881 172961 2909 172989
rect 2943 172961 2971 172989
rect 18117 298578 18145 298606
rect 18179 298578 18207 298606
rect 18241 298578 18269 298606
rect 18303 298578 18331 298606
rect 18117 298516 18145 298544
rect 18179 298516 18207 298544
rect 18241 298516 18269 298544
rect 18303 298516 18331 298544
rect 18117 298454 18145 298482
rect 18179 298454 18207 298482
rect 18241 298454 18269 298482
rect 18303 298454 18331 298482
rect 18117 298392 18145 298420
rect 18179 298392 18207 298420
rect 18241 298392 18269 298420
rect 18303 298392 18331 298420
rect 18117 290147 18145 290175
rect 18179 290147 18207 290175
rect 18241 290147 18269 290175
rect 18303 290147 18331 290175
rect 18117 290085 18145 290113
rect 18179 290085 18207 290113
rect 18241 290085 18269 290113
rect 18303 290085 18331 290113
rect 18117 290023 18145 290051
rect 18179 290023 18207 290051
rect 18241 290023 18269 290051
rect 18303 290023 18331 290051
rect 18117 289961 18145 289989
rect 18179 289961 18207 289989
rect 18241 289961 18269 289989
rect 18303 289961 18331 289989
rect 18117 281147 18145 281175
rect 18179 281147 18207 281175
rect 18241 281147 18269 281175
rect 18303 281147 18331 281175
rect 18117 281085 18145 281113
rect 18179 281085 18207 281113
rect 18241 281085 18269 281113
rect 18303 281085 18331 281113
rect 18117 281023 18145 281051
rect 18179 281023 18207 281051
rect 18241 281023 18269 281051
rect 18303 281023 18331 281051
rect 18117 280961 18145 280989
rect 18179 280961 18207 280989
rect 18241 280961 18269 280989
rect 18303 280961 18331 280989
rect 18117 272147 18145 272175
rect 18179 272147 18207 272175
rect 18241 272147 18269 272175
rect 18303 272147 18331 272175
rect 18117 272085 18145 272113
rect 18179 272085 18207 272113
rect 18241 272085 18269 272113
rect 18303 272085 18331 272113
rect 18117 272023 18145 272051
rect 18179 272023 18207 272051
rect 18241 272023 18269 272051
rect 18303 272023 18331 272051
rect 18117 271961 18145 271989
rect 18179 271961 18207 271989
rect 18241 271961 18269 271989
rect 18303 271961 18331 271989
rect 18117 263147 18145 263175
rect 18179 263147 18207 263175
rect 18241 263147 18269 263175
rect 18303 263147 18331 263175
rect 18117 263085 18145 263113
rect 18179 263085 18207 263113
rect 18241 263085 18269 263113
rect 18303 263085 18331 263113
rect 18117 263023 18145 263051
rect 18179 263023 18207 263051
rect 18241 263023 18269 263051
rect 18303 263023 18331 263051
rect 18117 262961 18145 262989
rect 18179 262961 18207 262989
rect 18241 262961 18269 262989
rect 18303 262961 18331 262989
rect 18117 254147 18145 254175
rect 18179 254147 18207 254175
rect 18241 254147 18269 254175
rect 18303 254147 18331 254175
rect 18117 254085 18145 254113
rect 18179 254085 18207 254113
rect 18241 254085 18269 254113
rect 18303 254085 18331 254113
rect 18117 254023 18145 254051
rect 18179 254023 18207 254051
rect 18241 254023 18269 254051
rect 18303 254023 18331 254051
rect 18117 253961 18145 253989
rect 18179 253961 18207 253989
rect 18241 253961 18269 253989
rect 18303 253961 18331 253989
rect 18117 245147 18145 245175
rect 18179 245147 18207 245175
rect 18241 245147 18269 245175
rect 18303 245147 18331 245175
rect 18117 245085 18145 245113
rect 18179 245085 18207 245113
rect 18241 245085 18269 245113
rect 18303 245085 18331 245113
rect 18117 245023 18145 245051
rect 18179 245023 18207 245051
rect 18241 245023 18269 245051
rect 18303 245023 18331 245051
rect 18117 244961 18145 244989
rect 18179 244961 18207 244989
rect 18241 244961 18269 244989
rect 18303 244961 18331 244989
rect 18117 236147 18145 236175
rect 18179 236147 18207 236175
rect 18241 236147 18269 236175
rect 18303 236147 18331 236175
rect 18117 236085 18145 236113
rect 18179 236085 18207 236113
rect 18241 236085 18269 236113
rect 18303 236085 18331 236113
rect 18117 236023 18145 236051
rect 18179 236023 18207 236051
rect 18241 236023 18269 236051
rect 18303 236023 18331 236051
rect 18117 235961 18145 235989
rect 18179 235961 18207 235989
rect 18241 235961 18269 235989
rect 18303 235961 18331 235989
rect 18117 227147 18145 227175
rect 18179 227147 18207 227175
rect 18241 227147 18269 227175
rect 18303 227147 18331 227175
rect 18117 227085 18145 227113
rect 18179 227085 18207 227113
rect 18241 227085 18269 227113
rect 18303 227085 18331 227113
rect 18117 227023 18145 227051
rect 18179 227023 18207 227051
rect 18241 227023 18269 227051
rect 18303 227023 18331 227051
rect 18117 226961 18145 226989
rect 18179 226961 18207 226989
rect 18241 226961 18269 226989
rect 18303 226961 18331 226989
rect 18117 218147 18145 218175
rect 18179 218147 18207 218175
rect 18241 218147 18269 218175
rect 18303 218147 18331 218175
rect 18117 218085 18145 218113
rect 18179 218085 18207 218113
rect 18241 218085 18269 218113
rect 18303 218085 18331 218113
rect 18117 218023 18145 218051
rect 18179 218023 18207 218051
rect 18241 218023 18269 218051
rect 18303 218023 18331 218051
rect 18117 217961 18145 217989
rect 18179 217961 18207 217989
rect 18241 217961 18269 217989
rect 18303 217961 18331 217989
rect 18117 209147 18145 209175
rect 18179 209147 18207 209175
rect 18241 209147 18269 209175
rect 18303 209147 18331 209175
rect 18117 209085 18145 209113
rect 18179 209085 18207 209113
rect 18241 209085 18269 209113
rect 18303 209085 18331 209113
rect 18117 209023 18145 209051
rect 18179 209023 18207 209051
rect 18241 209023 18269 209051
rect 18303 209023 18331 209051
rect 18117 208961 18145 208989
rect 18179 208961 18207 208989
rect 18241 208961 18269 208989
rect 18303 208961 18331 208989
rect 18117 200147 18145 200175
rect 18179 200147 18207 200175
rect 18241 200147 18269 200175
rect 18303 200147 18331 200175
rect 18117 200085 18145 200113
rect 18179 200085 18207 200113
rect 18241 200085 18269 200113
rect 18303 200085 18331 200113
rect 18117 200023 18145 200051
rect 18179 200023 18207 200051
rect 18241 200023 18269 200051
rect 18303 200023 18331 200051
rect 18117 199961 18145 199989
rect 18179 199961 18207 199989
rect 18241 199961 18269 199989
rect 18303 199961 18331 199989
rect 18117 191147 18145 191175
rect 18179 191147 18207 191175
rect 18241 191147 18269 191175
rect 18303 191147 18331 191175
rect 18117 191085 18145 191113
rect 18179 191085 18207 191113
rect 18241 191085 18269 191113
rect 18303 191085 18331 191113
rect 18117 191023 18145 191051
rect 18179 191023 18207 191051
rect 18241 191023 18269 191051
rect 18303 191023 18331 191051
rect 18117 190961 18145 190989
rect 18179 190961 18207 190989
rect 18241 190961 18269 190989
rect 18303 190961 18331 190989
rect 18117 182147 18145 182175
rect 18179 182147 18207 182175
rect 18241 182147 18269 182175
rect 18303 182147 18331 182175
rect 18117 182085 18145 182113
rect 18179 182085 18207 182113
rect 18241 182085 18269 182113
rect 18303 182085 18331 182113
rect 18117 182023 18145 182051
rect 18179 182023 18207 182051
rect 18241 182023 18269 182051
rect 18303 182023 18331 182051
rect 18117 181961 18145 181989
rect 18179 181961 18207 181989
rect 18241 181961 18269 181989
rect 18303 181961 18331 181989
rect 8259 173147 8287 173175
rect 8321 173147 8349 173175
rect 8259 173085 8287 173113
rect 8321 173085 8349 173113
rect 8259 173023 8287 173051
rect 8321 173023 8349 173051
rect 8259 172961 8287 172989
rect 8321 172961 8349 172989
rect 18117 173147 18145 173175
rect 18179 173147 18207 173175
rect 18241 173147 18269 173175
rect 18303 173147 18331 173175
rect 18117 173085 18145 173113
rect 18179 173085 18207 173113
rect 18241 173085 18269 173113
rect 18303 173085 18331 173113
rect 18117 173023 18145 173051
rect 18179 173023 18207 173051
rect 18241 173023 18269 173051
rect 18303 173023 18331 173051
rect 18117 172961 18145 172989
rect 18179 172961 18207 172989
rect 18241 172961 18269 172989
rect 18303 172961 18331 172989
rect 4617 167147 4645 167175
rect 4679 167147 4707 167175
rect 4741 167147 4769 167175
rect 4803 167147 4831 167175
rect 4617 167085 4645 167113
rect 4679 167085 4707 167113
rect 4741 167085 4769 167113
rect 4803 167085 4831 167113
rect 4617 167023 4645 167051
rect 4679 167023 4707 167051
rect 4741 167023 4769 167051
rect 4803 167023 4831 167051
rect 4617 166961 4645 166989
rect 4679 166961 4707 166989
rect 4741 166961 4769 166989
rect 4803 166961 4831 166989
rect 2757 164147 2785 164175
rect 2819 164147 2847 164175
rect 2881 164147 2909 164175
rect 2943 164147 2971 164175
rect 2757 164085 2785 164113
rect 2819 164085 2847 164113
rect 2881 164085 2909 164113
rect 2943 164085 2971 164113
rect 2757 164023 2785 164051
rect 2819 164023 2847 164051
rect 2881 164023 2909 164051
rect 2943 164023 2971 164051
rect 2757 163961 2785 163989
rect 2819 163961 2847 163989
rect 2881 163961 2909 163989
rect 2943 163961 2971 163989
rect 2757 155147 2785 155175
rect 2819 155147 2847 155175
rect 2881 155147 2909 155175
rect 2943 155147 2971 155175
rect 2757 155085 2785 155113
rect 2819 155085 2847 155113
rect 2881 155085 2909 155113
rect 2943 155085 2971 155113
rect 2757 155023 2785 155051
rect 2819 155023 2847 155051
rect 2881 155023 2909 155051
rect 2943 155023 2971 155051
rect 2757 154961 2785 154989
rect 2819 154961 2847 154989
rect 2881 154961 2909 154989
rect 2943 154961 2971 154989
rect 15939 167147 15967 167175
rect 16001 167147 16029 167175
rect 15939 167085 15967 167113
rect 16001 167085 16029 167113
rect 15939 167023 15967 167051
rect 16001 167023 16029 167051
rect 15939 166961 15967 166989
rect 16001 166961 16029 166989
rect 8259 164147 8287 164175
rect 8321 164147 8349 164175
rect 8259 164085 8287 164113
rect 8321 164085 8349 164113
rect 8259 164023 8287 164051
rect 8321 164023 8349 164051
rect 8259 163961 8287 163989
rect 8321 163961 8349 163989
rect 18117 164147 18145 164175
rect 18179 164147 18207 164175
rect 18241 164147 18269 164175
rect 18303 164147 18331 164175
rect 18117 164085 18145 164113
rect 18179 164085 18207 164113
rect 18241 164085 18269 164113
rect 18303 164085 18331 164113
rect 18117 164023 18145 164051
rect 18179 164023 18207 164051
rect 18241 164023 18269 164051
rect 18303 164023 18331 164051
rect 18117 163961 18145 163989
rect 18179 163961 18207 163989
rect 18241 163961 18269 163989
rect 18303 163961 18331 163989
rect 4617 158147 4645 158175
rect 4679 158147 4707 158175
rect 4741 158147 4769 158175
rect 4803 158147 4831 158175
rect 4617 158085 4645 158113
rect 4679 158085 4707 158113
rect 4741 158085 4769 158113
rect 4803 158085 4831 158113
rect 4617 158023 4645 158051
rect 4679 158023 4707 158051
rect 4741 158023 4769 158051
rect 4803 158023 4831 158051
rect 4617 157961 4645 157989
rect 4679 157961 4707 157989
rect 4741 157961 4769 157989
rect 4803 157961 4831 157989
rect 2757 146147 2785 146175
rect 2819 146147 2847 146175
rect 2881 146147 2909 146175
rect 2943 146147 2971 146175
rect 2757 146085 2785 146113
rect 2819 146085 2847 146113
rect 2881 146085 2909 146113
rect 2943 146085 2971 146113
rect 2757 146023 2785 146051
rect 2819 146023 2847 146051
rect 2881 146023 2909 146051
rect 2943 146023 2971 146051
rect 2757 145961 2785 145989
rect 2819 145961 2847 145989
rect 2881 145961 2909 145989
rect 2943 145961 2971 145989
rect 15939 158147 15967 158175
rect 16001 158147 16029 158175
rect 15939 158085 15967 158113
rect 16001 158085 16029 158113
rect 15939 158023 15967 158051
rect 16001 158023 16029 158051
rect 15939 157961 15967 157989
rect 16001 157961 16029 157989
rect 8259 155147 8287 155175
rect 8321 155147 8349 155175
rect 8259 155085 8287 155113
rect 8321 155085 8349 155113
rect 8259 155023 8287 155051
rect 8321 155023 8349 155051
rect 8259 154961 8287 154989
rect 8321 154961 8349 154989
rect 18117 155147 18145 155175
rect 18179 155147 18207 155175
rect 18241 155147 18269 155175
rect 18303 155147 18331 155175
rect 18117 155085 18145 155113
rect 18179 155085 18207 155113
rect 18241 155085 18269 155113
rect 18303 155085 18331 155113
rect 18117 155023 18145 155051
rect 18179 155023 18207 155051
rect 18241 155023 18269 155051
rect 18303 155023 18331 155051
rect 18117 154961 18145 154989
rect 18179 154961 18207 154989
rect 18241 154961 18269 154989
rect 18303 154961 18331 154989
rect 4617 149147 4645 149175
rect 4679 149147 4707 149175
rect 4741 149147 4769 149175
rect 4803 149147 4831 149175
rect 4617 149085 4645 149113
rect 4679 149085 4707 149113
rect 4741 149085 4769 149113
rect 4803 149085 4831 149113
rect 4617 149023 4645 149051
rect 4679 149023 4707 149051
rect 4741 149023 4769 149051
rect 4803 149023 4831 149051
rect 4617 148961 4645 148989
rect 4679 148961 4707 148989
rect 4741 148961 4769 148989
rect 4803 148961 4831 148989
rect 15939 149147 15967 149175
rect 16001 149147 16029 149175
rect 15939 149085 15967 149113
rect 16001 149085 16029 149113
rect 15939 149023 15967 149051
rect 16001 149023 16029 149051
rect 15939 148961 15967 148989
rect 16001 148961 16029 148989
rect 8259 146147 8287 146175
rect 8321 146147 8349 146175
rect 8259 146085 8287 146113
rect 8321 146085 8349 146113
rect 8259 146023 8287 146051
rect 8321 146023 8349 146051
rect 8259 145961 8287 145989
rect 8321 145961 8349 145989
rect 18117 146147 18145 146175
rect 18179 146147 18207 146175
rect 18241 146147 18269 146175
rect 18303 146147 18331 146175
rect 18117 146085 18145 146113
rect 18179 146085 18207 146113
rect 18241 146085 18269 146113
rect 18303 146085 18331 146113
rect 18117 146023 18145 146051
rect 18179 146023 18207 146051
rect 18241 146023 18269 146051
rect 18303 146023 18331 146051
rect 18117 145961 18145 145989
rect 18179 145961 18207 145989
rect 18241 145961 18269 145989
rect 18303 145961 18331 145989
rect 4617 140147 4645 140175
rect 4679 140147 4707 140175
rect 4741 140147 4769 140175
rect 4803 140147 4831 140175
rect 4617 140085 4645 140113
rect 4679 140085 4707 140113
rect 4741 140085 4769 140113
rect 4803 140085 4831 140113
rect 4617 140023 4645 140051
rect 4679 140023 4707 140051
rect 4741 140023 4769 140051
rect 4803 140023 4831 140051
rect 4617 139961 4645 139989
rect 4679 139961 4707 139989
rect 4741 139961 4769 139989
rect 4803 139961 4831 139989
rect 2757 137147 2785 137175
rect 2819 137147 2847 137175
rect 2881 137147 2909 137175
rect 2943 137147 2971 137175
rect 2757 137085 2785 137113
rect 2819 137085 2847 137113
rect 2881 137085 2909 137113
rect 2943 137085 2971 137113
rect 2757 137023 2785 137051
rect 2819 137023 2847 137051
rect 2881 137023 2909 137051
rect 2943 137023 2971 137051
rect 2757 136961 2785 136989
rect 2819 136961 2847 136989
rect 2881 136961 2909 136989
rect 2943 136961 2971 136989
rect 15939 140147 15967 140175
rect 16001 140147 16029 140175
rect 15939 140085 15967 140113
rect 16001 140085 16029 140113
rect 15939 140023 15967 140051
rect 16001 140023 16029 140051
rect 15939 139961 15967 139989
rect 16001 139961 16029 139989
rect 8259 137147 8287 137175
rect 8321 137147 8349 137175
rect 8259 137085 8287 137113
rect 8321 137085 8349 137113
rect 8259 137023 8287 137051
rect 8321 137023 8349 137051
rect 8259 136961 8287 136989
rect 8321 136961 8349 136989
rect 18117 137147 18145 137175
rect 18179 137147 18207 137175
rect 18241 137147 18269 137175
rect 18303 137147 18331 137175
rect 18117 137085 18145 137113
rect 18179 137085 18207 137113
rect 18241 137085 18269 137113
rect 18303 137085 18331 137113
rect 18117 137023 18145 137051
rect 18179 137023 18207 137051
rect 18241 137023 18269 137051
rect 18303 137023 18331 137051
rect 18117 136961 18145 136989
rect 18179 136961 18207 136989
rect 18241 136961 18269 136989
rect 18303 136961 18331 136989
rect 4617 131147 4645 131175
rect 4679 131147 4707 131175
rect 4741 131147 4769 131175
rect 4803 131147 4831 131175
rect 4617 131085 4645 131113
rect 4679 131085 4707 131113
rect 4741 131085 4769 131113
rect 4803 131085 4831 131113
rect 4617 131023 4645 131051
rect 4679 131023 4707 131051
rect 4741 131023 4769 131051
rect 4803 131023 4831 131051
rect 4617 130961 4645 130989
rect 4679 130961 4707 130989
rect 4741 130961 4769 130989
rect 4803 130961 4831 130989
rect 2757 128147 2785 128175
rect 2819 128147 2847 128175
rect 2881 128147 2909 128175
rect 2943 128147 2971 128175
rect 2757 128085 2785 128113
rect 2819 128085 2847 128113
rect 2881 128085 2909 128113
rect 2943 128085 2971 128113
rect 2757 128023 2785 128051
rect 2819 128023 2847 128051
rect 2881 128023 2909 128051
rect 2943 128023 2971 128051
rect 2757 127961 2785 127989
rect 2819 127961 2847 127989
rect 2881 127961 2909 127989
rect 2943 127961 2971 127989
rect 2757 119147 2785 119175
rect 2819 119147 2847 119175
rect 2881 119147 2909 119175
rect 2943 119147 2971 119175
rect 2757 119085 2785 119113
rect 2819 119085 2847 119113
rect 2881 119085 2909 119113
rect 2943 119085 2971 119113
rect 2757 119023 2785 119051
rect 2819 119023 2847 119051
rect 2881 119023 2909 119051
rect 2943 119023 2971 119051
rect 2757 118961 2785 118989
rect 2819 118961 2847 118989
rect 2881 118961 2909 118989
rect 2943 118961 2971 118989
rect -430 110147 -402 110175
rect -368 110147 -340 110175
rect -306 110147 -278 110175
rect -244 110147 -216 110175
rect -430 110085 -402 110113
rect -368 110085 -340 110113
rect -306 110085 -278 110113
rect -244 110085 -216 110113
rect -430 110023 -402 110051
rect -368 110023 -340 110051
rect -306 110023 -278 110051
rect -244 110023 -216 110051
rect -430 109961 -402 109989
rect -368 109961 -340 109989
rect -306 109961 -278 109989
rect -244 109961 -216 109989
rect -430 101147 -402 101175
rect -368 101147 -340 101175
rect -306 101147 -278 101175
rect -244 101147 -216 101175
rect -430 101085 -402 101113
rect -368 101085 -340 101113
rect -306 101085 -278 101113
rect -244 101085 -216 101113
rect -430 101023 -402 101051
rect -368 101023 -340 101051
rect -306 101023 -278 101051
rect -244 101023 -216 101051
rect -430 100961 -402 100989
rect -368 100961 -340 100989
rect -306 100961 -278 100989
rect -244 100961 -216 100989
rect 15939 131147 15967 131175
rect 16001 131147 16029 131175
rect 15939 131085 15967 131113
rect 16001 131085 16029 131113
rect 15939 131023 15967 131051
rect 16001 131023 16029 131051
rect 15939 130961 15967 130989
rect 16001 130961 16029 130989
rect 8259 128147 8287 128175
rect 8321 128147 8349 128175
rect 8259 128085 8287 128113
rect 8321 128085 8349 128113
rect 8259 128023 8287 128051
rect 8321 128023 8349 128051
rect 8259 127961 8287 127989
rect 8321 127961 8349 127989
rect 18117 128147 18145 128175
rect 18179 128147 18207 128175
rect 18241 128147 18269 128175
rect 18303 128147 18331 128175
rect 18117 128085 18145 128113
rect 18179 128085 18207 128113
rect 18241 128085 18269 128113
rect 18303 128085 18331 128113
rect 18117 128023 18145 128051
rect 18179 128023 18207 128051
rect 18241 128023 18269 128051
rect 18303 128023 18331 128051
rect 18117 127961 18145 127989
rect 18179 127961 18207 127989
rect 18241 127961 18269 127989
rect 18303 127961 18331 127989
rect 4617 122147 4645 122175
rect 4679 122147 4707 122175
rect 4741 122147 4769 122175
rect 4803 122147 4831 122175
rect 4617 122085 4645 122113
rect 4679 122085 4707 122113
rect 4741 122085 4769 122113
rect 4803 122085 4831 122113
rect 4617 122023 4645 122051
rect 4679 122023 4707 122051
rect 4741 122023 4769 122051
rect 4803 122023 4831 122051
rect 4617 121961 4645 121989
rect 4679 121961 4707 121989
rect 4741 121961 4769 121989
rect 4803 121961 4831 121989
rect 2757 110147 2785 110175
rect 2819 110147 2847 110175
rect 2881 110147 2909 110175
rect 2943 110147 2971 110175
rect 2757 110085 2785 110113
rect 2819 110085 2847 110113
rect 2881 110085 2909 110113
rect 2943 110085 2971 110113
rect 2757 110023 2785 110051
rect 2819 110023 2847 110051
rect 2881 110023 2909 110051
rect 2943 110023 2971 110051
rect 2757 109961 2785 109989
rect 2819 109961 2847 109989
rect 2881 109961 2909 109989
rect 2943 109961 2971 109989
rect 15939 122147 15967 122175
rect 16001 122147 16029 122175
rect 15939 122085 15967 122113
rect 16001 122085 16029 122113
rect 15939 122023 15967 122051
rect 16001 122023 16029 122051
rect 15939 121961 15967 121989
rect 16001 121961 16029 121989
rect 8259 119147 8287 119175
rect 8321 119147 8349 119175
rect 8259 119085 8287 119113
rect 8321 119085 8349 119113
rect 8259 119023 8287 119051
rect 8321 119023 8349 119051
rect 8259 118961 8287 118989
rect 8321 118961 8349 118989
rect 18117 119147 18145 119175
rect 18179 119147 18207 119175
rect 18241 119147 18269 119175
rect 18303 119147 18331 119175
rect 18117 119085 18145 119113
rect 18179 119085 18207 119113
rect 18241 119085 18269 119113
rect 18303 119085 18331 119113
rect 18117 119023 18145 119051
rect 18179 119023 18207 119051
rect 18241 119023 18269 119051
rect 18303 119023 18331 119051
rect 18117 118961 18145 118989
rect 18179 118961 18207 118989
rect 18241 118961 18269 118989
rect 18303 118961 18331 118989
rect 4617 113147 4645 113175
rect 4679 113147 4707 113175
rect 4741 113147 4769 113175
rect 4803 113147 4831 113175
rect 4617 113085 4645 113113
rect 4679 113085 4707 113113
rect 4741 113085 4769 113113
rect 4803 113085 4831 113113
rect 4617 113023 4645 113051
rect 4679 113023 4707 113051
rect 4741 113023 4769 113051
rect 4803 113023 4831 113051
rect 4617 112961 4645 112989
rect 4679 112961 4707 112989
rect 4741 112961 4769 112989
rect 4803 112961 4831 112989
rect 15939 113147 15967 113175
rect 16001 113147 16029 113175
rect 15939 113085 15967 113113
rect 16001 113085 16029 113113
rect 15939 113023 15967 113051
rect 16001 113023 16029 113051
rect 15939 112961 15967 112989
rect 16001 112961 16029 112989
rect 8259 110147 8287 110175
rect 8321 110147 8349 110175
rect 8259 110085 8287 110113
rect 8321 110085 8349 110113
rect 8259 110023 8287 110051
rect 8321 110023 8349 110051
rect 8259 109961 8287 109989
rect 8321 109961 8349 109989
rect 18117 110147 18145 110175
rect 18179 110147 18207 110175
rect 18241 110147 18269 110175
rect 18303 110147 18331 110175
rect 18117 110085 18145 110113
rect 18179 110085 18207 110113
rect 18241 110085 18269 110113
rect 18303 110085 18331 110113
rect 18117 110023 18145 110051
rect 18179 110023 18207 110051
rect 18241 110023 18269 110051
rect 18303 110023 18331 110051
rect 18117 109961 18145 109989
rect 18179 109961 18207 109989
rect 18241 109961 18269 109989
rect 18303 109961 18331 109989
rect 4617 104147 4645 104175
rect 4679 104147 4707 104175
rect 4741 104147 4769 104175
rect 4803 104147 4831 104175
rect 4617 104085 4645 104113
rect 4679 104085 4707 104113
rect 4741 104085 4769 104113
rect 4803 104085 4831 104113
rect 4617 104023 4645 104051
rect 4679 104023 4707 104051
rect 4741 104023 4769 104051
rect 4803 104023 4831 104051
rect 4617 103961 4645 103989
rect 4679 103961 4707 103989
rect 4741 103961 4769 103989
rect 4803 103961 4831 103989
rect 2757 101147 2785 101175
rect 2819 101147 2847 101175
rect 2881 101147 2909 101175
rect 2943 101147 2971 101175
rect 2757 101085 2785 101113
rect 2819 101085 2847 101113
rect 2881 101085 2909 101113
rect 2943 101085 2971 101113
rect 2757 101023 2785 101051
rect 2819 101023 2847 101051
rect 2881 101023 2909 101051
rect 2943 101023 2971 101051
rect 2757 100961 2785 100989
rect 2819 100961 2847 100989
rect 2881 100961 2909 100989
rect 2943 100961 2971 100989
rect -430 92147 -402 92175
rect -368 92147 -340 92175
rect -306 92147 -278 92175
rect -244 92147 -216 92175
rect -430 92085 -402 92113
rect -368 92085 -340 92113
rect -306 92085 -278 92113
rect -244 92085 -216 92113
rect -430 92023 -402 92051
rect -368 92023 -340 92051
rect -306 92023 -278 92051
rect -244 92023 -216 92051
rect -430 91961 -402 91989
rect -368 91961 -340 91989
rect -306 91961 -278 91989
rect -244 91961 -216 91989
rect 2757 92147 2785 92175
rect 2819 92147 2847 92175
rect 2881 92147 2909 92175
rect 2943 92147 2971 92175
rect 2757 92085 2785 92113
rect 2819 92085 2847 92113
rect 2881 92085 2909 92113
rect 2943 92085 2971 92113
rect 2757 92023 2785 92051
rect 2819 92023 2847 92051
rect 2881 92023 2909 92051
rect 2943 92023 2971 92051
rect 2757 91961 2785 91989
rect 2819 91961 2847 91989
rect 2881 91961 2909 91989
rect 2943 91961 2971 91989
rect -430 83147 -402 83175
rect -368 83147 -340 83175
rect -306 83147 -278 83175
rect -244 83147 -216 83175
rect -430 83085 -402 83113
rect -368 83085 -340 83113
rect -306 83085 -278 83113
rect -244 83085 -216 83113
rect -430 83023 -402 83051
rect -368 83023 -340 83051
rect -306 83023 -278 83051
rect -244 83023 -216 83051
rect -430 82961 -402 82989
rect -368 82961 -340 82989
rect -306 82961 -278 82989
rect -244 82961 -216 82989
rect 2757 83147 2785 83175
rect 2819 83147 2847 83175
rect 2881 83147 2909 83175
rect 2943 83147 2971 83175
rect 2757 83085 2785 83113
rect 2819 83085 2847 83113
rect 2881 83085 2909 83113
rect 2943 83085 2971 83113
rect 2757 83023 2785 83051
rect 2819 83023 2847 83051
rect 2881 83023 2909 83051
rect 2943 83023 2971 83051
rect 2757 82961 2785 82989
rect 2819 82961 2847 82989
rect 2881 82961 2909 82989
rect 2943 82961 2971 82989
rect -430 74147 -402 74175
rect -368 74147 -340 74175
rect -306 74147 -278 74175
rect -244 74147 -216 74175
rect -430 74085 -402 74113
rect -368 74085 -340 74113
rect -306 74085 -278 74113
rect -244 74085 -216 74113
rect -430 74023 -402 74051
rect -368 74023 -340 74051
rect -306 74023 -278 74051
rect -244 74023 -216 74051
rect -430 73961 -402 73989
rect -368 73961 -340 73989
rect -306 73961 -278 73989
rect -244 73961 -216 73989
rect -430 65147 -402 65175
rect -368 65147 -340 65175
rect -306 65147 -278 65175
rect -244 65147 -216 65175
rect -430 65085 -402 65113
rect -368 65085 -340 65113
rect -306 65085 -278 65113
rect -244 65085 -216 65113
rect -430 65023 -402 65051
rect -368 65023 -340 65051
rect -306 65023 -278 65051
rect -244 65023 -216 65051
rect -430 64961 -402 64989
rect -368 64961 -340 64989
rect -306 64961 -278 64989
rect -244 64961 -216 64989
rect -430 56147 -402 56175
rect -368 56147 -340 56175
rect -306 56147 -278 56175
rect -244 56147 -216 56175
rect -430 56085 -402 56113
rect -368 56085 -340 56113
rect -306 56085 -278 56113
rect -244 56085 -216 56113
rect -430 56023 -402 56051
rect -368 56023 -340 56051
rect -306 56023 -278 56051
rect -244 56023 -216 56051
rect -430 55961 -402 55989
rect -368 55961 -340 55989
rect -306 55961 -278 55989
rect -244 55961 -216 55989
rect -430 47147 -402 47175
rect -368 47147 -340 47175
rect -306 47147 -278 47175
rect -244 47147 -216 47175
rect -430 47085 -402 47113
rect -368 47085 -340 47113
rect -306 47085 -278 47113
rect -244 47085 -216 47113
rect -430 47023 -402 47051
rect -368 47023 -340 47051
rect -306 47023 -278 47051
rect -244 47023 -216 47051
rect -430 46961 -402 46989
rect -368 46961 -340 46989
rect -306 46961 -278 46989
rect -244 46961 -216 46989
rect -430 38147 -402 38175
rect -368 38147 -340 38175
rect -306 38147 -278 38175
rect -244 38147 -216 38175
rect -430 38085 -402 38113
rect -368 38085 -340 38113
rect -306 38085 -278 38113
rect -244 38085 -216 38113
rect -430 38023 -402 38051
rect -368 38023 -340 38051
rect -306 38023 -278 38051
rect -244 38023 -216 38051
rect -430 37961 -402 37989
rect -368 37961 -340 37989
rect -306 37961 -278 37989
rect -244 37961 -216 37989
rect -430 29147 -402 29175
rect -368 29147 -340 29175
rect -306 29147 -278 29175
rect -244 29147 -216 29175
rect -430 29085 -402 29113
rect -368 29085 -340 29113
rect -306 29085 -278 29113
rect -244 29085 -216 29113
rect -430 29023 -402 29051
rect -368 29023 -340 29051
rect -306 29023 -278 29051
rect -244 29023 -216 29051
rect -430 28961 -402 28989
rect -368 28961 -340 28989
rect -306 28961 -278 28989
rect -244 28961 -216 28989
rect 15939 104147 15967 104175
rect 16001 104147 16029 104175
rect 15939 104085 15967 104113
rect 16001 104085 16029 104113
rect 15939 104023 15967 104051
rect 16001 104023 16029 104051
rect 15939 103961 15967 103989
rect 16001 103961 16029 103989
rect 8259 101147 8287 101175
rect 8321 101147 8349 101175
rect 8259 101085 8287 101113
rect 8321 101085 8349 101113
rect 8259 101023 8287 101051
rect 8321 101023 8349 101051
rect 8259 100961 8287 100989
rect 8321 100961 8349 100989
rect 18117 101147 18145 101175
rect 18179 101147 18207 101175
rect 18241 101147 18269 101175
rect 18303 101147 18331 101175
rect 18117 101085 18145 101113
rect 18179 101085 18207 101113
rect 18241 101085 18269 101113
rect 18303 101085 18331 101113
rect 18117 101023 18145 101051
rect 18179 101023 18207 101051
rect 18241 101023 18269 101051
rect 18303 101023 18331 101051
rect 18117 100961 18145 100989
rect 18179 100961 18207 100989
rect 18241 100961 18269 100989
rect 18303 100961 18331 100989
rect 4617 95147 4645 95175
rect 4679 95147 4707 95175
rect 4741 95147 4769 95175
rect 4803 95147 4831 95175
rect 4617 95085 4645 95113
rect 4679 95085 4707 95113
rect 4741 95085 4769 95113
rect 4803 95085 4831 95113
rect 4617 95023 4645 95051
rect 4679 95023 4707 95051
rect 4741 95023 4769 95051
rect 4803 95023 4831 95051
rect 4617 94961 4645 94989
rect 4679 94961 4707 94989
rect 4741 94961 4769 94989
rect 4803 94961 4831 94989
rect 15939 95147 15967 95175
rect 16001 95147 16029 95175
rect 15939 95085 15967 95113
rect 16001 95085 16029 95113
rect 15939 95023 15967 95051
rect 16001 95023 16029 95051
rect 15939 94961 15967 94989
rect 16001 94961 16029 94989
rect 8259 92147 8287 92175
rect 8321 92147 8349 92175
rect 8259 92085 8287 92113
rect 8321 92085 8349 92113
rect 8259 92023 8287 92051
rect 8321 92023 8349 92051
rect 8259 91961 8287 91989
rect 8321 91961 8349 91989
rect 18117 92147 18145 92175
rect 18179 92147 18207 92175
rect 18241 92147 18269 92175
rect 18303 92147 18331 92175
rect 18117 92085 18145 92113
rect 18179 92085 18207 92113
rect 18241 92085 18269 92113
rect 18303 92085 18331 92113
rect 18117 92023 18145 92051
rect 18179 92023 18207 92051
rect 18241 92023 18269 92051
rect 18303 92023 18331 92051
rect 18117 91961 18145 91989
rect 18179 91961 18207 91989
rect 18241 91961 18269 91989
rect 18303 91961 18331 91989
rect 4617 86147 4645 86175
rect 4679 86147 4707 86175
rect 4741 86147 4769 86175
rect 4803 86147 4831 86175
rect 4617 86085 4645 86113
rect 4679 86085 4707 86113
rect 4741 86085 4769 86113
rect 4803 86085 4831 86113
rect 4617 86023 4645 86051
rect 4679 86023 4707 86051
rect 4741 86023 4769 86051
rect 4803 86023 4831 86051
rect 4617 85961 4645 85989
rect 4679 85961 4707 85989
rect 4741 85961 4769 85989
rect 4803 85961 4831 85989
rect 15939 86147 15967 86175
rect 16001 86147 16029 86175
rect 15939 86085 15967 86113
rect 16001 86085 16029 86113
rect 15939 86023 15967 86051
rect 16001 86023 16029 86051
rect 15939 85961 15967 85989
rect 16001 85961 16029 85989
rect 8259 83147 8287 83175
rect 8321 83147 8349 83175
rect 8259 83085 8287 83113
rect 8321 83085 8349 83113
rect 8259 83023 8287 83051
rect 8321 83023 8349 83051
rect 8259 82961 8287 82989
rect 8321 82961 8349 82989
rect 18117 83147 18145 83175
rect 18179 83147 18207 83175
rect 18241 83147 18269 83175
rect 18303 83147 18331 83175
rect 18117 83085 18145 83113
rect 18179 83085 18207 83113
rect 18241 83085 18269 83113
rect 18303 83085 18331 83113
rect 18117 83023 18145 83051
rect 18179 83023 18207 83051
rect 18241 83023 18269 83051
rect 18303 83023 18331 83051
rect 18117 82961 18145 82989
rect 18179 82961 18207 82989
rect 18241 82961 18269 82989
rect 18303 82961 18331 82989
rect 4617 77147 4645 77175
rect 4679 77147 4707 77175
rect 4741 77147 4769 77175
rect 4803 77147 4831 77175
rect 4617 77085 4645 77113
rect 4679 77085 4707 77113
rect 4741 77085 4769 77113
rect 4803 77085 4831 77113
rect 4617 77023 4645 77051
rect 4679 77023 4707 77051
rect 4741 77023 4769 77051
rect 4803 77023 4831 77051
rect 4617 76961 4645 76989
rect 4679 76961 4707 76989
rect 4741 76961 4769 76989
rect 4803 76961 4831 76989
rect 2757 74147 2785 74175
rect 2819 74147 2847 74175
rect 2881 74147 2909 74175
rect 2943 74147 2971 74175
rect 2757 74085 2785 74113
rect 2819 74085 2847 74113
rect 2881 74085 2909 74113
rect 2943 74085 2971 74113
rect 2757 74023 2785 74051
rect 2819 74023 2847 74051
rect 2881 74023 2909 74051
rect 2943 74023 2971 74051
rect 2757 73961 2785 73989
rect 2819 73961 2847 73989
rect 2881 73961 2909 73989
rect 2943 73961 2971 73989
rect 15939 77147 15967 77175
rect 16001 77147 16029 77175
rect 15939 77085 15967 77113
rect 16001 77085 16029 77113
rect 15939 77023 15967 77051
rect 16001 77023 16029 77051
rect 15939 76961 15967 76989
rect 16001 76961 16029 76989
rect 8259 74147 8287 74175
rect 8321 74147 8349 74175
rect 8259 74085 8287 74113
rect 8321 74085 8349 74113
rect 8259 74023 8287 74051
rect 8321 74023 8349 74051
rect 8259 73961 8287 73989
rect 8321 73961 8349 73989
rect 18117 74147 18145 74175
rect 18179 74147 18207 74175
rect 18241 74147 18269 74175
rect 18303 74147 18331 74175
rect 18117 74085 18145 74113
rect 18179 74085 18207 74113
rect 18241 74085 18269 74113
rect 18303 74085 18331 74113
rect 18117 74023 18145 74051
rect 18179 74023 18207 74051
rect 18241 74023 18269 74051
rect 18303 74023 18331 74051
rect 18117 73961 18145 73989
rect 18179 73961 18207 73989
rect 18241 73961 18269 73989
rect 18303 73961 18331 73989
rect 4617 68147 4645 68175
rect 4679 68147 4707 68175
rect 4741 68147 4769 68175
rect 4803 68147 4831 68175
rect 4617 68085 4645 68113
rect 4679 68085 4707 68113
rect 4741 68085 4769 68113
rect 4803 68085 4831 68113
rect 4617 68023 4645 68051
rect 4679 68023 4707 68051
rect 4741 68023 4769 68051
rect 4803 68023 4831 68051
rect 4617 67961 4645 67989
rect 4679 67961 4707 67989
rect 4741 67961 4769 67989
rect 4803 67961 4831 67989
rect 2757 65147 2785 65175
rect 2819 65147 2847 65175
rect 2881 65147 2909 65175
rect 2943 65147 2971 65175
rect 2757 65085 2785 65113
rect 2819 65085 2847 65113
rect 2881 65085 2909 65113
rect 2943 65085 2971 65113
rect 2757 65023 2785 65051
rect 2819 65023 2847 65051
rect 2881 65023 2909 65051
rect 2943 65023 2971 65051
rect 2757 64961 2785 64989
rect 2819 64961 2847 64989
rect 2881 64961 2909 64989
rect 2943 64961 2971 64989
rect 15939 68147 15967 68175
rect 16001 68147 16029 68175
rect 15939 68085 15967 68113
rect 16001 68085 16029 68113
rect 15939 68023 15967 68051
rect 16001 68023 16029 68051
rect 15939 67961 15967 67989
rect 16001 67961 16029 67989
rect 8259 65147 8287 65175
rect 8321 65147 8349 65175
rect 8259 65085 8287 65113
rect 8321 65085 8349 65113
rect 8259 65023 8287 65051
rect 8321 65023 8349 65051
rect 8259 64961 8287 64989
rect 8321 64961 8349 64989
rect 18117 65147 18145 65175
rect 18179 65147 18207 65175
rect 18241 65147 18269 65175
rect 18303 65147 18331 65175
rect 18117 65085 18145 65113
rect 18179 65085 18207 65113
rect 18241 65085 18269 65113
rect 18303 65085 18331 65113
rect 18117 65023 18145 65051
rect 18179 65023 18207 65051
rect 18241 65023 18269 65051
rect 18303 65023 18331 65051
rect 18117 64961 18145 64989
rect 18179 64961 18207 64989
rect 18241 64961 18269 64989
rect 18303 64961 18331 64989
rect 4617 59147 4645 59175
rect 4679 59147 4707 59175
rect 4741 59147 4769 59175
rect 4803 59147 4831 59175
rect 4617 59085 4645 59113
rect 4679 59085 4707 59113
rect 4741 59085 4769 59113
rect 4803 59085 4831 59113
rect 4617 59023 4645 59051
rect 4679 59023 4707 59051
rect 4741 59023 4769 59051
rect 4803 59023 4831 59051
rect 4617 58961 4645 58989
rect 4679 58961 4707 58989
rect 4741 58961 4769 58989
rect 4803 58961 4831 58989
rect 2757 56147 2785 56175
rect 2819 56147 2847 56175
rect 2881 56147 2909 56175
rect 2943 56147 2971 56175
rect 2757 56085 2785 56113
rect 2819 56085 2847 56113
rect 2881 56085 2909 56113
rect 2943 56085 2971 56113
rect 2757 56023 2785 56051
rect 2819 56023 2847 56051
rect 2881 56023 2909 56051
rect 2943 56023 2971 56051
rect 2757 55961 2785 55989
rect 2819 55961 2847 55989
rect 2881 55961 2909 55989
rect 2943 55961 2971 55989
rect 15939 59147 15967 59175
rect 16001 59147 16029 59175
rect 15939 59085 15967 59113
rect 16001 59085 16029 59113
rect 15939 59023 15967 59051
rect 16001 59023 16029 59051
rect 15939 58961 15967 58989
rect 16001 58961 16029 58989
rect 8259 56147 8287 56175
rect 8321 56147 8349 56175
rect 8259 56085 8287 56113
rect 8321 56085 8349 56113
rect 8259 56023 8287 56051
rect 8321 56023 8349 56051
rect 8259 55961 8287 55989
rect 8321 55961 8349 55989
rect 18117 56147 18145 56175
rect 18179 56147 18207 56175
rect 18241 56147 18269 56175
rect 18303 56147 18331 56175
rect 18117 56085 18145 56113
rect 18179 56085 18207 56113
rect 18241 56085 18269 56113
rect 18303 56085 18331 56113
rect 18117 56023 18145 56051
rect 18179 56023 18207 56051
rect 18241 56023 18269 56051
rect 18303 56023 18331 56051
rect 18117 55961 18145 55989
rect 18179 55961 18207 55989
rect 18241 55961 18269 55989
rect 18303 55961 18331 55989
rect 4617 50147 4645 50175
rect 4679 50147 4707 50175
rect 4741 50147 4769 50175
rect 4803 50147 4831 50175
rect 4617 50085 4645 50113
rect 4679 50085 4707 50113
rect 4741 50085 4769 50113
rect 4803 50085 4831 50113
rect 4617 50023 4645 50051
rect 4679 50023 4707 50051
rect 4741 50023 4769 50051
rect 4803 50023 4831 50051
rect 4617 49961 4645 49989
rect 4679 49961 4707 49989
rect 4741 49961 4769 49989
rect 4803 49961 4831 49989
rect 2757 47147 2785 47175
rect 2819 47147 2847 47175
rect 2881 47147 2909 47175
rect 2943 47147 2971 47175
rect 2757 47085 2785 47113
rect 2819 47085 2847 47113
rect 2881 47085 2909 47113
rect 2943 47085 2971 47113
rect 2757 47023 2785 47051
rect 2819 47023 2847 47051
rect 2881 47023 2909 47051
rect 2943 47023 2971 47051
rect 2757 46961 2785 46989
rect 2819 46961 2847 46989
rect 2881 46961 2909 46989
rect 2943 46961 2971 46989
rect 15939 50147 15967 50175
rect 16001 50147 16029 50175
rect 15939 50085 15967 50113
rect 16001 50085 16029 50113
rect 15939 50023 15967 50051
rect 16001 50023 16029 50051
rect 15939 49961 15967 49989
rect 16001 49961 16029 49989
rect 8259 47147 8287 47175
rect 8321 47147 8349 47175
rect 8259 47085 8287 47113
rect 8321 47085 8349 47113
rect 8259 47023 8287 47051
rect 8321 47023 8349 47051
rect 8259 46961 8287 46989
rect 8321 46961 8349 46989
rect 18117 47147 18145 47175
rect 18179 47147 18207 47175
rect 18241 47147 18269 47175
rect 18303 47147 18331 47175
rect 18117 47085 18145 47113
rect 18179 47085 18207 47113
rect 18241 47085 18269 47113
rect 18303 47085 18331 47113
rect 18117 47023 18145 47051
rect 18179 47023 18207 47051
rect 18241 47023 18269 47051
rect 18303 47023 18331 47051
rect 18117 46961 18145 46989
rect 18179 46961 18207 46989
rect 18241 46961 18269 46989
rect 18303 46961 18331 46989
rect 4617 41147 4645 41175
rect 4679 41147 4707 41175
rect 4741 41147 4769 41175
rect 4803 41147 4831 41175
rect 4617 41085 4645 41113
rect 4679 41085 4707 41113
rect 4741 41085 4769 41113
rect 4803 41085 4831 41113
rect 4617 41023 4645 41051
rect 4679 41023 4707 41051
rect 4741 41023 4769 41051
rect 4803 41023 4831 41051
rect 4617 40961 4645 40989
rect 4679 40961 4707 40989
rect 4741 40961 4769 40989
rect 4803 40961 4831 40989
rect 2757 38147 2785 38175
rect 2819 38147 2847 38175
rect 2881 38147 2909 38175
rect 2943 38147 2971 38175
rect 2757 38085 2785 38113
rect 2819 38085 2847 38113
rect 2881 38085 2909 38113
rect 2943 38085 2971 38113
rect 2757 38023 2785 38051
rect 2819 38023 2847 38051
rect 2881 38023 2909 38051
rect 2943 38023 2971 38051
rect 2757 37961 2785 37989
rect 2819 37961 2847 37989
rect 2881 37961 2909 37989
rect 2943 37961 2971 37989
rect 2757 29147 2785 29175
rect 2819 29147 2847 29175
rect 2881 29147 2909 29175
rect 2943 29147 2971 29175
rect 2757 29085 2785 29113
rect 2819 29085 2847 29113
rect 2881 29085 2909 29113
rect 2943 29085 2971 29113
rect 2757 29023 2785 29051
rect 2819 29023 2847 29051
rect 2881 29023 2909 29051
rect 2943 29023 2971 29051
rect 2757 28961 2785 28989
rect 2819 28961 2847 28989
rect 2881 28961 2909 28989
rect 2943 28961 2971 28989
rect -430 20147 -402 20175
rect -368 20147 -340 20175
rect -306 20147 -278 20175
rect -244 20147 -216 20175
rect -430 20085 -402 20113
rect -368 20085 -340 20113
rect -306 20085 -278 20113
rect -244 20085 -216 20113
rect -430 20023 -402 20051
rect -368 20023 -340 20051
rect -306 20023 -278 20051
rect -244 20023 -216 20051
rect -430 19961 -402 19989
rect -368 19961 -340 19989
rect -306 19961 -278 19989
rect -244 19961 -216 19989
rect 15939 41147 15967 41175
rect 16001 41147 16029 41175
rect 15939 41085 15967 41113
rect 16001 41085 16029 41113
rect 15939 41023 15967 41051
rect 16001 41023 16029 41051
rect 15939 40961 15967 40989
rect 16001 40961 16029 40989
rect 8259 38147 8287 38175
rect 8321 38147 8349 38175
rect 8259 38085 8287 38113
rect 8321 38085 8349 38113
rect 8259 38023 8287 38051
rect 8321 38023 8349 38051
rect 8259 37961 8287 37989
rect 8321 37961 8349 37989
rect 18117 38147 18145 38175
rect 18179 38147 18207 38175
rect 18241 38147 18269 38175
rect 18303 38147 18331 38175
rect 18117 38085 18145 38113
rect 18179 38085 18207 38113
rect 18241 38085 18269 38113
rect 18303 38085 18331 38113
rect 18117 38023 18145 38051
rect 18179 38023 18207 38051
rect 18241 38023 18269 38051
rect 18303 38023 18331 38051
rect 18117 37961 18145 37989
rect 18179 37961 18207 37989
rect 18241 37961 18269 37989
rect 18303 37961 18331 37989
rect 4617 32147 4645 32175
rect 4679 32147 4707 32175
rect 4741 32147 4769 32175
rect 4803 32147 4831 32175
rect 4617 32085 4645 32113
rect 4679 32085 4707 32113
rect 4741 32085 4769 32113
rect 4803 32085 4831 32113
rect 4617 32023 4645 32051
rect 4679 32023 4707 32051
rect 4741 32023 4769 32051
rect 4803 32023 4831 32051
rect 4617 31961 4645 31989
rect 4679 31961 4707 31989
rect 4741 31961 4769 31989
rect 4803 31961 4831 31989
rect 15939 32147 15967 32175
rect 16001 32147 16029 32175
rect 15939 32085 15967 32113
rect 16001 32085 16029 32113
rect 15939 32023 15967 32051
rect 16001 32023 16029 32051
rect 15939 31961 15967 31989
rect 16001 31961 16029 31989
rect 8259 29147 8287 29175
rect 8321 29147 8349 29175
rect 8259 29085 8287 29113
rect 8321 29085 8349 29113
rect 8259 29023 8287 29051
rect 8321 29023 8349 29051
rect 8259 28961 8287 28989
rect 8321 28961 8349 28989
rect 18117 29147 18145 29175
rect 18179 29147 18207 29175
rect 18241 29147 18269 29175
rect 18303 29147 18331 29175
rect 18117 29085 18145 29113
rect 18179 29085 18207 29113
rect 18241 29085 18269 29113
rect 18303 29085 18331 29113
rect 18117 29023 18145 29051
rect 18179 29023 18207 29051
rect 18241 29023 18269 29051
rect 18303 29023 18331 29051
rect 18117 28961 18145 28989
rect 18179 28961 18207 28989
rect 18241 28961 18269 28989
rect 18303 28961 18331 28989
rect 4617 23147 4645 23175
rect 4679 23147 4707 23175
rect 4741 23147 4769 23175
rect 4803 23147 4831 23175
rect 4617 23085 4645 23113
rect 4679 23085 4707 23113
rect 4741 23085 4769 23113
rect 4803 23085 4831 23113
rect 4617 23023 4645 23051
rect 4679 23023 4707 23051
rect 4741 23023 4769 23051
rect 4803 23023 4831 23051
rect 4617 22961 4645 22989
rect 4679 22961 4707 22989
rect 4741 22961 4769 22989
rect 4803 22961 4831 22989
rect 2757 20147 2785 20175
rect 2819 20147 2847 20175
rect 2881 20147 2909 20175
rect 2943 20147 2971 20175
rect 2757 20085 2785 20113
rect 2819 20085 2847 20113
rect 2881 20085 2909 20113
rect 2943 20085 2971 20113
rect 2757 20023 2785 20051
rect 2819 20023 2847 20051
rect 2881 20023 2909 20051
rect 2943 20023 2971 20051
rect 2757 19961 2785 19989
rect 2819 19961 2847 19989
rect 2881 19961 2909 19989
rect 2943 19961 2971 19989
rect -430 11147 -402 11175
rect -368 11147 -340 11175
rect -306 11147 -278 11175
rect -244 11147 -216 11175
rect -430 11085 -402 11113
rect -368 11085 -340 11113
rect -306 11085 -278 11113
rect -244 11085 -216 11113
rect -430 11023 -402 11051
rect -368 11023 -340 11051
rect -306 11023 -278 11051
rect -244 11023 -216 11051
rect -430 10961 -402 10989
rect -368 10961 -340 10989
rect -306 10961 -278 10989
rect -244 10961 -216 10989
rect -430 2147 -402 2175
rect -368 2147 -340 2175
rect -306 2147 -278 2175
rect -244 2147 -216 2175
rect -430 2085 -402 2113
rect -368 2085 -340 2113
rect -306 2085 -278 2113
rect -244 2085 -216 2113
rect -430 2023 -402 2051
rect -368 2023 -340 2051
rect -306 2023 -278 2051
rect -244 2023 -216 2051
rect -430 1961 -402 1989
rect -368 1961 -340 1989
rect -306 1961 -278 1989
rect -244 1961 -216 1989
rect -430 -108 -402 -80
rect -368 -108 -340 -80
rect -306 -108 -278 -80
rect -244 -108 -216 -80
rect -430 -170 -402 -142
rect -368 -170 -340 -142
rect -306 -170 -278 -142
rect -244 -170 -216 -142
rect -430 -232 -402 -204
rect -368 -232 -340 -204
rect -306 -232 -278 -204
rect -244 -232 -216 -204
rect -430 -294 -402 -266
rect -368 -294 -340 -266
rect -306 -294 -278 -266
rect -244 -294 -216 -266
rect 2757 11147 2785 11175
rect 2819 11147 2847 11175
rect 2881 11147 2909 11175
rect 2943 11147 2971 11175
rect 2757 11085 2785 11113
rect 2819 11085 2847 11113
rect 2881 11085 2909 11113
rect 2943 11085 2971 11113
rect 2757 11023 2785 11051
rect 2819 11023 2847 11051
rect 2881 11023 2909 11051
rect 2943 11023 2971 11051
rect 2757 10961 2785 10989
rect 2819 10961 2847 10989
rect 2881 10961 2909 10989
rect 2943 10961 2971 10989
rect 15939 23147 15967 23175
rect 16001 23147 16029 23175
rect 15939 23085 15967 23113
rect 16001 23085 16029 23113
rect 15939 23023 15967 23051
rect 16001 23023 16029 23051
rect 15939 22961 15967 22989
rect 16001 22961 16029 22989
rect 8259 20147 8287 20175
rect 8321 20147 8349 20175
rect 8259 20085 8287 20113
rect 8321 20085 8349 20113
rect 8259 20023 8287 20051
rect 8321 20023 8349 20051
rect 8259 19961 8287 19989
rect 8321 19961 8349 19989
rect 18117 20147 18145 20175
rect 18179 20147 18207 20175
rect 18241 20147 18269 20175
rect 18303 20147 18331 20175
rect 18117 20085 18145 20113
rect 18179 20085 18207 20113
rect 18241 20085 18269 20113
rect 18303 20085 18331 20113
rect 18117 20023 18145 20051
rect 18179 20023 18207 20051
rect 18241 20023 18269 20051
rect 18303 20023 18331 20051
rect 18117 19961 18145 19989
rect 18179 19961 18207 19989
rect 18241 19961 18269 19989
rect 18303 19961 18331 19989
rect 4617 14147 4645 14175
rect 4679 14147 4707 14175
rect 4741 14147 4769 14175
rect 4803 14147 4831 14175
rect 4617 14085 4645 14113
rect 4679 14085 4707 14113
rect 4741 14085 4769 14113
rect 4803 14085 4831 14113
rect 4617 14023 4645 14051
rect 4679 14023 4707 14051
rect 4741 14023 4769 14051
rect 4803 14023 4831 14051
rect 4617 13961 4645 13989
rect 4679 13961 4707 13989
rect 4741 13961 4769 13989
rect 4803 13961 4831 13989
rect 15939 14147 15967 14175
rect 16001 14147 16029 14175
rect 15939 14085 15967 14113
rect 16001 14085 16029 14113
rect 15939 14023 15967 14051
rect 16001 14023 16029 14051
rect 15939 13961 15967 13989
rect 16001 13961 16029 13989
rect 8259 11147 8287 11175
rect 8321 11147 8349 11175
rect 8259 11085 8287 11113
rect 8321 11085 8349 11113
rect 8259 11023 8287 11051
rect 8321 11023 8349 11051
rect 8259 10961 8287 10989
rect 8321 10961 8349 10989
rect 18117 11147 18145 11175
rect 18179 11147 18207 11175
rect 18241 11147 18269 11175
rect 18303 11147 18331 11175
rect 18117 11085 18145 11113
rect 18179 11085 18207 11113
rect 18241 11085 18269 11113
rect 18303 11085 18331 11113
rect 18117 11023 18145 11051
rect 18179 11023 18207 11051
rect 18241 11023 18269 11051
rect 18303 11023 18331 11051
rect 18117 10961 18145 10989
rect 18179 10961 18207 10989
rect 18241 10961 18269 10989
rect 18303 10961 18331 10989
rect 4617 5147 4645 5175
rect 4679 5147 4707 5175
rect 4741 5147 4769 5175
rect 4803 5147 4831 5175
rect 4617 5085 4645 5113
rect 4679 5085 4707 5113
rect 4741 5085 4769 5113
rect 4803 5085 4831 5113
rect 4617 5023 4645 5051
rect 4679 5023 4707 5051
rect 4741 5023 4769 5051
rect 4803 5023 4831 5051
rect 4617 4961 4645 4989
rect 4679 4961 4707 4989
rect 4741 4961 4769 4989
rect 4803 4961 4831 4989
rect 2757 2147 2785 2175
rect 2819 2147 2847 2175
rect 2881 2147 2909 2175
rect 2943 2147 2971 2175
rect 2757 2085 2785 2113
rect 2819 2085 2847 2113
rect 2881 2085 2909 2113
rect 2943 2085 2971 2113
rect 2757 2023 2785 2051
rect 2819 2023 2847 2051
rect 2881 2023 2909 2051
rect 2943 2023 2971 2051
rect 2757 1961 2785 1989
rect 2819 1961 2847 1989
rect 2881 1961 2909 1989
rect 2943 1961 2971 1989
rect 2757 -108 2785 -80
rect 2819 -108 2847 -80
rect 2881 -108 2909 -80
rect 2943 -108 2971 -80
rect 2757 -170 2785 -142
rect 2819 -170 2847 -142
rect 2881 -170 2909 -142
rect 2943 -170 2971 -142
rect 2757 -232 2785 -204
rect 2819 -232 2847 -204
rect 2881 -232 2909 -204
rect 2943 -232 2971 -204
rect 2757 -294 2785 -266
rect 2819 -294 2847 -266
rect 2881 -294 2909 -266
rect 2943 -294 2971 -266
rect -910 -588 -882 -560
rect -848 -588 -820 -560
rect -786 -588 -758 -560
rect -724 -588 -696 -560
rect -910 -650 -882 -622
rect -848 -650 -820 -622
rect -786 -650 -758 -622
rect -724 -650 -696 -622
rect -910 -712 -882 -684
rect -848 -712 -820 -684
rect -786 -712 -758 -684
rect -724 -712 -696 -684
rect -910 -774 -882 -746
rect -848 -774 -820 -746
rect -786 -774 -758 -746
rect -724 -774 -696 -746
rect 15939 5147 15967 5175
rect 16001 5147 16029 5175
rect 15939 5085 15967 5113
rect 16001 5085 16029 5113
rect 15939 5023 15967 5051
rect 16001 5023 16029 5051
rect 15939 4961 15967 4989
rect 16001 4961 16029 4989
rect 4617 -588 4645 -560
rect 4679 -588 4707 -560
rect 4741 -588 4769 -560
rect 4803 -588 4831 -560
rect 4617 -650 4645 -622
rect 4679 -650 4707 -622
rect 4741 -650 4769 -622
rect 4803 -650 4831 -622
rect 4617 -712 4645 -684
rect 4679 -712 4707 -684
rect 4741 -712 4769 -684
rect 4803 -712 4831 -684
rect 4617 -774 4645 -746
rect 4679 -774 4707 -746
rect 4741 -774 4769 -746
rect 4803 -774 4831 -746
rect 18117 2147 18145 2175
rect 18179 2147 18207 2175
rect 18241 2147 18269 2175
rect 18303 2147 18331 2175
rect 18117 2085 18145 2113
rect 18179 2085 18207 2113
rect 18241 2085 18269 2113
rect 18303 2085 18331 2113
rect 18117 2023 18145 2051
rect 18179 2023 18207 2051
rect 18241 2023 18269 2051
rect 18303 2023 18331 2051
rect 18117 1961 18145 1989
rect 18179 1961 18207 1989
rect 18241 1961 18269 1989
rect 18303 1961 18331 1989
rect 18117 -108 18145 -80
rect 18179 -108 18207 -80
rect 18241 -108 18269 -80
rect 18303 -108 18331 -80
rect 18117 -170 18145 -142
rect 18179 -170 18207 -142
rect 18241 -170 18269 -142
rect 18303 -170 18331 -142
rect 18117 -232 18145 -204
rect 18179 -232 18207 -204
rect 18241 -232 18269 -204
rect 18303 -232 18331 -204
rect 18117 -294 18145 -266
rect 18179 -294 18207 -266
rect 18241 -294 18269 -266
rect 18303 -294 18331 -266
rect 19977 299058 20005 299086
rect 20039 299058 20067 299086
rect 20101 299058 20129 299086
rect 20163 299058 20191 299086
rect 19977 298996 20005 299024
rect 20039 298996 20067 299024
rect 20101 298996 20129 299024
rect 20163 298996 20191 299024
rect 19977 298934 20005 298962
rect 20039 298934 20067 298962
rect 20101 298934 20129 298962
rect 20163 298934 20191 298962
rect 19977 298872 20005 298900
rect 20039 298872 20067 298900
rect 20101 298872 20129 298900
rect 20163 298872 20191 298900
rect 19977 293147 20005 293175
rect 20039 293147 20067 293175
rect 20101 293147 20129 293175
rect 20163 293147 20191 293175
rect 19977 293085 20005 293113
rect 20039 293085 20067 293113
rect 20101 293085 20129 293113
rect 20163 293085 20191 293113
rect 19977 293023 20005 293051
rect 20039 293023 20067 293051
rect 20101 293023 20129 293051
rect 20163 293023 20191 293051
rect 19977 292961 20005 292989
rect 20039 292961 20067 292989
rect 20101 292961 20129 292989
rect 20163 292961 20191 292989
rect 19977 284147 20005 284175
rect 20039 284147 20067 284175
rect 20101 284147 20129 284175
rect 20163 284147 20191 284175
rect 19977 284085 20005 284113
rect 20039 284085 20067 284113
rect 20101 284085 20129 284113
rect 20163 284085 20191 284113
rect 19977 284023 20005 284051
rect 20039 284023 20067 284051
rect 20101 284023 20129 284051
rect 20163 284023 20191 284051
rect 19977 283961 20005 283989
rect 20039 283961 20067 283989
rect 20101 283961 20129 283989
rect 20163 283961 20191 283989
rect 19977 275147 20005 275175
rect 20039 275147 20067 275175
rect 20101 275147 20129 275175
rect 20163 275147 20191 275175
rect 19977 275085 20005 275113
rect 20039 275085 20067 275113
rect 20101 275085 20129 275113
rect 20163 275085 20191 275113
rect 19977 275023 20005 275051
rect 20039 275023 20067 275051
rect 20101 275023 20129 275051
rect 20163 275023 20191 275051
rect 19977 274961 20005 274989
rect 20039 274961 20067 274989
rect 20101 274961 20129 274989
rect 20163 274961 20191 274989
rect 19977 266147 20005 266175
rect 20039 266147 20067 266175
rect 20101 266147 20129 266175
rect 20163 266147 20191 266175
rect 19977 266085 20005 266113
rect 20039 266085 20067 266113
rect 20101 266085 20129 266113
rect 20163 266085 20191 266113
rect 19977 266023 20005 266051
rect 20039 266023 20067 266051
rect 20101 266023 20129 266051
rect 20163 266023 20191 266051
rect 19977 265961 20005 265989
rect 20039 265961 20067 265989
rect 20101 265961 20129 265989
rect 20163 265961 20191 265989
rect 19977 257147 20005 257175
rect 20039 257147 20067 257175
rect 20101 257147 20129 257175
rect 20163 257147 20191 257175
rect 19977 257085 20005 257113
rect 20039 257085 20067 257113
rect 20101 257085 20129 257113
rect 20163 257085 20191 257113
rect 19977 257023 20005 257051
rect 20039 257023 20067 257051
rect 20101 257023 20129 257051
rect 20163 257023 20191 257051
rect 19977 256961 20005 256989
rect 20039 256961 20067 256989
rect 20101 256961 20129 256989
rect 20163 256961 20191 256989
rect 19977 248147 20005 248175
rect 20039 248147 20067 248175
rect 20101 248147 20129 248175
rect 20163 248147 20191 248175
rect 19977 248085 20005 248113
rect 20039 248085 20067 248113
rect 20101 248085 20129 248113
rect 20163 248085 20191 248113
rect 19977 248023 20005 248051
rect 20039 248023 20067 248051
rect 20101 248023 20129 248051
rect 20163 248023 20191 248051
rect 19977 247961 20005 247989
rect 20039 247961 20067 247989
rect 20101 247961 20129 247989
rect 20163 247961 20191 247989
rect 19977 239147 20005 239175
rect 20039 239147 20067 239175
rect 20101 239147 20129 239175
rect 20163 239147 20191 239175
rect 19977 239085 20005 239113
rect 20039 239085 20067 239113
rect 20101 239085 20129 239113
rect 20163 239085 20191 239113
rect 19977 239023 20005 239051
rect 20039 239023 20067 239051
rect 20101 239023 20129 239051
rect 20163 239023 20191 239051
rect 19977 238961 20005 238989
rect 20039 238961 20067 238989
rect 20101 238961 20129 238989
rect 20163 238961 20191 238989
rect 19977 230147 20005 230175
rect 20039 230147 20067 230175
rect 20101 230147 20129 230175
rect 20163 230147 20191 230175
rect 19977 230085 20005 230113
rect 20039 230085 20067 230113
rect 20101 230085 20129 230113
rect 20163 230085 20191 230113
rect 19977 230023 20005 230051
rect 20039 230023 20067 230051
rect 20101 230023 20129 230051
rect 20163 230023 20191 230051
rect 19977 229961 20005 229989
rect 20039 229961 20067 229989
rect 20101 229961 20129 229989
rect 20163 229961 20191 229989
rect 19977 221147 20005 221175
rect 20039 221147 20067 221175
rect 20101 221147 20129 221175
rect 20163 221147 20191 221175
rect 19977 221085 20005 221113
rect 20039 221085 20067 221113
rect 20101 221085 20129 221113
rect 20163 221085 20191 221113
rect 19977 221023 20005 221051
rect 20039 221023 20067 221051
rect 20101 221023 20129 221051
rect 20163 221023 20191 221051
rect 19977 220961 20005 220989
rect 20039 220961 20067 220989
rect 20101 220961 20129 220989
rect 20163 220961 20191 220989
rect 19977 212147 20005 212175
rect 20039 212147 20067 212175
rect 20101 212147 20129 212175
rect 20163 212147 20191 212175
rect 19977 212085 20005 212113
rect 20039 212085 20067 212113
rect 20101 212085 20129 212113
rect 20163 212085 20191 212113
rect 19977 212023 20005 212051
rect 20039 212023 20067 212051
rect 20101 212023 20129 212051
rect 20163 212023 20191 212051
rect 19977 211961 20005 211989
rect 20039 211961 20067 211989
rect 20101 211961 20129 211989
rect 20163 211961 20191 211989
rect 19977 203147 20005 203175
rect 20039 203147 20067 203175
rect 20101 203147 20129 203175
rect 20163 203147 20191 203175
rect 19977 203085 20005 203113
rect 20039 203085 20067 203113
rect 20101 203085 20129 203113
rect 20163 203085 20191 203113
rect 19977 203023 20005 203051
rect 20039 203023 20067 203051
rect 20101 203023 20129 203051
rect 20163 203023 20191 203051
rect 19977 202961 20005 202989
rect 20039 202961 20067 202989
rect 20101 202961 20129 202989
rect 20163 202961 20191 202989
rect 19977 194147 20005 194175
rect 20039 194147 20067 194175
rect 20101 194147 20129 194175
rect 20163 194147 20191 194175
rect 19977 194085 20005 194113
rect 20039 194085 20067 194113
rect 20101 194085 20129 194113
rect 20163 194085 20191 194113
rect 19977 194023 20005 194051
rect 20039 194023 20067 194051
rect 20101 194023 20129 194051
rect 20163 194023 20191 194051
rect 19977 193961 20005 193989
rect 20039 193961 20067 193989
rect 20101 193961 20129 193989
rect 20163 193961 20191 193989
rect 19977 185147 20005 185175
rect 20039 185147 20067 185175
rect 20101 185147 20129 185175
rect 20163 185147 20191 185175
rect 19977 185085 20005 185113
rect 20039 185085 20067 185113
rect 20101 185085 20129 185113
rect 20163 185085 20191 185113
rect 19977 185023 20005 185051
rect 20039 185023 20067 185051
rect 20101 185023 20129 185051
rect 20163 185023 20191 185051
rect 19977 184961 20005 184989
rect 20039 184961 20067 184989
rect 20101 184961 20129 184989
rect 20163 184961 20191 184989
rect 19977 176147 20005 176175
rect 20039 176147 20067 176175
rect 20101 176147 20129 176175
rect 20163 176147 20191 176175
rect 19977 176085 20005 176113
rect 20039 176085 20067 176113
rect 20101 176085 20129 176113
rect 20163 176085 20191 176113
rect 19977 176023 20005 176051
rect 20039 176023 20067 176051
rect 20101 176023 20129 176051
rect 20163 176023 20191 176051
rect 19977 175961 20005 175989
rect 20039 175961 20067 175989
rect 20101 175961 20129 175989
rect 20163 175961 20191 175989
rect 33477 298578 33505 298606
rect 33539 298578 33567 298606
rect 33601 298578 33629 298606
rect 33663 298578 33691 298606
rect 33477 298516 33505 298544
rect 33539 298516 33567 298544
rect 33601 298516 33629 298544
rect 33663 298516 33691 298544
rect 33477 298454 33505 298482
rect 33539 298454 33567 298482
rect 33601 298454 33629 298482
rect 33663 298454 33691 298482
rect 33477 298392 33505 298420
rect 33539 298392 33567 298420
rect 33601 298392 33629 298420
rect 33663 298392 33691 298420
rect 33477 290147 33505 290175
rect 33539 290147 33567 290175
rect 33601 290147 33629 290175
rect 33663 290147 33691 290175
rect 33477 290085 33505 290113
rect 33539 290085 33567 290113
rect 33601 290085 33629 290113
rect 33663 290085 33691 290113
rect 33477 290023 33505 290051
rect 33539 290023 33567 290051
rect 33601 290023 33629 290051
rect 33663 290023 33691 290051
rect 33477 289961 33505 289989
rect 33539 289961 33567 289989
rect 33601 289961 33629 289989
rect 33663 289961 33691 289989
rect 33477 281147 33505 281175
rect 33539 281147 33567 281175
rect 33601 281147 33629 281175
rect 33663 281147 33691 281175
rect 33477 281085 33505 281113
rect 33539 281085 33567 281113
rect 33601 281085 33629 281113
rect 33663 281085 33691 281113
rect 33477 281023 33505 281051
rect 33539 281023 33567 281051
rect 33601 281023 33629 281051
rect 33663 281023 33691 281051
rect 33477 280961 33505 280989
rect 33539 280961 33567 280989
rect 33601 280961 33629 280989
rect 33663 280961 33691 280989
rect 33477 272147 33505 272175
rect 33539 272147 33567 272175
rect 33601 272147 33629 272175
rect 33663 272147 33691 272175
rect 33477 272085 33505 272113
rect 33539 272085 33567 272113
rect 33601 272085 33629 272113
rect 33663 272085 33691 272113
rect 33477 272023 33505 272051
rect 33539 272023 33567 272051
rect 33601 272023 33629 272051
rect 33663 272023 33691 272051
rect 33477 271961 33505 271989
rect 33539 271961 33567 271989
rect 33601 271961 33629 271989
rect 33663 271961 33691 271989
rect 33477 263147 33505 263175
rect 33539 263147 33567 263175
rect 33601 263147 33629 263175
rect 33663 263147 33691 263175
rect 33477 263085 33505 263113
rect 33539 263085 33567 263113
rect 33601 263085 33629 263113
rect 33663 263085 33691 263113
rect 33477 263023 33505 263051
rect 33539 263023 33567 263051
rect 33601 263023 33629 263051
rect 33663 263023 33691 263051
rect 33477 262961 33505 262989
rect 33539 262961 33567 262989
rect 33601 262961 33629 262989
rect 33663 262961 33691 262989
rect 33477 254147 33505 254175
rect 33539 254147 33567 254175
rect 33601 254147 33629 254175
rect 33663 254147 33691 254175
rect 33477 254085 33505 254113
rect 33539 254085 33567 254113
rect 33601 254085 33629 254113
rect 33663 254085 33691 254113
rect 33477 254023 33505 254051
rect 33539 254023 33567 254051
rect 33601 254023 33629 254051
rect 33663 254023 33691 254051
rect 33477 253961 33505 253989
rect 33539 253961 33567 253989
rect 33601 253961 33629 253989
rect 33663 253961 33691 253989
rect 33477 245147 33505 245175
rect 33539 245147 33567 245175
rect 33601 245147 33629 245175
rect 33663 245147 33691 245175
rect 33477 245085 33505 245113
rect 33539 245085 33567 245113
rect 33601 245085 33629 245113
rect 33663 245085 33691 245113
rect 33477 245023 33505 245051
rect 33539 245023 33567 245051
rect 33601 245023 33629 245051
rect 33663 245023 33691 245051
rect 33477 244961 33505 244989
rect 33539 244961 33567 244989
rect 33601 244961 33629 244989
rect 33663 244961 33691 244989
rect 33477 236147 33505 236175
rect 33539 236147 33567 236175
rect 33601 236147 33629 236175
rect 33663 236147 33691 236175
rect 33477 236085 33505 236113
rect 33539 236085 33567 236113
rect 33601 236085 33629 236113
rect 33663 236085 33691 236113
rect 33477 236023 33505 236051
rect 33539 236023 33567 236051
rect 33601 236023 33629 236051
rect 33663 236023 33691 236051
rect 33477 235961 33505 235989
rect 33539 235961 33567 235989
rect 33601 235961 33629 235989
rect 33663 235961 33691 235989
rect 33477 227147 33505 227175
rect 33539 227147 33567 227175
rect 33601 227147 33629 227175
rect 33663 227147 33691 227175
rect 33477 227085 33505 227113
rect 33539 227085 33567 227113
rect 33601 227085 33629 227113
rect 33663 227085 33691 227113
rect 33477 227023 33505 227051
rect 33539 227023 33567 227051
rect 33601 227023 33629 227051
rect 33663 227023 33691 227051
rect 33477 226961 33505 226989
rect 33539 226961 33567 226989
rect 33601 226961 33629 226989
rect 33663 226961 33691 226989
rect 33477 218147 33505 218175
rect 33539 218147 33567 218175
rect 33601 218147 33629 218175
rect 33663 218147 33691 218175
rect 33477 218085 33505 218113
rect 33539 218085 33567 218113
rect 33601 218085 33629 218113
rect 33663 218085 33691 218113
rect 33477 218023 33505 218051
rect 33539 218023 33567 218051
rect 33601 218023 33629 218051
rect 33663 218023 33691 218051
rect 33477 217961 33505 217989
rect 33539 217961 33567 217989
rect 33601 217961 33629 217989
rect 33663 217961 33691 217989
rect 33477 209147 33505 209175
rect 33539 209147 33567 209175
rect 33601 209147 33629 209175
rect 33663 209147 33691 209175
rect 33477 209085 33505 209113
rect 33539 209085 33567 209113
rect 33601 209085 33629 209113
rect 33663 209085 33691 209113
rect 33477 209023 33505 209051
rect 33539 209023 33567 209051
rect 33601 209023 33629 209051
rect 33663 209023 33691 209051
rect 33477 208961 33505 208989
rect 33539 208961 33567 208989
rect 33601 208961 33629 208989
rect 33663 208961 33691 208989
rect 33477 200147 33505 200175
rect 33539 200147 33567 200175
rect 33601 200147 33629 200175
rect 33663 200147 33691 200175
rect 33477 200085 33505 200113
rect 33539 200085 33567 200113
rect 33601 200085 33629 200113
rect 33663 200085 33691 200113
rect 33477 200023 33505 200051
rect 33539 200023 33567 200051
rect 33601 200023 33629 200051
rect 33663 200023 33691 200051
rect 33477 199961 33505 199989
rect 33539 199961 33567 199989
rect 33601 199961 33629 199989
rect 33663 199961 33691 199989
rect 33477 191147 33505 191175
rect 33539 191147 33567 191175
rect 33601 191147 33629 191175
rect 33663 191147 33691 191175
rect 33477 191085 33505 191113
rect 33539 191085 33567 191113
rect 33601 191085 33629 191113
rect 33663 191085 33691 191113
rect 33477 191023 33505 191051
rect 33539 191023 33567 191051
rect 33601 191023 33629 191051
rect 33663 191023 33691 191051
rect 33477 190961 33505 190989
rect 33539 190961 33567 190989
rect 33601 190961 33629 190989
rect 33663 190961 33691 190989
rect 33477 182147 33505 182175
rect 33539 182147 33567 182175
rect 33601 182147 33629 182175
rect 33663 182147 33691 182175
rect 33477 182085 33505 182113
rect 33539 182085 33567 182113
rect 33601 182085 33629 182113
rect 33663 182085 33691 182113
rect 33477 182023 33505 182051
rect 33539 182023 33567 182051
rect 33601 182023 33629 182051
rect 33663 182023 33691 182051
rect 33477 181961 33505 181989
rect 33539 181961 33567 181989
rect 33601 181961 33629 181989
rect 33663 181961 33691 181989
rect 23619 173147 23647 173175
rect 23681 173147 23709 173175
rect 23619 173085 23647 173113
rect 23681 173085 23709 173113
rect 23619 173023 23647 173051
rect 23681 173023 23709 173051
rect 23619 172961 23647 172989
rect 23681 172961 23709 172989
rect 33477 173147 33505 173175
rect 33539 173147 33567 173175
rect 33601 173147 33629 173175
rect 33663 173147 33691 173175
rect 33477 173085 33505 173113
rect 33539 173085 33567 173113
rect 33601 173085 33629 173113
rect 33663 173085 33691 173113
rect 33477 173023 33505 173051
rect 33539 173023 33567 173051
rect 33601 173023 33629 173051
rect 33663 173023 33691 173051
rect 33477 172961 33505 172989
rect 33539 172961 33567 172989
rect 33601 172961 33629 172989
rect 33663 172961 33691 172989
rect 19977 167147 20005 167175
rect 20039 167147 20067 167175
rect 20101 167147 20129 167175
rect 20163 167147 20191 167175
rect 19977 167085 20005 167113
rect 20039 167085 20067 167113
rect 20101 167085 20129 167113
rect 20163 167085 20191 167113
rect 19977 167023 20005 167051
rect 20039 167023 20067 167051
rect 20101 167023 20129 167051
rect 20163 167023 20191 167051
rect 19977 166961 20005 166989
rect 20039 166961 20067 166989
rect 20101 166961 20129 166989
rect 20163 166961 20191 166989
rect 31299 167147 31327 167175
rect 31361 167147 31389 167175
rect 31299 167085 31327 167113
rect 31361 167085 31389 167113
rect 31299 167023 31327 167051
rect 31361 167023 31389 167051
rect 31299 166961 31327 166989
rect 31361 166961 31389 166989
rect 23619 164147 23647 164175
rect 23681 164147 23709 164175
rect 23619 164085 23647 164113
rect 23681 164085 23709 164113
rect 23619 164023 23647 164051
rect 23681 164023 23709 164051
rect 23619 163961 23647 163989
rect 23681 163961 23709 163989
rect 33477 164147 33505 164175
rect 33539 164147 33567 164175
rect 33601 164147 33629 164175
rect 33663 164147 33691 164175
rect 33477 164085 33505 164113
rect 33539 164085 33567 164113
rect 33601 164085 33629 164113
rect 33663 164085 33691 164113
rect 33477 164023 33505 164051
rect 33539 164023 33567 164051
rect 33601 164023 33629 164051
rect 33663 164023 33691 164051
rect 33477 163961 33505 163989
rect 33539 163961 33567 163989
rect 33601 163961 33629 163989
rect 33663 163961 33691 163989
rect 19977 158147 20005 158175
rect 20039 158147 20067 158175
rect 20101 158147 20129 158175
rect 20163 158147 20191 158175
rect 19977 158085 20005 158113
rect 20039 158085 20067 158113
rect 20101 158085 20129 158113
rect 20163 158085 20191 158113
rect 19977 158023 20005 158051
rect 20039 158023 20067 158051
rect 20101 158023 20129 158051
rect 20163 158023 20191 158051
rect 19977 157961 20005 157989
rect 20039 157961 20067 157989
rect 20101 157961 20129 157989
rect 20163 157961 20191 157989
rect 31299 158147 31327 158175
rect 31361 158147 31389 158175
rect 31299 158085 31327 158113
rect 31361 158085 31389 158113
rect 31299 158023 31327 158051
rect 31361 158023 31389 158051
rect 31299 157961 31327 157989
rect 31361 157961 31389 157989
rect 23619 155147 23647 155175
rect 23681 155147 23709 155175
rect 23619 155085 23647 155113
rect 23681 155085 23709 155113
rect 23619 155023 23647 155051
rect 23681 155023 23709 155051
rect 23619 154961 23647 154989
rect 23681 154961 23709 154989
rect 33477 155147 33505 155175
rect 33539 155147 33567 155175
rect 33601 155147 33629 155175
rect 33663 155147 33691 155175
rect 33477 155085 33505 155113
rect 33539 155085 33567 155113
rect 33601 155085 33629 155113
rect 33663 155085 33691 155113
rect 33477 155023 33505 155051
rect 33539 155023 33567 155051
rect 33601 155023 33629 155051
rect 33663 155023 33691 155051
rect 33477 154961 33505 154989
rect 33539 154961 33567 154989
rect 33601 154961 33629 154989
rect 33663 154961 33691 154989
rect 19977 149147 20005 149175
rect 20039 149147 20067 149175
rect 20101 149147 20129 149175
rect 20163 149147 20191 149175
rect 19977 149085 20005 149113
rect 20039 149085 20067 149113
rect 20101 149085 20129 149113
rect 20163 149085 20191 149113
rect 19977 149023 20005 149051
rect 20039 149023 20067 149051
rect 20101 149023 20129 149051
rect 20163 149023 20191 149051
rect 19977 148961 20005 148989
rect 20039 148961 20067 148989
rect 20101 148961 20129 148989
rect 20163 148961 20191 148989
rect 31299 149147 31327 149175
rect 31361 149147 31389 149175
rect 31299 149085 31327 149113
rect 31361 149085 31389 149113
rect 31299 149023 31327 149051
rect 31361 149023 31389 149051
rect 31299 148961 31327 148989
rect 31361 148961 31389 148989
rect 23619 146147 23647 146175
rect 23681 146147 23709 146175
rect 23619 146085 23647 146113
rect 23681 146085 23709 146113
rect 23619 146023 23647 146051
rect 23681 146023 23709 146051
rect 23619 145961 23647 145989
rect 23681 145961 23709 145989
rect 33477 146147 33505 146175
rect 33539 146147 33567 146175
rect 33601 146147 33629 146175
rect 33663 146147 33691 146175
rect 33477 146085 33505 146113
rect 33539 146085 33567 146113
rect 33601 146085 33629 146113
rect 33663 146085 33691 146113
rect 33477 146023 33505 146051
rect 33539 146023 33567 146051
rect 33601 146023 33629 146051
rect 33663 146023 33691 146051
rect 33477 145961 33505 145989
rect 33539 145961 33567 145989
rect 33601 145961 33629 145989
rect 33663 145961 33691 145989
rect 19977 140147 20005 140175
rect 20039 140147 20067 140175
rect 20101 140147 20129 140175
rect 20163 140147 20191 140175
rect 19977 140085 20005 140113
rect 20039 140085 20067 140113
rect 20101 140085 20129 140113
rect 20163 140085 20191 140113
rect 19977 140023 20005 140051
rect 20039 140023 20067 140051
rect 20101 140023 20129 140051
rect 20163 140023 20191 140051
rect 19977 139961 20005 139989
rect 20039 139961 20067 139989
rect 20101 139961 20129 139989
rect 20163 139961 20191 139989
rect 31299 140147 31327 140175
rect 31361 140147 31389 140175
rect 31299 140085 31327 140113
rect 31361 140085 31389 140113
rect 31299 140023 31327 140051
rect 31361 140023 31389 140051
rect 31299 139961 31327 139989
rect 31361 139961 31389 139989
rect 23619 137147 23647 137175
rect 23681 137147 23709 137175
rect 23619 137085 23647 137113
rect 23681 137085 23709 137113
rect 23619 137023 23647 137051
rect 23681 137023 23709 137051
rect 23619 136961 23647 136989
rect 23681 136961 23709 136989
rect 33477 137147 33505 137175
rect 33539 137147 33567 137175
rect 33601 137147 33629 137175
rect 33663 137147 33691 137175
rect 33477 137085 33505 137113
rect 33539 137085 33567 137113
rect 33601 137085 33629 137113
rect 33663 137085 33691 137113
rect 33477 137023 33505 137051
rect 33539 137023 33567 137051
rect 33601 137023 33629 137051
rect 33663 137023 33691 137051
rect 33477 136961 33505 136989
rect 33539 136961 33567 136989
rect 33601 136961 33629 136989
rect 33663 136961 33691 136989
rect 19977 131147 20005 131175
rect 20039 131147 20067 131175
rect 20101 131147 20129 131175
rect 20163 131147 20191 131175
rect 19977 131085 20005 131113
rect 20039 131085 20067 131113
rect 20101 131085 20129 131113
rect 20163 131085 20191 131113
rect 19977 131023 20005 131051
rect 20039 131023 20067 131051
rect 20101 131023 20129 131051
rect 20163 131023 20191 131051
rect 19977 130961 20005 130989
rect 20039 130961 20067 130989
rect 20101 130961 20129 130989
rect 20163 130961 20191 130989
rect 31299 131147 31327 131175
rect 31361 131147 31389 131175
rect 31299 131085 31327 131113
rect 31361 131085 31389 131113
rect 31299 131023 31327 131051
rect 31361 131023 31389 131051
rect 31299 130961 31327 130989
rect 31361 130961 31389 130989
rect 23619 128147 23647 128175
rect 23681 128147 23709 128175
rect 23619 128085 23647 128113
rect 23681 128085 23709 128113
rect 23619 128023 23647 128051
rect 23681 128023 23709 128051
rect 23619 127961 23647 127989
rect 23681 127961 23709 127989
rect 33477 128147 33505 128175
rect 33539 128147 33567 128175
rect 33601 128147 33629 128175
rect 33663 128147 33691 128175
rect 33477 128085 33505 128113
rect 33539 128085 33567 128113
rect 33601 128085 33629 128113
rect 33663 128085 33691 128113
rect 33477 128023 33505 128051
rect 33539 128023 33567 128051
rect 33601 128023 33629 128051
rect 33663 128023 33691 128051
rect 33477 127961 33505 127989
rect 33539 127961 33567 127989
rect 33601 127961 33629 127989
rect 33663 127961 33691 127989
rect 19977 122147 20005 122175
rect 20039 122147 20067 122175
rect 20101 122147 20129 122175
rect 20163 122147 20191 122175
rect 19977 122085 20005 122113
rect 20039 122085 20067 122113
rect 20101 122085 20129 122113
rect 20163 122085 20191 122113
rect 19977 122023 20005 122051
rect 20039 122023 20067 122051
rect 20101 122023 20129 122051
rect 20163 122023 20191 122051
rect 19977 121961 20005 121989
rect 20039 121961 20067 121989
rect 20101 121961 20129 121989
rect 20163 121961 20191 121989
rect 31299 122147 31327 122175
rect 31361 122147 31389 122175
rect 31299 122085 31327 122113
rect 31361 122085 31389 122113
rect 31299 122023 31327 122051
rect 31361 122023 31389 122051
rect 31299 121961 31327 121989
rect 31361 121961 31389 121989
rect 23619 119147 23647 119175
rect 23681 119147 23709 119175
rect 23619 119085 23647 119113
rect 23681 119085 23709 119113
rect 23619 119023 23647 119051
rect 23681 119023 23709 119051
rect 23619 118961 23647 118989
rect 23681 118961 23709 118989
rect 33477 119147 33505 119175
rect 33539 119147 33567 119175
rect 33601 119147 33629 119175
rect 33663 119147 33691 119175
rect 33477 119085 33505 119113
rect 33539 119085 33567 119113
rect 33601 119085 33629 119113
rect 33663 119085 33691 119113
rect 33477 119023 33505 119051
rect 33539 119023 33567 119051
rect 33601 119023 33629 119051
rect 33663 119023 33691 119051
rect 33477 118961 33505 118989
rect 33539 118961 33567 118989
rect 33601 118961 33629 118989
rect 33663 118961 33691 118989
rect 19977 113147 20005 113175
rect 20039 113147 20067 113175
rect 20101 113147 20129 113175
rect 20163 113147 20191 113175
rect 19977 113085 20005 113113
rect 20039 113085 20067 113113
rect 20101 113085 20129 113113
rect 20163 113085 20191 113113
rect 19977 113023 20005 113051
rect 20039 113023 20067 113051
rect 20101 113023 20129 113051
rect 20163 113023 20191 113051
rect 19977 112961 20005 112989
rect 20039 112961 20067 112989
rect 20101 112961 20129 112989
rect 20163 112961 20191 112989
rect 31299 113147 31327 113175
rect 31361 113147 31389 113175
rect 31299 113085 31327 113113
rect 31361 113085 31389 113113
rect 31299 113023 31327 113051
rect 31361 113023 31389 113051
rect 31299 112961 31327 112989
rect 31361 112961 31389 112989
rect 23619 110147 23647 110175
rect 23681 110147 23709 110175
rect 23619 110085 23647 110113
rect 23681 110085 23709 110113
rect 23619 110023 23647 110051
rect 23681 110023 23709 110051
rect 23619 109961 23647 109989
rect 23681 109961 23709 109989
rect 33477 110147 33505 110175
rect 33539 110147 33567 110175
rect 33601 110147 33629 110175
rect 33663 110147 33691 110175
rect 33477 110085 33505 110113
rect 33539 110085 33567 110113
rect 33601 110085 33629 110113
rect 33663 110085 33691 110113
rect 33477 110023 33505 110051
rect 33539 110023 33567 110051
rect 33601 110023 33629 110051
rect 33663 110023 33691 110051
rect 33477 109961 33505 109989
rect 33539 109961 33567 109989
rect 33601 109961 33629 109989
rect 33663 109961 33691 109989
rect 19977 104147 20005 104175
rect 20039 104147 20067 104175
rect 20101 104147 20129 104175
rect 20163 104147 20191 104175
rect 19977 104085 20005 104113
rect 20039 104085 20067 104113
rect 20101 104085 20129 104113
rect 20163 104085 20191 104113
rect 19977 104023 20005 104051
rect 20039 104023 20067 104051
rect 20101 104023 20129 104051
rect 20163 104023 20191 104051
rect 19977 103961 20005 103989
rect 20039 103961 20067 103989
rect 20101 103961 20129 103989
rect 20163 103961 20191 103989
rect 31299 104147 31327 104175
rect 31361 104147 31389 104175
rect 31299 104085 31327 104113
rect 31361 104085 31389 104113
rect 31299 104023 31327 104051
rect 31361 104023 31389 104051
rect 31299 103961 31327 103989
rect 31361 103961 31389 103989
rect 23619 101147 23647 101175
rect 23681 101147 23709 101175
rect 23619 101085 23647 101113
rect 23681 101085 23709 101113
rect 23619 101023 23647 101051
rect 23681 101023 23709 101051
rect 23619 100961 23647 100989
rect 23681 100961 23709 100989
rect 33477 101147 33505 101175
rect 33539 101147 33567 101175
rect 33601 101147 33629 101175
rect 33663 101147 33691 101175
rect 33477 101085 33505 101113
rect 33539 101085 33567 101113
rect 33601 101085 33629 101113
rect 33663 101085 33691 101113
rect 33477 101023 33505 101051
rect 33539 101023 33567 101051
rect 33601 101023 33629 101051
rect 33663 101023 33691 101051
rect 33477 100961 33505 100989
rect 33539 100961 33567 100989
rect 33601 100961 33629 100989
rect 33663 100961 33691 100989
rect 19977 95147 20005 95175
rect 20039 95147 20067 95175
rect 20101 95147 20129 95175
rect 20163 95147 20191 95175
rect 19977 95085 20005 95113
rect 20039 95085 20067 95113
rect 20101 95085 20129 95113
rect 20163 95085 20191 95113
rect 19977 95023 20005 95051
rect 20039 95023 20067 95051
rect 20101 95023 20129 95051
rect 20163 95023 20191 95051
rect 19977 94961 20005 94989
rect 20039 94961 20067 94989
rect 20101 94961 20129 94989
rect 20163 94961 20191 94989
rect 31299 95147 31327 95175
rect 31361 95147 31389 95175
rect 31299 95085 31327 95113
rect 31361 95085 31389 95113
rect 31299 95023 31327 95051
rect 31361 95023 31389 95051
rect 31299 94961 31327 94989
rect 31361 94961 31389 94989
rect 23619 92147 23647 92175
rect 23681 92147 23709 92175
rect 23619 92085 23647 92113
rect 23681 92085 23709 92113
rect 23619 92023 23647 92051
rect 23681 92023 23709 92051
rect 23619 91961 23647 91989
rect 23681 91961 23709 91989
rect 33477 92147 33505 92175
rect 33539 92147 33567 92175
rect 33601 92147 33629 92175
rect 33663 92147 33691 92175
rect 33477 92085 33505 92113
rect 33539 92085 33567 92113
rect 33601 92085 33629 92113
rect 33663 92085 33691 92113
rect 33477 92023 33505 92051
rect 33539 92023 33567 92051
rect 33601 92023 33629 92051
rect 33663 92023 33691 92051
rect 33477 91961 33505 91989
rect 33539 91961 33567 91989
rect 33601 91961 33629 91989
rect 33663 91961 33691 91989
rect 19977 86147 20005 86175
rect 20039 86147 20067 86175
rect 20101 86147 20129 86175
rect 20163 86147 20191 86175
rect 19977 86085 20005 86113
rect 20039 86085 20067 86113
rect 20101 86085 20129 86113
rect 20163 86085 20191 86113
rect 19977 86023 20005 86051
rect 20039 86023 20067 86051
rect 20101 86023 20129 86051
rect 20163 86023 20191 86051
rect 19977 85961 20005 85989
rect 20039 85961 20067 85989
rect 20101 85961 20129 85989
rect 20163 85961 20191 85989
rect 31299 86147 31327 86175
rect 31361 86147 31389 86175
rect 31299 86085 31327 86113
rect 31361 86085 31389 86113
rect 31299 86023 31327 86051
rect 31361 86023 31389 86051
rect 31299 85961 31327 85989
rect 31361 85961 31389 85989
rect 23619 83147 23647 83175
rect 23681 83147 23709 83175
rect 23619 83085 23647 83113
rect 23681 83085 23709 83113
rect 23619 83023 23647 83051
rect 23681 83023 23709 83051
rect 23619 82961 23647 82989
rect 23681 82961 23709 82989
rect 33477 83147 33505 83175
rect 33539 83147 33567 83175
rect 33601 83147 33629 83175
rect 33663 83147 33691 83175
rect 33477 83085 33505 83113
rect 33539 83085 33567 83113
rect 33601 83085 33629 83113
rect 33663 83085 33691 83113
rect 33477 83023 33505 83051
rect 33539 83023 33567 83051
rect 33601 83023 33629 83051
rect 33663 83023 33691 83051
rect 33477 82961 33505 82989
rect 33539 82961 33567 82989
rect 33601 82961 33629 82989
rect 33663 82961 33691 82989
rect 19977 77147 20005 77175
rect 20039 77147 20067 77175
rect 20101 77147 20129 77175
rect 20163 77147 20191 77175
rect 19977 77085 20005 77113
rect 20039 77085 20067 77113
rect 20101 77085 20129 77113
rect 20163 77085 20191 77113
rect 19977 77023 20005 77051
rect 20039 77023 20067 77051
rect 20101 77023 20129 77051
rect 20163 77023 20191 77051
rect 19977 76961 20005 76989
rect 20039 76961 20067 76989
rect 20101 76961 20129 76989
rect 20163 76961 20191 76989
rect 31299 77147 31327 77175
rect 31361 77147 31389 77175
rect 31299 77085 31327 77113
rect 31361 77085 31389 77113
rect 31299 77023 31327 77051
rect 31361 77023 31389 77051
rect 31299 76961 31327 76989
rect 31361 76961 31389 76989
rect 23619 74147 23647 74175
rect 23681 74147 23709 74175
rect 23619 74085 23647 74113
rect 23681 74085 23709 74113
rect 23619 74023 23647 74051
rect 23681 74023 23709 74051
rect 23619 73961 23647 73989
rect 23681 73961 23709 73989
rect 33477 74147 33505 74175
rect 33539 74147 33567 74175
rect 33601 74147 33629 74175
rect 33663 74147 33691 74175
rect 33477 74085 33505 74113
rect 33539 74085 33567 74113
rect 33601 74085 33629 74113
rect 33663 74085 33691 74113
rect 33477 74023 33505 74051
rect 33539 74023 33567 74051
rect 33601 74023 33629 74051
rect 33663 74023 33691 74051
rect 33477 73961 33505 73989
rect 33539 73961 33567 73989
rect 33601 73961 33629 73989
rect 33663 73961 33691 73989
rect 19977 68147 20005 68175
rect 20039 68147 20067 68175
rect 20101 68147 20129 68175
rect 20163 68147 20191 68175
rect 19977 68085 20005 68113
rect 20039 68085 20067 68113
rect 20101 68085 20129 68113
rect 20163 68085 20191 68113
rect 19977 68023 20005 68051
rect 20039 68023 20067 68051
rect 20101 68023 20129 68051
rect 20163 68023 20191 68051
rect 19977 67961 20005 67989
rect 20039 67961 20067 67989
rect 20101 67961 20129 67989
rect 20163 67961 20191 67989
rect 31299 68147 31327 68175
rect 31361 68147 31389 68175
rect 31299 68085 31327 68113
rect 31361 68085 31389 68113
rect 31299 68023 31327 68051
rect 31361 68023 31389 68051
rect 31299 67961 31327 67989
rect 31361 67961 31389 67989
rect 23619 65147 23647 65175
rect 23681 65147 23709 65175
rect 23619 65085 23647 65113
rect 23681 65085 23709 65113
rect 23619 65023 23647 65051
rect 23681 65023 23709 65051
rect 23619 64961 23647 64989
rect 23681 64961 23709 64989
rect 33477 65147 33505 65175
rect 33539 65147 33567 65175
rect 33601 65147 33629 65175
rect 33663 65147 33691 65175
rect 33477 65085 33505 65113
rect 33539 65085 33567 65113
rect 33601 65085 33629 65113
rect 33663 65085 33691 65113
rect 33477 65023 33505 65051
rect 33539 65023 33567 65051
rect 33601 65023 33629 65051
rect 33663 65023 33691 65051
rect 33477 64961 33505 64989
rect 33539 64961 33567 64989
rect 33601 64961 33629 64989
rect 33663 64961 33691 64989
rect 19977 59147 20005 59175
rect 20039 59147 20067 59175
rect 20101 59147 20129 59175
rect 20163 59147 20191 59175
rect 19977 59085 20005 59113
rect 20039 59085 20067 59113
rect 20101 59085 20129 59113
rect 20163 59085 20191 59113
rect 19977 59023 20005 59051
rect 20039 59023 20067 59051
rect 20101 59023 20129 59051
rect 20163 59023 20191 59051
rect 19977 58961 20005 58989
rect 20039 58961 20067 58989
rect 20101 58961 20129 58989
rect 20163 58961 20191 58989
rect 31299 59147 31327 59175
rect 31361 59147 31389 59175
rect 31299 59085 31327 59113
rect 31361 59085 31389 59113
rect 31299 59023 31327 59051
rect 31361 59023 31389 59051
rect 31299 58961 31327 58989
rect 31361 58961 31389 58989
rect 23619 56147 23647 56175
rect 23681 56147 23709 56175
rect 23619 56085 23647 56113
rect 23681 56085 23709 56113
rect 23619 56023 23647 56051
rect 23681 56023 23709 56051
rect 23619 55961 23647 55989
rect 23681 55961 23709 55989
rect 33477 56147 33505 56175
rect 33539 56147 33567 56175
rect 33601 56147 33629 56175
rect 33663 56147 33691 56175
rect 33477 56085 33505 56113
rect 33539 56085 33567 56113
rect 33601 56085 33629 56113
rect 33663 56085 33691 56113
rect 33477 56023 33505 56051
rect 33539 56023 33567 56051
rect 33601 56023 33629 56051
rect 33663 56023 33691 56051
rect 33477 55961 33505 55989
rect 33539 55961 33567 55989
rect 33601 55961 33629 55989
rect 33663 55961 33691 55989
rect 19977 50147 20005 50175
rect 20039 50147 20067 50175
rect 20101 50147 20129 50175
rect 20163 50147 20191 50175
rect 19977 50085 20005 50113
rect 20039 50085 20067 50113
rect 20101 50085 20129 50113
rect 20163 50085 20191 50113
rect 19977 50023 20005 50051
rect 20039 50023 20067 50051
rect 20101 50023 20129 50051
rect 20163 50023 20191 50051
rect 19977 49961 20005 49989
rect 20039 49961 20067 49989
rect 20101 49961 20129 49989
rect 20163 49961 20191 49989
rect 31299 50147 31327 50175
rect 31361 50147 31389 50175
rect 31299 50085 31327 50113
rect 31361 50085 31389 50113
rect 31299 50023 31327 50051
rect 31361 50023 31389 50051
rect 31299 49961 31327 49989
rect 31361 49961 31389 49989
rect 23619 47147 23647 47175
rect 23681 47147 23709 47175
rect 23619 47085 23647 47113
rect 23681 47085 23709 47113
rect 23619 47023 23647 47051
rect 23681 47023 23709 47051
rect 23619 46961 23647 46989
rect 23681 46961 23709 46989
rect 33477 47147 33505 47175
rect 33539 47147 33567 47175
rect 33601 47147 33629 47175
rect 33663 47147 33691 47175
rect 33477 47085 33505 47113
rect 33539 47085 33567 47113
rect 33601 47085 33629 47113
rect 33663 47085 33691 47113
rect 33477 47023 33505 47051
rect 33539 47023 33567 47051
rect 33601 47023 33629 47051
rect 33663 47023 33691 47051
rect 33477 46961 33505 46989
rect 33539 46961 33567 46989
rect 33601 46961 33629 46989
rect 33663 46961 33691 46989
rect 19977 41147 20005 41175
rect 20039 41147 20067 41175
rect 20101 41147 20129 41175
rect 20163 41147 20191 41175
rect 19977 41085 20005 41113
rect 20039 41085 20067 41113
rect 20101 41085 20129 41113
rect 20163 41085 20191 41113
rect 19977 41023 20005 41051
rect 20039 41023 20067 41051
rect 20101 41023 20129 41051
rect 20163 41023 20191 41051
rect 19977 40961 20005 40989
rect 20039 40961 20067 40989
rect 20101 40961 20129 40989
rect 20163 40961 20191 40989
rect 31299 41147 31327 41175
rect 31361 41147 31389 41175
rect 31299 41085 31327 41113
rect 31361 41085 31389 41113
rect 31299 41023 31327 41051
rect 31361 41023 31389 41051
rect 31299 40961 31327 40989
rect 31361 40961 31389 40989
rect 23619 38147 23647 38175
rect 23681 38147 23709 38175
rect 23619 38085 23647 38113
rect 23681 38085 23709 38113
rect 23619 38023 23647 38051
rect 23681 38023 23709 38051
rect 23619 37961 23647 37989
rect 23681 37961 23709 37989
rect 33477 38147 33505 38175
rect 33539 38147 33567 38175
rect 33601 38147 33629 38175
rect 33663 38147 33691 38175
rect 33477 38085 33505 38113
rect 33539 38085 33567 38113
rect 33601 38085 33629 38113
rect 33663 38085 33691 38113
rect 33477 38023 33505 38051
rect 33539 38023 33567 38051
rect 33601 38023 33629 38051
rect 33663 38023 33691 38051
rect 33477 37961 33505 37989
rect 33539 37961 33567 37989
rect 33601 37961 33629 37989
rect 33663 37961 33691 37989
rect 19977 32147 20005 32175
rect 20039 32147 20067 32175
rect 20101 32147 20129 32175
rect 20163 32147 20191 32175
rect 19977 32085 20005 32113
rect 20039 32085 20067 32113
rect 20101 32085 20129 32113
rect 20163 32085 20191 32113
rect 19977 32023 20005 32051
rect 20039 32023 20067 32051
rect 20101 32023 20129 32051
rect 20163 32023 20191 32051
rect 19977 31961 20005 31989
rect 20039 31961 20067 31989
rect 20101 31961 20129 31989
rect 20163 31961 20191 31989
rect 31299 32147 31327 32175
rect 31361 32147 31389 32175
rect 31299 32085 31327 32113
rect 31361 32085 31389 32113
rect 31299 32023 31327 32051
rect 31361 32023 31389 32051
rect 31299 31961 31327 31989
rect 31361 31961 31389 31989
rect 23619 29147 23647 29175
rect 23681 29147 23709 29175
rect 23619 29085 23647 29113
rect 23681 29085 23709 29113
rect 23619 29023 23647 29051
rect 23681 29023 23709 29051
rect 23619 28961 23647 28989
rect 23681 28961 23709 28989
rect 33477 29147 33505 29175
rect 33539 29147 33567 29175
rect 33601 29147 33629 29175
rect 33663 29147 33691 29175
rect 33477 29085 33505 29113
rect 33539 29085 33567 29113
rect 33601 29085 33629 29113
rect 33663 29085 33691 29113
rect 33477 29023 33505 29051
rect 33539 29023 33567 29051
rect 33601 29023 33629 29051
rect 33663 29023 33691 29051
rect 33477 28961 33505 28989
rect 33539 28961 33567 28989
rect 33601 28961 33629 28989
rect 33663 28961 33691 28989
rect 19977 23147 20005 23175
rect 20039 23147 20067 23175
rect 20101 23147 20129 23175
rect 20163 23147 20191 23175
rect 19977 23085 20005 23113
rect 20039 23085 20067 23113
rect 20101 23085 20129 23113
rect 20163 23085 20191 23113
rect 19977 23023 20005 23051
rect 20039 23023 20067 23051
rect 20101 23023 20129 23051
rect 20163 23023 20191 23051
rect 19977 22961 20005 22989
rect 20039 22961 20067 22989
rect 20101 22961 20129 22989
rect 20163 22961 20191 22989
rect 31299 23147 31327 23175
rect 31361 23147 31389 23175
rect 31299 23085 31327 23113
rect 31361 23085 31389 23113
rect 31299 23023 31327 23051
rect 31361 23023 31389 23051
rect 31299 22961 31327 22989
rect 31361 22961 31389 22989
rect 23619 20147 23647 20175
rect 23681 20147 23709 20175
rect 23619 20085 23647 20113
rect 23681 20085 23709 20113
rect 23619 20023 23647 20051
rect 23681 20023 23709 20051
rect 23619 19961 23647 19989
rect 23681 19961 23709 19989
rect 33477 20147 33505 20175
rect 33539 20147 33567 20175
rect 33601 20147 33629 20175
rect 33663 20147 33691 20175
rect 33477 20085 33505 20113
rect 33539 20085 33567 20113
rect 33601 20085 33629 20113
rect 33663 20085 33691 20113
rect 33477 20023 33505 20051
rect 33539 20023 33567 20051
rect 33601 20023 33629 20051
rect 33663 20023 33691 20051
rect 33477 19961 33505 19989
rect 33539 19961 33567 19989
rect 33601 19961 33629 19989
rect 33663 19961 33691 19989
rect 19977 14147 20005 14175
rect 20039 14147 20067 14175
rect 20101 14147 20129 14175
rect 20163 14147 20191 14175
rect 19977 14085 20005 14113
rect 20039 14085 20067 14113
rect 20101 14085 20129 14113
rect 20163 14085 20191 14113
rect 19977 14023 20005 14051
rect 20039 14023 20067 14051
rect 20101 14023 20129 14051
rect 20163 14023 20191 14051
rect 19977 13961 20005 13989
rect 20039 13961 20067 13989
rect 20101 13961 20129 13989
rect 20163 13961 20191 13989
rect 31299 14147 31327 14175
rect 31361 14147 31389 14175
rect 31299 14085 31327 14113
rect 31361 14085 31389 14113
rect 31299 14023 31327 14051
rect 31361 14023 31389 14051
rect 31299 13961 31327 13989
rect 31361 13961 31389 13989
rect 23619 11147 23647 11175
rect 23681 11147 23709 11175
rect 23619 11085 23647 11113
rect 23681 11085 23709 11113
rect 23619 11023 23647 11051
rect 23681 11023 23709 11051
rect 23619 10961 23647 10989
rect 23681 10961 23709 10989
rect 33477 11147 33505 11175
rect 33539 11147 33567 11175
rect 33601 11147 33629 11175
rect 33663 11147 33691 11175
rect 33477 11085 33505 11113
rect 33539 11085 33567 11113
rect 33601 11085 33629 11113
rect 33663 11085 33691 11113
rect 33477 11023 33505 11051
rect 33539 11023 33567 11051
rect 33601 11023 33629 11051
rect 33663 11023 33691 11051
rect 33477 10961 33505 10989
rect 33539 10961 33567 10989
rect 33601 10961 33629 10989
rect 33663 10961 33691 10989
rect 19977 5147 20005 5175
rect 20039 5147 20067 5175
rect 20101 5147 20129 5175
rect 20163 5147 20191 5175
rect 19977 5085 20005 5113
rect 20039 5085 20067 5113
rect 20101 5085 20129 5113
rect 20163 5085 20191 5113
rect 19977 5023 20005 5051
rect 20039 5023 20067 5051
rect 20101 5023 20129 5051
rect 20163 5023 20191 5051
rect 19977 4961 20005 4989
rect 20039 4961 20067 4989
rect 20101 4961 20129 4989
rect 20163 4961 20191 4989
rect 31299 5147 31327 5175
rect 31361 5147 31389 5175
rect 31299 5085 31327 5113
rect 31361 5085 31389 5113
rect 31299 5023 31327 5051
rect 31361 5023 31389 5051
rect 31299 4961 31327 4989
rect 31361 4961 31389 4989
rect 19977 -588 20005 -560
rect 20039 -588 20067 -560
rect 20101 -588 20129 -560
rect 20163 -588 20191 -560
rect 19977 -650 20005 -622
rect 20039 -650 20067 -622
rect 20101 -650 20129 -622
rect 20163 -650 20191 -622
rect 19977 -712 20005 -684
rect 20039 -712 20067 -684
rect 20101 -712 20129 -684
rect 20163 -712 20191 -684
rect 19977 -774 20005 -746
rect 20039 -774 20067 -746
rect 20101 -774 20129 -746
rect 20163 -774 20191 -746
rect 33477 2147 33505 2175
rect 33539 2147 33567 2175
rect 33601 2147 33629 2175
rect 33663 2147 33691 2175
rect 33477 2085 33505 2113
rect 33539 2085 33567 2113
rect 33601 2085 33629 2113
rect 33663 2085 33691 2113
rect 33477 2023 33505 2051
rect 33539 2023 33567 2051
rect 33601 2023 33629 2051
rect 33663 2023 33691 2051
rect 33477 1961 33505 1989
rect 33539 1961 33567 1989
rect 33601 1961 33629 1989
rect 33663 1961 33691 1989
rect 33477 -108 33505 -80
rect 33539 -108 33567 -80
rect 33601 -108 33629 -80
rect 33663 -108 33691 -80
rect 33477 -170 33505 -142
rect 33539 -170 33567 -142
rect 33601 -170 33629 -142
rect 33663 -170 33691 -142
rect 33477 -232 33505 -204
rect 33539 -232 33567 -204
rect 33601 -232 33629 -204
rect 33663 -232 33691 -204
rect 33477 -294 33505 -266
rect 33539 -294 33567 -266
rect 33601 -294 33629 -266
rect 33663 -294 33691 -266
rect 35337 299058 35365 299086
rect 35399 299058 35427 299086
rect 35461 299058 35489 299086
rect 35523 299058 35551 299086
rect 35337 298996 35365 299024
rect 35399 298996 35427 299024
rect 35461 298996 35489 299024
rect 35523 298996 35551 299024
rect 35337 298934 35365 298962
rect 35399 298934 35427 298962
rect 35461 298934 35489 298962
rect 35523 298934 35551 298962
rect 35337 298872 35365 298900
rect 35399 298872 35427 298900
rect 35461 298872 35489 298900
rect 35523 298872 35551 298900
rect 35337 293147 35365 293175
rect 35399 293147 35427 293175
rect 35461 293147 35489 293175
rect 35523 293147 35551 293175
rect 35337 293085 35365 293113
rect 35399 293085 35427 293113
rect 35461 293085 35489 293113
rect 35523 293085 35551 293113
rect 35337 293023 35365 293051
rect 35399 293023 35427 293051
rect 35461 293023 35489 293051
rect 35523 293023 35551 293051
rect 35337 292961 35365 292989
rect 35399 292961 35427 292989
rect 35461 292961 35489 292989
rect 35523 292961 35551 292989
rect 35337 284147 35365 284175
rect 35399 284147 35427 284175
rect 35461 284147 35489 284175
rect 35523 284147 35551 284175
rect 35337 284085 35365 284113
rect 35399 284085 35427 284113
rect 35461 284085 35489 284113
rect 35523 284085 35551 284113
rect 35337 284023 35365 284051
rect 35399 284023 35427 284051
rect 35461 284023 35489 284051
rect 35523 284023 35551 284051
rect 35337 283961 35365 283989
rect 35399 283961 35427 283989
rect 35461 283961 35489 283989
rect 35523 283961 35551 283989
rect 35337 275147 35365 275175
rect 35399 275147 35427 275175
rect 35461 275147 35489 275175
rect 35523 275147 35551 275175
rect 35337 275085 35365 275113
rect 35399 275085 35427 275113
rect 35461 275085 35489 275113
rect 35523 275085 35551 275113
rect 35337 275023 35365 275051
rect 35399 275023 35427 275051
rect 35461 275023 35489 275051
rect 35523 275023 35551 275051
rect 35337 274961 35365 274989
rect 35399 274961 35427 274989
rect 35461 274961 35489 274989
rect 35523 274961 35551 274989
rect 35337 266147 35365 266175
rect 35399 266147 35427 266175
rect 35461 266147 35489 266175
rect 35523 266147 35551 266175
rect 35337 266085 35365 266113
rect 35399 266085 35427 266113
rect 35461 266085 35489 266113
rect 35523 266085 35551 266113
rect 35337 266023 35365 266051
rect 35399 266023 35427 266051
rect 35461 266023 35489 266051
rect 35523 266023 35551 266051
rect 35337 265961 35365 265989
rect 35399 265961 35427 265989
rect 35461 265961 35489 265989
rect 35523 265961 35551 265989
rect 35337 257147 35365 257175
rect 35399 257147 35427 257175
rect 35461 257147 35489 257175
rect 35523 257147 35551 257175
rect 35337 257085 35365 257113
rect 35399 257085 35427 257113
rect 35461 257085 35489 257113
rect 35523 257085 35551 257113
rect 35337 257023 35365 257051
rect 35399 257023 35427 257051
rect 35461 257023 35489 257051
rect 35523 257023 35551 257051
rect 35337 256961 35365 256989
rect 35399 256961 35427 256989
rect 35461 256961 35489 256989
rect 35523 256961 35551 256989
rect 35337 248147 35365 248175
rect 35399 248147 35427 248175
rect 35461 248147 35489 248175
rect 35523 248147 35551 248175
rect 35337 248085 35365 248113
rect 35399 248085 35427 248113
rect 35461 248085 35489 248113
rect 35523 248085 35551 248113
rect 35337 248023 35365 248051
rect 35399 248023 35427 248051
rect 35461 248023 35489 248051
rect 35523 248023 35551 248051
rect 35337 247961 35365 247989
rect 35399 247961 35427 247989
rect 35461 247961 35489 247989
rect 35523 247961 35551 247989
rect 35337 239147 35365 239175
rect 35399 239147 35427 239175
rect 35461 239147 35489 239175
rect 35523 239147 35551 239175
rect 35337 239085 35365 239113
rect 35399 239085 35427 239113
rect 35461 239085 35489 239113
rect 35523 239085 35551 239113
rect 35337 239023 35365 239051
rect 35399 239023 35427 239051
rect 35461 239023 35489 239051
rect 35523 239023 35551 239051
rect 35337 238961 35365 238989
rect 35399 238961 35427 238989
rect 35461 238961 35489 238989
rect 35523 238961 35551 238989
rect 35337 230147 35365 230175
rect 35399 230147 35427 230175
rect 35461 230147 35489 230175
rect 35523 230147 35551 230175
rect 35337 230085 35365 230113
rect 35399 230085 35427 230113
rect 35461 230085 35489 230113
rect 35523 230085 35551 230113
rect 35337 230023 35365 230051
rect 35399 230023 35427 230051
rect 35461 230023 35489 230051
rect 35523 230023 35551 230051
rect 35337 229961 35365 229989
rect 35399 229961 35427 229989
rect 35461 229961 35489 229989
rect 35523 229961 35551 229989
rect 35337 221147 35365 221175
rect 35399 221147 35427 221175
rect 35461 221147 35489 221175
rect 35523 221147 35551 221175
rect 35337 221085 35365 221113
rect 35399 221085 35427 221113
rect 35461 221085 35489 221113
rect 35523 221085 35551 221113
rect 35337 221023 35365 221051
rect 35399 221023 35427 221051
rect 35461 221023 35489 221051
rect 35523 221023 35551 221051
rect 35337 220961 35365 220989
rect 35399 220961 35427 220989
rect 35461 220961 35489 220989
rect 35523 220961 35551 220989
rect 35337 212147 35365 212175
rect 35399 212147 35427 212175
rect 35461 212147 35489 212175
rect 35523 212147 35551 212175
rect 35337 212085 35365 212113
rect 35399 212085 35427 212113
rect 35461 212085 35489 212113
rect 35523 212085 35551 212113
rect 35337 212023 35365 212051
rect 35399 212023 35427 212051
rect 35461 212023 35489 212051
rect 35523 212023 35551 212051
rect 35337 211961 35365 211989
rect 35399 211961 35427 211989
rect 35461 211961 35489 211989
rect 35523 211961 35551 211989
rect 35337 203147 35365 203175
rect 35399 203147 35427 203175
rect 35461 203147 35489 203175
rect 35523 203147 35551 203175
rect 35337 203085 35365 203113
rect 35399 203085 35427 203113
rect 35461 203085 35489 203113
rect 35523 203085 35551 203113
rect 35337 203023 35365 203051
rect 35399 203023 35427 203051
rect 35461 203023 35489 203051
rect 35523 203023 35551 203051
rect 35337 202961 35365 202989
rect 35399 202961 35427 202989
rect 35461 202961 35489 202989
rect 35523 202961 35551 202989
rect 35337 194147 35365 194175
rect 35399 194147 35427 194175
rect 35461 194147 35489 194175
rect 35523 194147 35551 194175
rect 35337 194085 35365 194113
rect 35399 194085 35427 194113
rect 35461 194085 35489 194113
rect 35523 194085 35551 194113
rect 35337 194023 35365 194051
rect 35399 194023 35427 194051
rect 35461 194023 35489 194051
rect 35523 194023 35551 194051
rect 35337 193961 35365 193989
rect 35399 193961 35427 193989
rect 35461 193961 35489 193989
rect 35523 193961 35551 193989
rect 35337 185147 35365 185175
rect 35399 185147 35427 185175
rect 35461 185147 35489 185175
rect 35523 185147 35551 185175
rect 35337 185085 35365 185113
rect 35399 185085 35427 185113
rect 35461 185085 35489 185113
rect 35523 185085 35551 185113
rect 35337 185023 35365 185051
rect 35399 185023 35427 185051
rect 35461 185023 35489 185051
rect 35523 185023 35551 185051
rect 35337 184961 35365 184989
rect 35399 184961 35427 184989
rect 35461 184961 35489 184989
rect 35523 184961 35551 184989
rect 35337 176147 35365 176175
rect 35399 176147 35427 176175
rect 35461 176147 35489 176175
rect 35523 176147 35551 176175
rect 35337 176085 35365 176113
rect 35399 176085 35427 176113
rect 35461 176085 35489 176113
rect 35523 176085 35551 176113
rect 35337 176023 35365 176051
rect 35399 176023 35427 176051
rect 35461 176023 35489 176051
rect 35523 176023 35551 176051
rect 35337 175961 35365 175989
rect 35399 175961 35427 175989
rect 35461 175961 35489 175989
rect 35523 175961 35551 175989
rect 48837 298578 48865 298606
rect 48899 298578 48927 298606
rect 48961 298578 48989 298606
rect 49023 298578 49051 298606
rect 48837 298516 48865 298544
rect 48899 298516 48927 298544
rect 48961 298516 48989 298544
rect 49023 298516 49051 298544
rect 48837 298454 48865 298482
rect 48899 298454 48927 298482
rect 48961 298454 48989 298482
rect 49023 298454 49051 298482
rect 48837 298392 48865 298420
rect 48899 298392 48927 298420
rect 48961 298392 48989 298420
rect 49023 298392 49051 298420
rect 48837 290147 48865 290175
rect 48899 290147 48927 290175
rect 48961 290147 48989 290175
rect 49023 290147 49051 290175
rect 48837 290085 48865 290113
rect 48899 290085 48927 290113
rect 48961 290085 48989 290113
rect 49023 290085 49051 290113
rect 48837 290023 48865 290051
rect 48899 290023 48927 290051
rect 48961 290023 48989 290051
rect 49023 290023 49051 290051
rect 48837 289961 48865 289989
rect 48899 289961 48927 289989
rect 48961 289961 48989 289989
rect 49023 289961 49051 289989
rect 48837 281147 48865 281175
rect 48899 281147 48927 281175
rect 48961 281147 48989 281175
rect 49023 281147 49051 281175
rect 48837 281085 48865 281113
rect 48899 281085 48927 281113
rect 48961 281085 48989 281113
rect 49023 281085 49051 281113
rect 48837 281023 48865 281051
rect 48899 281023 48927 281051
rect 48961 281023 48989 281051
rect 49023 281023 49051 281051
rect 48837 280961 48865 280989
rect 48899 280961 48927 280989
rect 48961 280961 48989 280989
rect 49023 280961 49051 280989
rect 48837 272147 48865 272175
rect 48899 272147 48927 272175
rect 48961 272147 48989 272175
rect 49023 272147 49051 272175
rect 48837 272085 48865 272113
rect 48899 272085 48927 272113
rect 48961 272085 48989 272113
rect 49023 272085 49051 272113
rect 48837 272023 48865 272051
rect 48899 272023 48927 272051
rect 48961 272023 48989 272051
rect 49023 272023 49051 272051
rect 48837 271961 48865 271989
rect 48899 271961 48927 271989
rect 48961 271961 48989 271989
rect 49023 271961 49051 271989
rect 48837 263147 48865 263175
rect 48899 263147 48927 263175
rect 48961 263147 48989 263175
rect 49023 263147 49051 263175
rect 48837 263085 48865 263113
rect 48899 263085 48927 263113
rect 48961 263085 48989 263113
rect 49023 263085 49051 263113
rect 48837 263023 48865 263051
rect 48899 263023 48927 263051
rect 48961 263023 48989 263051
rect 49023 263023 49051 263051
rect 48837 262961 48865 262989
rect 48899 262961 48927 262989
rect 48961 262961 48989 262989
rect 49023 262961 49051 262989
rect 48837 254147 48865 254175
rect 48899 254147 48927 254175
rect 48961 254147 48989 254175
rect 49023 254147 49051 254175
rect 48837 254085 48865 254113
rect 48899 254085 48927 254113
rect 48961 254085 48989 254113
rect 49023 254085 49051 254113
rect 48837 254023 48865 254051
rect 48899 254023 48927 254051
rect 48961 254023 48989 254051
rect 49023 254023 49051 254051
rect 48837 253961 48865 253989
rect 48899 253961 48927 253989
rect 48961 253961 48989 253989
rect 49023 253961 49051 253989
rect 48837 245147 48865 245175
rect 48899 245147 48927 245175
rect 48961 245147 48989 245175
rect 49023 245147 49051 245175
rect 48837 245085 48865 245113
rect 48899 245085 48927 245113
rect 48961 245085 48989 245113
rect 49023 245085 49051 245113
rect 48837 245023 48865 245051
rect 48899 245023 48927 245051
rect 48961 245023 48989 245051
rect 49023 245023 49051 245051
rect 48837 244961 48865 244989
rect 48899 244961 48927 244989
rect 48961 244961 48989 244989
rect 49023 244961 49051 244989
rect 48837 236147 48865 236175
rect 48899 236147 48927 236175
rect 48961 236147 48989 236175
rect 49023 236147 49051 236175
rect 48837 236085 48865 236113
rect 48899 236085 48927 236113
rect 48961 236085 48989 236113
rect 49023 236085 49051 236113
rect 48837 236023 48865 236051
rect 48899 236023 48927 236051
rect 48961 236023 48989 236051
rect 49023 236023 49051 236051
rect 48837 235961 48865 235989
rect 48899 235961 48927 235989
rect 48961 235961 48989 235989
rect 49023 235961 49051 235989
rect 48837 227147 48865 227175
rect 48899 227147 48927 227175
rect 48961 227147 48989 227175
rect 49023 227147 49051 227175
rect 48837 227085 48865 227113
rect 48899 227085 48927 227113
rect 48961 227085 48989 227113
rect 49023 227085 49051 227113
rect 48837 227023 48865 227051
rect 48899 227023 48927 227051
rect 48961 227023 48989 227051
rect 49023 227023 49051 227051
rect 48837 226961 48865 226989
rect 48899 226961 48927 226989
rect 48961 226961 48989 226989
rect 49023 226961 49051 226989
rect 48837 218147 48865 218175
rect 48899 218147 48927 218175
rect 48961 218147 48989 218175
rect 49023 218147 49051 218175
rect 48837 218085 48865 218113
rect 48899 218085 48927 218113
rect 48961 218085 48989 218113
rect 49023 218085 49051 218113
rect 48837 218023 48865 218051
rect 48899 218023 48927 218051
rect 48961 218023 48989 218051
rect 49023 218023 49051 218051
rect 48837 217961 48865 217989
rect 48899 217961 48927 217989
rect 48961 217961 48989 217989
rect 49023 217961 49051 217989
rect 48837 209147 48865 209175
rect 48899 209147 48927 209175
rect 48961 209147 48989 209175
rect 49023 209147 49051 209175
rect 48837 209085 48865 209113
rect 48899 209085 48927 209113
rect 48961 209085 48989 209113
rect 49023 209085 49051 209113
rect 48837 209023 48865 209051
rect 48899 209023 48927 209051
rect 48961 209023 48989 209051
rect 49023 209023 49051 209051
rect 48837 208961 48865 208989
rect 48899 208961 48927 208989
rect 48961 208961 48989 208989
rect 49023 208961 49051 208989
rect 48837 200147 48865 200175
rect 48899 200147 48927 200175
rect 48961 200147 48989 200175
rect 49023 200147 49051 200175
rect 48837 200085 48865 200113
rect 48899 200085 48927 200113
rect 48961 200085 48989 200113
rect 49023 200085 49051 200113
rect 48837 200023 48865 200051
rect 48899 200023 48927 200051
rect 48961 200023 48989 200051
rect 49023 200023 49051 200051
rect 48837 199961 48865 199989
rect 48899 199961 48927 199989
rect 48961 199961 48989 199989
rect 49023 199961 49051 199989
rect 48837 191147 48865 191175
rect 48899 191147 48927 191175
rect 48961 191147 48989 191175
rect 49023 191147 49051 191175
rect 48837 191085 48865 191113
rect 48899 191085 48927 191113
rect 48961 191085 48989 191113
rect 49023 191085 49051 191113
rect 48837 191023 48865 191051
rect 48899 191023 48927 191051
rect 48961 191023 48989 191051
rect 49023 191023 49051 191051
rect 48837 190961 48865 190989
rect 48899 190961 48927 190989
rect 48961 190961 48989 190989
rect 49023 190961 49051 190989
rect 48837 182147 48865 182175
rect 48899 182147 48927 182175
rect 48961 182147 48989 182175
rect 49023 182147 49051 182175
rect 48837 182085 48865 182113
rect 48899 182085 48927 182113
rect 48961 182085 48989 182113
rect 49023 182085 49051 182113
rect 48837 182023 48865 182051
rect 48899 182023 48927 182051
rect 48961 182023 48989 182051
rect 49023 182023 49051 182051
rect 48837 181961 48865 181989
rect 48899 181961 48927 181989
rect 48961 181961 48989 181989
rect 49023 181961 49051 181989
rect 38979 173147 39007 173175
rect 39041 173147 39069 173175
rect 38979 173085 39007 173113
rect 39041 173085 39069 173113
rect 38979 173023 39007 173051
rect 39041 173023 39069 173051
rect 38979 172961 39007 172989
rect 39041 172961 39069 172989
rect 48837 173147 48865 173175
rect 48899 173147 48927 173175
rect 48961 173147 48989 173175
rect 49023 173147 49051 173175
rect 48837 173085 48865 173113
rect 48899 173085 48927 173113
rect 48961 173085 48989 173113
rect 49023 173085 49051 173113
rect 48837 173023 48865 173051
rect 48899 173023 48927 173051
rect 48961 173023 48989 173051
rect 49023 173023 49051 173051
rect 48837 172961 48865 172989
rect 48899 172961 48927 172989
rect 48961 172961 48989 172989
rect 49023 172961 49051 172989
rect 35337 167147 35365 167175
rect 35399 167147 35427 167175
rect 35461 167147 35489 167175
rect 35523 167147 35551 167175
rect 35337 167085 35365 167113
rect 35399 167085 35427 167113
rect 35461 167085 35489 167113
rect 35523 167085 35551 167113
rect 35337 167023 35365 167051
rect 35399 167023 35427 167051
rect 35461 167023 35489 167051
rect 35523 167023 35551 167051
rect 35337 166961 35365 166989
rect 35399 166961 35427 166989
rect 35461 166961 35489 166989
rect 35523 166961 35551 166989
rect 46659 167147 46687 167175
rect 46721 167147 46749 167175
rect 46659 167085 46687 167113
rect 46721 167085 46749 167113
rect 46659 167023 46687 167051
rect 46721 167023 46749 167051
rect 46659 166961 46687 166989
rect 46721 166961 46749 166989
rect 38979 164147 39007 164175
rect 39041 164147 39069 164175
rect 38979 164085 39007 164113
rect 39041 164085 39069 164113
rect 38979 164023 39007 164051
rect 39041 164023 39069 164051
rect 38979 163961 39007 163989
rect 39041 163961 39069 163989
rect 48837 164147 48865 164175
rect 48899 164147 48927 164175
rect 48961 164147 48989 164175
rect 49023 164147 49051 164175
rect 48837 164085 48865 164113
rect 48899 164085 48927 164113
rect 48961 164085 48989 164113
rect 49023 164085 49051 164113
rect 48837 164023 48865 164051
rect 48899 164023 48927 164051
rect 48961 164023 48989 164051
rect 49023 164023 49051 164051
rect 48837 163961 48865 163989
rect 48899 163961 48927 163989
rect 48961 163961 48989 163989
rect 49023 163961 49051 163989
rect 35337 158147 35365 158175
rect 35399 158147 35427 158175
rect 35461 158147 35489 158175
rect 35523 158147 35551 158175
rect 35337 158085 35365 158113
rect 35399 158085 35427 158113
rect 35461 158085 35489 158113
rect 35523 158085 35551 158113
rect 35337 158023 35365 158051
rect 35399 158023 35427 158051
rect 35461 158023 35489 158051
rect 35523 158023 35551 158051
rect 35337 157961 35365 157989
rect 35399 157961 35427 157989
rect 35461 157961 35489 157989
rect 35523 157961 35551 157989
rect 46659 158147 46687 158175
rect 46721 158147 46749 158175
rect 46659 158085 46687 158113
rect 46721 158085 46749 158113
rect 46659 158023 46687 158051
rect 46721 158023 46749 158051
rect 46659 157961 46687 157989
rect 46721 157961 46749 157989
rect 38979 155147 39007 155175
rect 39041 155147 39069 155175
rect 38979 155085 39007 155113
rect 39041 155085 39069 155113
rect 38979 155023 39007 155051
rect 39041 155023 39069 155051
rect 38979 154961 39007 154989
rect 39041 154961 39069 154989
rect 48837 155147 48865 155175
rect 48899 155147 48927 155175
rect 48961 155147 48989 155175
rect 49023 155147 49051 155175
rect 48837 155085 48865 155113
rect 48899 155085 48927 155113
rect 48961 155085 48989 155113
rect 49023 155085 49051 155113
rect 48837 155023 48865 155051
rect 48899 155023 48927 155051
rect 48961 155023 48989 155051
rect 49023 155023 49051 155051
rect 48837 154961 48865 154989
rect 48899 154961 48927 154989
rect 48961 154961 48989 154989
rect 49023 154961 49051 154989
rect 35337 149147 35365 149175
rect 35399 149147 35427 149175
rect 35461 149147 35489 149175
rect 35523 149147 35551 149175
rect 35337 149085 35365 149113
rect 35399 149085 35427 149113
rect 35461 149085 35489 149113
rect 35523 149085 35551 149113
rect 35337 149023 35365 149051
rect 35399 149023 35427 149051
rect 35461 149023 35489 149051
rect 35523 149023 35551 149051
rect 35337 148961 35365 148989
rect 35399 148961 35427 148989
rect 35461 148961 35489 148989
rect 35523 148961 35551 148989
rect 46659 149147 46687 149175
rect 46721 149147 46749 149175
rect 46659 149085 46687 149113
rect 46721 149085 46749 149113
rect 46659 149023 46687 149051
rect 46721 149023 46749 149051
rect 46659 148961 46687 148989
rect 46721 148961 46749 148989
rect 38979 146147 39007 146175
rect 39041 146147 39069 146175
rect 38979 146085 39007 146113
rect 39041 146085 39069 146113
rect 38979 146023 39007 146051
rect 39041 146023 39069 146051
rect 38979 145961 39007 145989
rect 39041 145961 39069 145989
rect 48837 146147 48865 146175
rect 48899 146147 48927 146175
rect 48961 146147 48989 146175
rect 49023 146147 49051 146175
rect 48837 146085 48865 146113
rect 48899 146085 48927 146113
rect 48961 146085 48989 146113
rect 49023 146085 49051 146113
rect 48837 146023 48865 146051
rect 48899 146023 48927 146051
rect 48961 146023 48989 146051
rect 49023 146023 49051 146051
rect 48837 145961 48865 145989
rect 48899 145961 48927 145989
rect 48961 145961 48989 145989
rect 49023 145961 49051 145989
rect 35337 140147 35365 140175
rect 35399 140147 35427 140175
rect 35461 140147 35489 140175
rect 35523 140147 35551 140175
rect 35337 140085 35365 140113
rect 35399 140085 35427 140113
rect 35461 140085 35489 140113
rect 35523 140085 35551 140113
rect 35337 140023 35365 140051
rect 35399 140023 35427 140051
rect 35461 140023 35489 140051
rect 35523 140023 35551 140051
rect 35337 139961 35365 139989
rect 35399 139961 35427 139989
rect 35461 139961 35489 139989
rect 35523 139961 35551 139989
rect 46659 140147 46687 140175
rect 46721 140147 46749 140175
rect 46659 140085 46687 140113
rect 46721 140085 46749 140113
rect 46659 140023 46687 140051
rect 46721 140023 46749 140051
rect 46659 139961 46687 139989
rect 46721 139961 46749 139989
rect 38979 137147 39007 137175
rect 39041 137147 39069 137175
rect 38979 137085 39007 137113
rect 39041 137085 39069 137113
rect 38979 137023 39007 137051
rect 39041 137023 39069 137051
rect 38979 136961 39007 136989
rect 39041 136961 39069 136989
rect 48837 137147 48865 137175
rect 48899 137147 48927 137175
rect 48961 137147 48989 137175
rect 49023 137147 49051 137175
rect 48837 137085 48865 137113
rect 48899 137085 48927 137113
rect 48961 137085 48989 137113
rect 49023 137085 49051 137113
rect 48837 137023 48865 137051
rect 48899 137023 48927 137051
rect 48961 137023 48989 137051
rect 49023 137023 49051 137051
rect 48837 136961 48865 136989
rect 48899 136961 48927 136989
rect 48961 136961 48989 136989
rect 49023 136961 49051 136989
rect 35337 131147 35365 131175
rect 35399 131147 35427 131175
rect 35461 131147 35489 131175
rect 35523 131147 35551 131175
rect 35337 131085 35365 131113
rect 35399 131085 35427 131113
rect 35461 131085 35489 131113
rect 35523 131085 35551 131113
rect 35337 131023 35365 131051
rect 35399 131023 35427 131051
rect 35461 131023 35489 131051
rect 35523 131023 35551 131051
rect 35337 130961 35365 130989
rect 35399 130961 35427 130989
rect 35461 130961 35489 130989
rect 35523 130961 35551 130989
rect 46659 131147 46687 131175
rect 46721 131147 46749 131175
rect 46659 131085 46687 131113
rect 46721 131085 46749 131113
rect 46659 131023 46687 131051
rect 46721 131023 46749 131051
rect 46659 130961 46687 130989
rect 46721 130961 46749 130989
rect 38979 128147 39007 128175
rect 39041 128147 39069 128175
rect 38979 128085 39007 128113
rect 39041 128085 39069 128113
rect 38979 128023 39007 128051
rect 39041 128023 39069 128051
rect 38979 127961 39007 127989
rect 39041 127961 39069 127989
rect 48837 128147 48865 128175
rect 48899 128147 48927 128175
rect 48961 128147 48989 128175
rect 49023 128147 49051 128175
rect 48837 128085 48865 128113
rect 48899 128085 48927 128113
rect 48961 128085 48989 128113
rect 49023 128085 49051 128113
rect 48837 128023 48865 128051
rect 48899 128023 48927 128051
rect 48961 128023 48989 128051
rect 49023 128023 49051 128051
rect 48837 127961 48865 127989
rect 48899 127961 48927 127989
rect 48961 127961 48989 127989
rect 49023 127961 49051 127989
rect 35337 122147 35365 122175
rect 35399 122147 35427 122175
rect 35461 122147 35489 122175
rect 35523 122147 35551 122175
rect 35337 122085 35365 122113
rect 35399 122085 35427 122113
rect 35461 122085 35489 122113
rect 35523 122085 35551 122113
rect 35337 122023 35365 122051
rect 35399 122023 35427 122051
rect 35461 122023 35489 122051
rect 35523 122023 35551 122051
rect 35337 121961 35365 121989
rect 35399 121961 35427 121989
rect 35461 121961 35489 121989
rect 35523 121961 35551 121989
rect 46659 122147 46687 122175
rect 46721 122147 46749 122175
rect 46659 122085 46687 122113
rect 46721 122085 46749 122113
rect 46659 122023 46687 122051
rect 46721 122023 46749 122051
rect 46659 121961 46687 121989
rect 46721 121961 46749 121989
rect 38979 119147 39007 119175
rect 39041 119147 39069 119175
rect 38979 119085 39007 119113
rect 39041 119085 39069 119113
rect 38979 119023 39007 119051
rect 39041 119023 39069 119051
rect 38979 118961 39007 118989
rect 39041 118961 39069 118989
rect 48837 119147 48865 119175
rect 48899 119147 48927 119175
rect 48961 119147 48989 119175
rect 49023 119147 49051 119175
rect 48837 119085 48865 119113
rect 48899 119085 48927 119113
rect 48961 119085 48989 119113
rect 49023 119085 49051 119113
rect 48837 119023 48865 119051
rect 48899 119023 48927 119051
rect 48961 119023 48989 119051
rect 49023 119023 49051 119051
rect 48837 118961 48865 118989
rect 48899 118961 48927 118989
rect 48961 118961 48989 118989
rect 49023 118961 49051 118989
rect 35337 113147 35365 113175
rect 35399 113147 35427 113175
rect 35461 113147 35489 113175
rect 35523 113147 35551 113175
rect 35337 113085 35365 113113
rect 35399 113085 35427 113113
rect 35461 113085 35489 113113
rect 35523 113085 35551 113113
rect 35337 113023 35365 113051
rect 35399 113023 35427 113051
rect 35461 113023 35489 113051
rect 35523 113023 35551 113051
rect 35337 112961 35365 112989
rect 35399 112961 35427 112989
rect 35461 112961 35489 112989
rect 35523 112961 35551 112989
rect 46659 113147 46687 113175
rect 46721 113147 46749 113175
rect 46659 113085 46687 113113
rect 46721 113085 46749 113113
rect 46659 113023 46687 113051
rect 46721 113023 46749 113051
rect 46659 112961 46687 112989
rect 46721 112961 46749 112989
rect 38979 110147 39007 110175
rect 39041 110147 39069 110175
rect 38979 110085 39007 110113
rect 39041 110085 39069 110113
rect 38979 110023 39007 110051
rect 39041 110023 39069 110051
rect 38979 109961 39007 109989
rect 39041 109961 39069 109989
rect 48837 110147 48865 110175
rect 48899 110147 48927 110175
rect 48961 110147 48989 110175
rect 49023 110147 49051 110175
rect 48837 110085 48865 110113
rect 48899 110085 48927 110113
rect 48961 110085 48989 110113
rect 49023 110085 49051 110113
rect 48837 110023 48865 110051
rect 48899 110023 48927 110051
rect 48961 110023 48989 110051
rect 49023 110023 49051 110051
rect 48837 109961 48865 109989
rect 48899 109961 48927 109989
rect 48961 109961 48989 109989
rect 49023 109961 49051 109989
rect 35337 104147 35365 104175
rect 35399 104147 35427 104175
rect 35461 104147 35489 104175
rect 35523 104147 35551 104175
rect 35337 104085 35365 104113
rect 35399 104085 35427 104113
rect 35461 104085 35489 104113
rect 35523 104085 35551 104113
rect 35337 104023 35365 104051
rect 35399 104023 35427 104051
rect 35461 104023 35489 104051
rect 35523 104023 35551 104051
rect 35337 103961 35365 103989
rect 35399 103961 35427 103989
rect 35461 103961 35489 103989
rect 35523 103961 35551 103989
rect 46659 104147 46687 104175
rect 46721 104147 46749 104175
rect 46659 104085 46687 104113
rect 46721 104085 46749 104113
rect 46659 104023 46687 104051
rect 46721 104023 46749 104051
rect 46659 103961 46687 103989
rect 46721 103961 46749 103989
rect 38979 101147 39007 101175
rect 39041 101147 39069 101175
rect 38979 101085 39007 101113
rect 39041 101085 39069 101113
rect 38979 101023 39007 101051
rect 39041 101023 39069 101051
rect 38979 100961 39007 100989
rect 39041 100961 39069 100989
rect 48837 101147 48865 101175
rect 48899 101147 48927 101175
rect 48961 101147 48989 101175
rect 49023 101147 49051 101175
rect 48837 101085 48865 101113
rect 48899 101085 48927 101113
rect 48961 101085 48989 101113
rect 49023 101085 49051 101113
rect 48837 101023 48865 101051
rect 48899 101023 48927 101051
rect 48961 101023 48989 101051
rect 49023 101023 49051 101051
rect 48837 100961 48865 100989
rect 48899 100961 48927 100989
rect 48961 100961 48989 100989
rect 49023 100961 49051 100989
rect 35337 95147 35365 95175
rect 35399 95147 35427 95175
rect 35461 95147 35489 95175
rect 35523 95147 35551 95175
rect 35337 95085 35365 95113
rect 35399 95085 35427 95113
rect 35461 95085 35489 95113
rect 35523 95085 35551 95113
rect 35337 95023 35365 95051
rect 35399 95023 35427 95051
rect 35461 95023 35489 95051
rect 35523 95023 35551 95051
rect 35337 94961 35365 94989
rect 35399 94961 35427 94989
rect 35461 94961 35489 94989
rect 35523 94961 35551 94989
rect 46659 95147 46687 95175
rect 46721 95147 46749 95175
rect 46659 95085 46687 95113
rect 46721 95085 46749 95113
rect 46659 95023 46687 95051
rect 46721 95023 46749 95051
rect 46659 94961 46687 94989
rect 46721 94961 46749 94989
rect 38979 92147 39007 92175
rect 39041 92147 39069 92175
rect 38979 92085 39007 92113
rect 39041 92085 39069 92113
rect 38979 92023 39007 92051
rect 39041 92023 39069 92051
rect 38979 91961 39007 91989
rect 39041 91961 39069 91989
rect 48837 92147 48865 92175
rect 48899 92147 48927 92175
rect 48961 92147 48989 92175
rect 49023 92147 49051 92175
rect 48837 92085 48865 92113
rect 48899 92085 48927 92113
rect 48961 92085 48989 92113
rect 49023 92085 49051 92113
rect 48837 92023 48865 92051
rect 48899 92023 48927 92051
rect 48961 92023 48989 92051
rect 49023 92023 49051 92051
rect 48837 91961 48865 91989
rect 48899 91961 48927 91989
rect 48961 91961 48989 91989
rect 49023 91961 49051 91989
rect 35337 86147 35365 86175
rect 35399 86147 35427 86175
rect 35461 86147 35489 86175
rect 35523 86147 35551 86175
rect 35337 86085 35365 86113
rect 35399 86085 35427 86113
rect 35461 86085 35489 86113
rect 35523 86085 35551 86113
rect 35337 86023 35365 86051
rect 35399 86023 35427 86051
rect 35461 86023 35489 86051
rect 35523 86023 35551 86051
rect 35337 85961 35365 85989
rect 35399 85961 35427 85989
rect 35461 85961 35489 85989
rect 35523 85961 35551 85989
rect 46659 86147 46687 86175
rect 46721 86147 46749 86175
rect 46659 86085 46687 86113
rect 46721 86085 46749 86113
rect 46659 86023 46687 86051
rect 46721 86023 46749 86051
rect 46659 85961 46687 85989
rect 46721 85961 46749 85989
rect 38979 83147 39007 83175
rect 39041 83147 39069 83175
rect 38979 83085 39007 83113
rect 39041 83085 39069 83113
rect 38979 83023 39007 83051
rect 39041 83023 39069 83051
rect 38979 82961 39007 82989
rect 39041 82961 39069 82989
rect 48837 83147 48865 83175
rect 48899 83147 48927 83175
rect 48961 83147 48989 83175
rect 49023 83147 49051 83175
rect 48837 83085 48865 83113
rect 48899 83085 48927 83113
rect 48961 83085 48989 83113
rect 49023 83085 49051 83113
rect 48837 83023 48865 83051
rect 48899 83023 48927 83051
rect 48961 83023 48989 83051
rect 49023 83023 49051 83051
rect 48837 82961 48865 82989
rect 48899 82961 48927 82989
rect 48961 82961 48989 82989
rect 49023 82961 49051 82989
rect 35337 77147 35365 77175
rect 35399 77147 35427 77175
rect 35461 77147 35489 77175
rect 35523 77147 35551 77175
rect 35337 77085 35365 77113
rect 35399 77085 35427 77113
rect 35461 77085 35489 77113
rect 35523 77085 35551 77113
rect 35337 77023 35365 77051
rect 35399 77023 35427 77051
rect 35461 77023 35489 77051
rect 35523 77023 35551 77051
rect 35337 76961 35365 76989
rect 35399 76961 35427 76989
rect 35461 76961 35489 76989
rect 35523 76961 35551 76989
rect 46659 77147 46687 77175
rect 46721 77147 46749 77175
rect 46659 77085 46687 77113
rect 46721 77085 46749 77113
rect 46659 77023 46687 77051
rect 46721 77023 46749 77051
rect 46659 76961 46687 76989
rect 46721 76961 46749 76989
rect 38979 74147 39007 74175
rect 39041 74147 39069 74175
rect 38979 74085 39007 74113
rect 39041 74085 39069 74113
rect 38979 74023 39007 74051
rect 39041 74023 39069 74051
rect 38979 73961 39007 73989
rect 39041 73961 39069 73989
rect 48837 74147 48865 74175
rect 48899 74147 48927 74175
rect 48961 74147 48989 74175
rect 49023 74147 49051 74175
rect 48837 74085 48865 74113
rect 48899 74085 48927 74113
rect 48961 74085 48989 74113
rect 49023 74085 49051 74113
rect 48837 74023 48865 74051
rect 48899 74023 48927 74051
rect 48961 74023 48989 74051
rect 49023 74023 49051 74051
rect 48837 73961 48865 73989
rect 48899 73961 48927 73989
rect 48961 73961 48989 73989
rect 49023 73961 49051 73989
rect 35337 68147 35365 68175
rect 35399 68147 35427 68175
rect 35461 68147 35489 68175
rect 35523 68147 35551 68175
rect 35337 68085 35365 68113
rect 35399 68085 35427 68113
rect 35461 68085 35489 68113
rect 35523 68085 35551 68113
rect 35337 68023 35365 68051
rect 35399 68023 35427 68051
rect 35461 68023 35489 68051
rect 35523 68023 35551 68051
rect 35337 67961 35365 67989
rect 35399 67961 35427 67989
rect 35461 67961 35489 67989
rect 35523 67961 35551 67989
rect 46659 68147 46687 68175
rect 46721 68147 46749 68175
rect 46659 68085 46687 68113
rect 46721 68085 46749 68113
rect 46659 68023 46687 68051
rect 46721 68023 46749 68051
rect 46659 67961 46687 67989
rect 46721 67961 46749 67989
rect 38979 65147 39007 65175
rect 39041 65147 39069 65175
rect 38979 65085 39007 65113
rect 39041 65085 39069 65113
rect 38979 65023 39007 65051
rect 39041 65023 39069 65051
rect 38979 64961 39007 64989
rect 39041 64961 39069 64989
rect 48837 65147 48865 65175
rect 48899 65147 48927 65175
rect 48961 65147 48989 65175
rect 49023 65147 49051 65175
rect 48837 65085 48865 65113
rect 48899 65085 48927 65113
rect 48961 65085 48989 65113
rect 49023 65085 49051 65113
rect 48837 65023 48865 65051
rect 48899 65023 48927 65051
rect 48961 65023 48989 65051
rect 49023 65023 49051 65051
rect 48837 64961 48865 64989
rect 48899 64961 48927 64989
rect 48961 64961 48989 64989
rect 49023 64961 49051 64989
rect 35337 59147 35365 59175
rect 35399 59147 35427 59175
rect 35461 59147 35489 59175
rect 35523 59147 35551 59175
rect 35337 59085 35365 59113
rect 35399 59085 35427 59113
rect 35461 59085 35489 59113
rect 35523 59085 35551 59113
rect 35337 59023 35365 59051
rect 35399 59023 35427 59051
rect 35461 59023 35489 59051
rect 35523 59023 35551 59051
rect 35337 58961 35365 58989
rect 35399 58961 35427 58989
rect 35461 58961 35489 58989
rect 35523 58961 35551 58989
rect 46659 59147 46687 59175
rect 46721 59147 46749 59175
rect 46659 59085 46687 59113
rect 46721 59085 46749 59113
rect 46659 59023 46687 59051
rect 46721 59023 46749 59051
rect 46659 58961 46687 58989
rect 46721 58961 46749 58989
rect 38979 56147 39007 56175
rect 39041 56147 39069 56175
rect 38979 56085 39007 56113
rect 39041 56085 39069 56113
rect 38979 56023 39007 56051
rect 39041 56023 39069 56051
rect 38979 55961 39007 55989
rect 39041 55961 39069 55989
rect 48837 56147 48865 56175
rect 48899 56147 48927 56175
rect 48961 56147 48989 56175
rect 49023 56147 49051 56175
rect 48837 56085 48865 56113
rect 48899 56085 48927 56113
rect 48961 56085 48989 56113
rect 49023 56085 49051 56113
rect 48837 56023 48865 56051
rect 48899 56023 48927 56051
rect 48961 56023 48989 56051
rect 49023 56023 49051 56051
rect 48837 55961 48865 55989
rect 48899 55961 48927 55989
rect 48961 55961 48989 55989
rect 49023 55961 49051 55989
rect 35337 50147 35365 50175
rect 35399 50147 35427 50175
rect 35461 50147 35489 50175
rect 35523 50147 35551 50175
rect 35337 50085 35365 50113
rect 35399 50085 35427 50113
rect 35461 50085 35489 50113
rect 35523 50085 35551 50113
rect 35337 50023 35365 50051
rect 35399 50023 35427 50051
rect 35461 50023 35489 50051
rect 35523 50023 35551 50051
rect 35337 49961 35365 49989
rect 35399 49961 35427 49989
rect 35461 49961 35489 49989
rect 35523 49961 35551 49989
rect 46659 50147 46687 50175
rect 46721 50147 46749 50175
rect 46659 50085 46687 50113
rect 46721 50085 46749 50113
rect 46659 50023 46687 50051
rect 46721 50023 46749 50051
rect 46659 49961 46687 49989
rect 46721 49961 46749 49989
rect 38979 47147 39007 47175
rect 39041 47147 39069 47175
rect 38979 47085 39007 47113
rect 39041 47085 39069 47113
rect 38979 47023 39007 47051
rect 39041 47023 39069 47051
rect 38979 46961 39007 46989
rect 39041 46961 39069 46989
rect 48837 47147 48865 47175
rect 48899 47147 48927 47175
rect 48961 47147 48989 47175
rect 49023 47147 49051 47175
rect 48837 47085 48865 47113
rect 48899 47085 48927 47113
rect 48961 47085 48989 47113
rect 49023 47085 49051 47113
rect 48837 47023 48865 47051
rect 48899 47023 48927 47051
rect 48961 47023 48989 47051
rect 49023 47023 49051 47051
rect 48837 46961 48865 46989
rect 48899 46961 48927 46989
rect 48961 46961 48989 46989
rect 49023 46961 49051 46989
rect 35337 41147 35365 41175
rect 35399 41147 35427 41175
rect 35461 41147 35489 41175
rect 35523 41147 35551 41175
rect 35337 41085 35365 41113
rect 35399 41085 35427 41113
rect 35461 41085 35489 41113
rect 35523 41085 35551 41113
rect 35337 41023 35365 41051
rect 35399 41023 35427 41051
rect 35461 41023 35489 41051
rect 35523 41023 35551 41051
rect 35337 40961 35365 40989
rect 35399 40961 35427 40989
rect 35461 40961 35489 40989
rect 35523 40961 35551 40989
rect 46659 41147 46687 41175
rect 46721 41147 46749 41175
rect 46659 41085 46687 41113
rect 46721 41085 46749 41113
rect 46659 41023 46687 41051
rect 46721 41023 46749 41051
rect 46659 40961 46687 40989
rect 46721 40961 46749 40989
rect 38979 38147 39007 38175
rect 39041 38147 39069 38175
rect 38979 38085 39007 38113
rect 39041 38085 39069 38113
rect 38979 38023 39007 38051
rect 39041 38023 39069 38051
rect 38979 37961 39007 37989
rect 39041 37961 39069 37989
rect 48837 38147 48865 38175
rect 48899 38147 48927 38175
rect 48961 38147 48989 38175
rect 49023 38147 49051 38175
rect 48837 38085 48865 38113
rect 48899 38085 48927 38113
rect 48961 38085 48989 38113
rect 49023 38085 49051 38113
rect 48837 38023 48865 38051
rect 48899 38023 48927 38051
rect 48961 38023 48989 38051
rect 49023 38023 49051 38051
rect 48837 37961 48865 37989
rect 48899 37961 48927 37989
rect 48961 37961 48989 37989
rect 49023 37961 49051 37989
rect 35337 32147 35365 32175
rect 35399 32147 35427 32175
rect 35461 32147 35489 32175
rect 35523 32147 35551 32175
rect 35337 32085 35365 32113
rect 35399 32085 35427 32113
rect 35461 32085 35489 32113
rect 35523 32085 35551 32113
rect 35337 32023 35365 32051
rect 35399 32023 35427 32051
rect 35461 32023 35489 32051
rect 35523 32023 35551 32051
rect 35337 31961 35365 31989
rect 35399 31961 35427 31989
rect 35461 31961 35489 31989
rect 35523 31961 35551 31989
rect 46659 32147 46687 32175
rect 46721 32147 46749 32175
rect 46659 32085 46687 32113
rect 46721 32085 46749 32113
rect 46659 32023 46687 32051
rect 46721 32023 46749 32051
rect 46659 31961 46687 31989
rect 46721 31961 46749 31989
rect 38979 29147 39007 29175
rect 39041 29147 39069 29175
rect 38979 29085 39007 29113
rect 39041 29085 39069 29113
rect 38979 29023 39007 29051
rect 39041 29023 39069 29051
rect 38979 28961 39007 28989
rect 39041 28961 39069 28989
rect 48837 29147 48865 29175
rect 48899 29147 48927 29175
rect 48961 29147 48989 29175
rect 49023 29147 49051 29175
rect 48837 29085 48865 29113
rect 48899 29085 48927 29113
rect 48961 29085 48989 29113
rect 49023 29085 49051 29113
rect 48837 29023 48865 29051
rect 48899 29023 48927 29051
rect 48961 29023 48989 29051
rect 49023 29023 49051 29051
rect 48837 28961 48865 28989
rect 48899 28961 48927 28989
rect 48961 28961 48989 28989
rect 49023 28961 49051 28989
rect 35337 23147 35365 23175
rect 35399 23147 35427 23175
rect 35461 23147 35489 23175
rect 35523 23147 35551 23175
rect 35337 23085 35365 23113
rect 35399 23085 35427 23113
rect 35461 23085 35489 23113
rect 35523 23085 35551 23113
rect 35337 23023 35365 23051
rect 35399 23023 35427 23051
rect 35461 23023 35489 23051
rect 35523 23023 35551 23051
rect 35337 22961 35365 22989
rect 35399 22961 35427 22989
rect 35461 22961 35489 22989
rect 35523 22961 35551 22989
rect 46659 23147 46687 23175
rect 46721 23147 46749 23175
rect 46659 23085 46687 23113
rect 46721 23085 46749 23113
rect 46659 23023 46687 23051
rect 46721 23023 46749 23051
rect 46659 22961 46687 22989
rect 46721 22961 46749 22989
rect 38979 20147 39007 20175
rect 39041 20147 39069 20175
rect 38979 20085 39007 20113
rect 39041 20085 39069 20113
rect 38979 20023 39007 20051
rect 39041 20023 39069 20051
rect 38979 19961 39007 19989
rect 39041 19961 39069 19989
rect 48837 20147 48865 20175
rect 48899 20147 48927 20175
rect 48961 20147 48989 20175
rect 49023 20147 49051 20175
rect 48837 20085 48865 20113
rect 48899 20085 48927 20113
rect 48961 20085 48989 20113
rect 49023 20085 49051 20113
rect 48837 20023 48865 20051
rect 48899 20023 48927 20051
rect 48961 20023 48989 20051
rect 49023 20023 49051 20051
rect 48837 19961 48865 19989
rect 48899 19961 48927 19989
rect 48961 19961 48989 19989
rect 49023 19961 49051 19989
rect 35337 14147 35365 14175
rect 35399 14147 35427 14175
rect 35461 14147 35489 14175
rect 35523 14147 35551 14175
rect 35337 14085 35365 14113
rect 35399 14085 35427 14113
rect 35461 14085 35489 14113
rect 35523 14085 35551 14113
rect 35337 14023 35365 14051
rect 35399 14023 35427 14051
rect 35461 14023 35489 14051
rect 35523 14023 35551 14051
rect 35337 13961 35365 13989
rect 35399 13961 35427 13989
rect 35461 13961 35489 13989
rect 35523 13961 35551 13989
rect 46659 14147 46687 14175
rect 46721 14147 46749 14175
rect 46659 14085 46687 14113
rect 46721 14085 46749 14113
rect 46659 14023 46687 14051
rect 46721 14023 46749 14051
rect 46659 13961 46687 13989
rect 46721 13961 46749 13989
rect 38979 11147 39007 11175
rect 39041 11147 39069 11175
rect 38979 11085 39007 11113
rect 39041 11085 39069 11113
rect 38979 11023 39007 11051
rect 39041 11023 39069 11051
rect 38979 10961 39007 10989
rect 39041 10961 39069 10989
rect 48837 11147 48865 11175
rect 48899 11147 48927 11175
rect 48961 11147 48989 11175
rect 49023 11147 49051 11175
rect 48837 11085 48865 11113
rect 48899 11085 48927 11113
rect 48961 11085 48989 11113
rect 49023 11085 49051 11113
rect 48837 11023 48865 11051
rect 48899 11023 48927 11051
rect 48961 11023 48989 11051
rect 49023 11023 49051 11051
rect 48837 10961 48865 10989
rect 48899 10961 48927 10989
rect 48961 10961 48989 10989
rect 49023 10961 49051 10989
rect 35337 5147 35365 5175
rect 35399 5147 35427 5175
rect 35461 5147 35489 5175
rect 35523 5147 35551 5175
rect 35337 5085 35365 5113
rect 35399 5085 35427 5113
rect 35461 5085 35489 5113
rect 35523 5085 35551 5113
rect 35337 5023 35365 5051
rect 35399 5023 35427 5051
rect 35461 5023 35489 5051
rect 35523 5023 35551 5051
rect 35337 4961 35365 4989
rect 35399 4961 35427 4989
rect 35461 4961 35489 4989
rect 35523 4961 35551 4989
rect 46659 5147 46687 5175
rect 46721 5147 46749 5175
rect 46659 5085 46687 5113
rect 46721 5085 46749 5113
rect 46659 5023 46687 5051
rect 46721 5023 46749 5051
rect 46659 4961 46687 4989
rect 46721 4961 46749 4989
rect 35337 -588 35365 -560
rect 35399 -588 35427 -560
rect 35461 -588 35489 -560
rect 35523 -588 35551 -560
rect 35337 -650 35365 -622
rect 35399 -650 35427 -622
rect 35461 -650 35489 -622
rect 35523 -650 35551 -622
rect 35337 -712 35365 -684
rect 35399 -712 35427 -684
rect 35461 -712 35489 -684
rect 35523 -712 35551 -684
rect 35337 -774 35365 -746
rect 35399 -774 35427 -746
rect 35461 -774 35489 -746
rect 35523 -774 35551 -746
rect 48837 2147 48865 2175
rect 48899 2147 48927 2175
rect 48961 2147 48989 2175
rect 49023 2147 49051 2175
rect 48837 2085 48865 2113
rect 48899 2085 48927 2113
rect 48961 2085 48989 2113
rect 49023 2085 49051 2113
rect 48837 2023 48865 2051
rect 48899 2023 48927 2051
rect 48961 2023 48989 2051
rect 49023 2023 49051 2051
rect 48837 1961 48865 1989
rect 48899 1961 48927 1989
rect 48961 1961 48989 1989
rect 49023 1961 49051 1989
rect 48837 -108 48865 -80
rect 48899 -108 48927 -80
rect 48961 -108 48989 -80
rect 49023 -108 49051 -80
rect 48837 -170 48865 -142
rect 48899 -170 48927 -142
rect 48961 -170 48989 -142
rect 49023 -170 49051 -142
rect 48837 -232 48865 -204
rect 48899 -232 48927 -204
rect 48961 -232 48989 -204
rect 49023 -232 49051 -204
rect 48837 -294 48865 -266
rect 48899 -294 48927 -266
rect 48961 -294 48989 -266
rect 49023 -294 49051 -266
rect 50697 299058 50725 299086
rect 50759 299058 50787 299086
rect 50821 299058 50849 299086
rect 50883 299058 50911 299086
rect 50697 298996 50725 299024
rect 50759 298996 50787 299024
rect 50821 298996 50849 299024
rect 50883 298996 50911 299024
rect 50697 298934 50725 298962
rect 50759 298934 50787 298962
rect 50821 298934 50849 298962
rect 50883 298934 50911 298962
rect 50697 298872 50725 298900
rect 50759 298872 50787 298900
rect 50821 298872 50849 298900
rect 50883 298872 50911 298900
rect 50697 293147 50725 293175
rect 50759 293147 50787 293175
rect 50821 293147 50849 293175
rect 50883 293147 50911 293175
rect 50697 293085 50725 293113
rect 50759 293085 50787 293113
rect 50821 293085 50849 293113
rect 50883 293085 50911 293113
rect 50697 293023 50725 293051
rect 50759 293023 50787 293051
rect 50821 293023 50849 293051
rect 50883 293023 50911 293051
rect 50697 292961 50725 292989
rect 50759 292961 50787 292989
rect 50821 292961 50849 292989
rect 50883 292961 50911 292989
rect 50697 284147 50725 284175
rect 50759 284147 50787 284175
rect 50821 284147 50849 284175
rect 50883 284147 50911 284175
rect 50697 284085 50725 284113
rect 50759 284085 50787 284113
rect 50821 284085 50849 284113
rect 50883 284085 50911 284113
rect 50697 284023 50725 284051
rect 50759 284023 50787 284051
rect 50821 284023 50849 284051
rect 50883 284023 50911 284051
rect 50697 283961 50725 283989
rect 50759 283961 50787 283989
rect 50821 283961 50849 283989
rect 50883 283961 50911 283989
rect 50697 275147 50725 275175
rect 50759 275147 50787 275175
rect 50821 275147 50849 275175
rect 50883 275147 50911 275175
rect 50697 275085 50725 275113
rect 50759 275085 50787 275113
rect 50821 275085 50849 275113
rect 50883 275085 50911 275113
rect 50697 275023 50725 275051
rect 50759 275023 50787 275051
rect 50821 275023 50849 275051
rect 50883 275023 50911 275051
rect 50697 274961 50725 274989
rect 50759 274961 50787 274989
rect 50821 274961 50849 274989
rect 50883 274961 50911 274989
rect 50697 266147 50725 266175
rect 50759 266147 50787 266175
rect 50821 266147 50849 266175
rect 50883 266147 50911 266175
rect 50697 266085 50725 266113
rect 50759 266085 50787 266113
rect 50821 266085 50849 266113
rect 50883 266085 50911 266113
rect 50697 266023 50725 266051
rect 50759 266023 50787 266051
rect 50821 266023 50849 266051
rect 50883 266023 50911 266051
rect 50697 265961 50725 265989
rect 50759 265961 50787 265989
rect 50821 265961 50849 265989
rect 50883 265961 50911 265989
rect 50697 257147 50725 257175
rect 50759 257147 50787 257175
rect 50821 257147 50849 257175
rect 50883 257147 50911 257175
rect 50697 257085 50725 257113
rect 50759 257085 50787 257113
rect 50821 257085 50849 257113
rect 50883 257085 50911 257113
rect 50697 257023 50725 257051
rect 50759 257023 50787 257051
rect 50821 257023 50849 257051
rect 50883 257023 50911 257051
rect 50697 256961 50725 256989
rect 50759 256961 50787 256989
rect 50821 256961 50849 256989
rect 50883 256961 50911 256989
rect 50697 248147 50725 248175
rect 50759 248147 50787 248175
rect 50821 248147 50849 248175
rect 50883 248147 50911 248175
rect 50697 248085 50725 248113
rect 50759 248085 50787 248113
rect 50821 248085 50849 248113
rect 50883 248085 50911 248113
rect 50697 248023 50725 248051
rect 50759 248023 50787 248051
rect 50821 248023 50849 248051
rect 50883 248023 50911 248051
rect 50697 247961 50725 247989
rect 50759 247961 50787 247989
rect 50821 247961 50849 247989
rect 50883 247961 50911 247989
rect 50697 239147 50725 239175
rect 50759 239147 50787 239175
rect 50821 239147 50849 239175
rect 50883 239147 50911 239175
rect 50697 239085 50725 239113
rect 50759 239085 50787 239113
rect 50821 239085 50849 239113
rect 50883 239085 50911 239113
rect 50697 239023 50725 239051
rect 50759 239023 50787 239051
rect 50821 239023 50849 239051
rect 50883 239023 50911 239051
rect 50697 238961 50725 238989
rect 50759 238961 50787 238989
rect 50821 238961 50849 238989
rect 50883 238961 50911 238989
rect 50697 230147 50725 230175
rect 50759 230147 50787 230175
rect 50821 230147 50849 230175
rect 50883 230147 50911 230175
rect 50697 230085 50725 230113
rect 50759 230085 50787 230113
rect 50821 230085 50849 230113
rect 50883 230085 50911 230113
rect 50697 230023 50725 230051
rect 50759 230023 50787 230051
rect 50821 230023 50849 230051
rect 50883 230023 50911 230051
rect 50697 229961 50725 229989
rect 50759 229961 50787 229989
rect 50821 229961 50849 229989
rect 50883 229961 50911 229989
rect 50697 221147 50725 221175
rect 50759 221147 50787 221175
rect 50821 221147 50849 221175
rect 50883 221147 50911 221175
rect 50697 221085 50725 221113
rect 50759 221085 50787 221113
rect 50821 221085 50849 221113
rect 50883 221085 50911 221113
rect 50697 221023 50725 221051
rect 50759 221023 50787 221051
rect 50821 221023 50849 221051
rect 50883 221023 50911 221051
rect 50697 220961 50725 220989
rect 50759 220961 50787 220989
rect 50821 220961 50849 220989
rect 50883 220961 50911 220989
rect 50697 212147 50725 212175
rect 50759 212147 50787 212175
rect 50821 212147 50849 212175
rect 50883 212147 50911 212175
rect 50697 212085 50725 212113
rect 50759 212085 50787 212113
rect 50821 212085 50849 212113
rect 50883 212085 50911 212113
rect 50697 212023 50725 212051
rect 50759 212023 50787 212051
rect 50821 212023 50849 212051
rect 50883 212023 50911 212051
rect 50697 211961 50725 211989
rect 50759 211961 50787 211989
rect 50821 211961 50849 211989
rect 50883 211961 50911 211989
rect 50697 203147 50725 203175
rect 50759 203147 50787 203175
rect 50821 203147 50849 203175
rect 50883 203147 50911 203175
rect 50697 203085 50725 203113
rect 50759 203085 50787 203113
rect 50821 203085 50849 203113
rect 50883 203085 50911 203113
rect 50697 203023 50725 203051
rect 50759 203023 50787 203051
rect 50821 203023 50849 203051
rect 50883 203023 50911 203051
rect 50697 202961 50725 202989
rect 50759 202961 50787 202989
rect 50821 202961 50849 202989
rect 50883 202961 50911 202989
rect 50697 194147 50725 194175
rect 50759 194147 50787 194175
rect 50821 194147 50849 194175
rect 50883 194147 50911 194175
rect 50697 194085 50725 194113
rect 50759 194085 50787 194113
rect 50821 194085 50849 194113
rect 50883 194085 50911 194113
rect 50697 194023 50725 194051
rect 50759 194023 50787 194051
rect 50821 194023 50849 194051
rect 50883 194023 50911 194051
rect 50697 193961 50725 193989
rect 50759 193961 50787 193989
rect 50821 193961 50849 193989
rect 50883 193961 50911 193989
rect 50697 185147 50725 185175
rect 50759 185147 50787 185175
rect 50821 185147 50849 185175
rect 50883 185147 50911 185175
rect 50697 185085 50725 185113
rect 50759 185085 50787 185113
rect 50821 185085 50849 185113
rect 50883 185085 50911 185113
rect 50697 185023 50725 185051
rect 50759 185023 50787 185051
rect 50821 185023 50849 185051
rect 50883 185023 50911 185051
rect 50697 184961 50725 184989
rect 50759 184961 50787 184989
rect 50821 184961 50849 184989
rect 50883 184961 50911 184989
rect 50697 176147 50725 176175
rect 50759 176147 50787 176175
rect 50821 176147 50849 176175
rect 50883 176147 50911 176175
rect 50697 176085 50725 176113
rect 50759 176085 50787 176113
rect 50821 176085 50849 176113
rect 50883 176085 50911 176113
rect 50697 176023 50725 176051
rect 50759 176023 50787 176051
rect 50821 176023 50849 176051
rect 50883 176023 50911 176051
rect 50697 175961 50725 175989
rect 50759 175961 50787 175989
rect 50821 175961 50849 175989
rect 50883 175961 50911 175989
rect 64197 298578 64225 298606
rect 64259 298578 64287 298606
rect 64321 298578 64349 298606
rect 64383 298578 64411 298606
rect 64197 298516 64225 298544
rect 64259 298516 64287 298544
rect 64321 298516 64349 298544
rect 64383 298516 64411 298544
rect 64197 298454 64225 298482
rect 64259 298454 64287 298482
rect 64321 298454 64349 298482
rect 64383 298454 64411 298482
rect 64197 298392 64225 298420
rect 64259 298392 64287 298420
rect 64321 298392 64349 298420
rect 64383 298392 64411 298420
rect 64197 290147 64225 290175
rect 64259 290147 64287 290175
rect 64321 290147 64349 290175
rect 64383 290147 64411 290175
rect 64197 290085 64225 290113
rect 64259 290085 64287 290113
rect 64321 290085 64349 290113
rect 64383 290085 64411 290113
rect 64197 290023 64225 290051
rect 64259 290023 64287 290051
rect 64321 290023 64349 290051
rect 64383 290023 64411 290051
rect 64197 289961 64225 289989
rect 64259 289961 64287 289989
rect 64321 289961 64349 289989
rect 64383 289961 64411 289989
rect 64197 281147 64225 281175
rect 64259 281147 64287 281175
rect 64321 281147 64349 281175
rect 64383 281147 64411 281175
rect 64197 281085 64225 281113
rect 64259 281085 64287 281113
rect 64321 281085 64349 281113
rect 64383 281085 64411 281113
rect 64197 281023 64225 281051
rect 64259 281023 64287 281051
rect 64321 281023 64349 281051
rect 64383 281023 64411 281051
rect 64197 280961 64225 280989
rect 64259 280961 64287 280989
rect 64321 280961 64349 280989
rect 64383 280961 64411 280989
rect 64197 272147 64225 272175
rect 64259 272147 64287 272175
rect 64321 272147 64349 272175
rect 64383 272147 64411 272175
rect 64197 272085 64225 272113
rect 64259 272085 64287 272113
rect 64321 272085 64349 272113
rect 64383 272085 64411 272113
rect 64197 272023 64225 272051
rect 64259 272023 64287 272051
rect 64321 272023 64349 272051
rect 64383 272023 64411 272051
rect 64197 271961 64225 271989
rect 64259 271961 64287 271989
rect 64321 271961 64349 271989
rect 64383 271961 64411 271989
rect 64197 263147 64225 263175
rect 64259 263147 64287 263175
rect 64321 263147 64349 263175
rect 64383 263147 64411 263175
rect 64197 263085 64225 263113
rect 64259 263085 64287 263113
rect 64321 263085 64349 263113
rect 64383 263085 64411 263113
rect 64197 263023 64225 263051
rect 64259 263023 64287 263051
rect 64321 263023 64349 263051
rect 64383 263023 64411 263051
rect 64197 262961 64225 262989
rect 64259 262961 64287 262989
rect 64321 262961 64349 262989
rect 64383 262961 64411 262989
rect 64197 254147 64225 254175
rect 64259 254147 64287 254175
rect 64321 254147 64349 254175
rect 64383 254147 64411 254175
rect 64197 254085 64225 254113
rect 64259 254085 64287 254113
rect 64321 254085 64349 254113
rect 64383 254085 64411 254113
rect 64197 254023 64225 254051
rect 64259 254023 64287 254051
rect 64321 254023 64349 254051
rect 64383 254023 64411 254051
rect 64197 253961 64225 253989
rect 64259 253961 64287 253989
rect 64321 253961 64349 253989
rect 64383 253961 64411 253989
rect 64197 245147 64225 245175
rect 64259 245147 64287 245175
rect 64321 245147 64349 245175
rect 64383 245147 64411 245175
rect 64197 245085 64225 245113
rect 64259 245085 64287 245113
rect 64321 245085 64349 245113
rect 64383 245085 64411 245113
rect 64197 245023 64225 245051
rect 64259 245023 64287 245051
rect 64321 245023 64349 245051
rect 64383 245023 64411 245051
rect 64197 244961 64225 244989
rect 64259 244961 64287 244989
rect 64321 244961 64349 244989
rect 64383 244961 64411 244989
rect 64197 236147 64225 236175
rect 64259 236147 64287 236175
rect 64321 236147 64349 236175
rect 64383 236147 64411 236175
rect 64197 236085 64225 236113
rect 64259 236085 64287 236113
rect 64321 236085 64349 236113
rect 64383 236085 64411 236113
rect 64197 236023 64225 236051
rect 64259 236023 64287 236051
rect 64321 236023 64349 236051
rect 64383 236023 64411 236051
rect 64197 235961 64225 235989
rect 64259 235961 64287 235989
rect 64321 235961 64349 235989
rect 64383 235961 64411 235989
rect 64197 227147 64225 227175
rect 64259 227147 64287 227175
rect 64321 227147 64349 227175
rect 64383 227147 64411 227175
rect 64197 227085 64225 227113
rect 64259 227085 64287 227113
rect 64321 227085 64349 227113
rect 64383 227085 64411 227113
rect 64197 227023 64225 227051
rect 64259 227023 64287 227051
rect 64321 227023 64349 227051
rect 64383 227023 64411 227051
rect 64197 226961 64225 226989
rect 64259 226961 64287 226989
rect 64321 226961 64349 226989
rect 64383 226961 64411 226989
rect 64197 218147 64225 218175
rect 64259 218147 64287 218175
rect 64321 218147 64349 218175
rect 64383 218147 64411 218175
rect 64197 218085 64225 218113
rect 64259 218085 64287 218113
rect 64321 218085 64349 218113
rect 64383 218085 64411 218113
rect 64197 218023 64225 218051
rect 64259 218023 64287 218051
rect 64321 218023 64349 218051
rect 64383 218023 64411 218051
rect 64197 217961 64225 217989
rect 64259 217961 64287 217989
rect 64321 217961 64349 217989
rect 64383 217961 64411 217989
rect 64197 209147 64225 209175
rect 64259 209147 64287 209175
rect 64321 209147 64349 209175
rect 64383 209147 64411 209175
rect 64197 209085 64225 209113
rect 64259 209085 64287 209113
rect 64321 209085 64349 209113
rect 64383 209085 64411 209113
rect 64197 209023 64225 209051
rect 64259 209023 64287 209051
rect 64321 209023 64349 209051
rect 64383 209023 64411 209051
rect 64197 208961 64225 208989
rect 64259 208961 64287 208989
rect 64321 208961 64349 208989
rect 64383 208961 64411 208989
rect 64197 200147 64225 200175
rect 64259 200147 64287 200175
rect 64321 200147 64349 200175
rect 64383 200147 64411 200175
rect 64197 200085 64225 200113
rect 64259 200085 64287 200113
rect 64321 200085 64349 200113
rect 64383 200085 64411 200113
rect 64197 200023 64225 200051
rect 64259 200023 64287 200051
rect 64321 200023 64349 200051
rect 64383 200023 64411 200051
rect 64197 199961 64225 199989
rect 64259 199961 64287 199989
rect 64321 199961 64349 199989
rect 64383 199961 64411 199989
rect 64197 191147 64225 191175
rect 64259 191147 64287 191175
rect 64321 191147 64349 191175
rect 64383 191147 64411 191175
rect 64197 191085 64225 191113
rect 64259 191085 64287 191113
rect 64321 191085 64349 191113
rect 64383 191085 64411 191113
rect 64197 191023 64225 191051
rect 64259 191023 64287 191051
rect 64321 191023 64349 191051
rect 64383 191023 64411 191051
rect 64197 190961 64225 190989
rect 64259 190961 64287 190989
rect 64321 190961 64349 190989
rect 64383 190961 64411 190989
rect 64197 182147 64225 182175
rect 64259 182147 64287 182175
rect 64321 182147 64349 182175
rect 64383 182147 64411 182175
rect 64197 182085 64225 182113
rect 64259 182085 64287 182113
rect 64321 182085 64349 182113
rect 64383 182085 64411 182113
rect 64197 182023 64225 182051
rect 64259 182023 64287 182051
rect 64321 182023 64349 182051
rect 64383 182023 64411 182051
rect 64197 181961 64225 181989
rect 64259 181961 64287 181989
rect 64321 181961 64349 181989
rect 64383 181961 64411 181989
rect 54339 173147 54367 173175
rect 54401 173147 54429 173175
rect 54339 173085 54367 173113
rect 54401 173085 54429 173113
rect 54339 173023 54367 173051
rect 54401 173023 54429 173051
rect 54339 172961 54367 172989
rect 54401 172961 54429 172989
rect 64197 173147 64225 173175
rect 64259 173147 64287 173175
rect 64321 173147 64349 173175
rect 64383 173147 64411 173175
rect 64197 173085 64225 173113
rect 64259 173085 64287 173113
rect 64321 173085 64349 173113
rect 64383 173085 64411 173113
rect 64197 173023 64225 173051
rect 64259 173023 64287 173051
rect 64321 173023 64349 173051
rect 64383 173023 64411 173051
rect 64197 172961 64225 172989
rect 64259 172961 64287 172989
rect 64321 172961 64349 172989
rect 64383 172961 64411 172989
rect 50697 167147 50725 167175
rect 50759 167147 50787 167175
rect 50821 167147 50849 167175
rect 50883 167147 50911 167175
rect 50697 167085 50725 167113
rect 50759 167085 50787 167113
rect 50821 167085 50849 167113
rect 50883 167085 50911 167113
rect 50697 167023 50725 167051
rect 50759 167023 50787 167051
rect 50821 167023 50849 167051
rect 50883 167023 50911 167051
rect 50697 166961 50725 166989
rect 50759 166961 50787 166989
rect 50821 166961 50849 166989
rect 50883 166961 50911 166989
rect 62019 167147 62047 167175
rect 62081 167147 62109 167175
rect 62019 167085 62047 167113
rect 62081 167085 62109 167113
rect 62019 167023 62047 167051
rect 62081 167023 62109 167051
rect 62019 166961 62047 166989
rect 62081 166961 62109 166989
rect 54339 164147 54367 164175
rect 54401 164147 54429 164175
rect 54339 164085 54367 164113
rect 54401 164085 54429 164113
rect 54339 164023 54367 164051
rect 54401 164023 54429 164051
rect 54339 163961 54367 163989
rect 54401 163961 54429 163989
rect 64197 164147 64225 164175
rect 64259 164147 64287 164175
rect 64321 164147 64349 164175
rect 64383 164147 64411 164175
rect 64197 164085 64225 164113
rect 64259 164085 64287 164113
rect 64321 164085 64349 164113
rect 64383 164085 64411 164113
rect 64197 164023 64225 164051
rect 64259 164023 64287 164051
rect 64321 164023 64349 164051
rect 64383 164023 64411 164051
rect 64197 163961 64225 163989
rect 64259 163961 64287 163989
rect 64321 163961 64349 163989
rect 64383 163961 64411 163989
rect 50697 158147 50725 158175
rect 50759 158147 50787 158175
rect 50821 158147 50849 158175
rect 50883 158147 50911 158175
rect 50697 158085 50725 158113
rect 50759 158085 50787 158113
rect 50821 158085 50849 158113
rect 50883 158085 50911 158113
rect 50697 158023 50725 158051
rect 50759 158023 50787 158051
rect 50821 158023 50849 158051
rect 50883 158023 50911 158051
rect 50697 157961 50725 157989
rect 50759 157961 50787 157989
rect 50821 157961 50849 157989
rect 50883 157961 50911 157989
rect 62019 158147 62047 158175
rect 62081 158147 62109 158175
rect 62019 158085 62047 158113
rect 62081 158085 62109 158113
rect 62019 158023 62047 158051
rect 62081 158023 62109 158051
rect 62019 157961 62047 157989
rect 62081 157961 62109 157989
rect 54339 155147 54367 155175
rect 54401 155147 54429 155175
rect 54339 155085 54367 155113
rect 54401 155085 54429 155113
rect 54339 155023 54367 155051
rect 54401 155023 54429 155051
rect 54339 154961 54367 154989
rect 54401 154961 54429 154989
rect 64197 155147 64225 155175
rect 64259 155147 64287 155175
rect 64321 155147 64349 155175
rect 64383 155147 64411 155175
rect 64197 155085 64225 155113
rect 64259 155085 64287 155113
rect 64321 155085 64349 155113
rect 64383 155085 64411 155113
rect 64197 155023 64225 155051
rect 64259 155023 64287 155051
rect 64321 155023 64349 155051
rect 64383 155023 64411 155051
rect 64197 154961 64225 154989
rect 64259 154961 64287 154989
rect 64321 154961 64349 154989
rect 64383 154961 64411 154989
rect 50697 149147 50725 149175
rect 50759 149147 50787 149175
rect 50821 149147 50849 149175
rect 50883 149147 50911 149175
rect 50697 149085 50725 149113
rect 50759 149085 50787 149113
rect 50821 149085 50849 149113
rect 50883 149085 50911 149113
rect 50697 149023 50725 149051
rect 50759 149023 50787 149051
rect 50821 149023 50849 149051
rect 50883 149023 50911 149051
rect 50697 148961 50725 148989
rect 50759 148961 50787 148989
rect 50821 148961 50849 148989
rect 50883 148961 50911 148989
rect 62019 149147 62047 149175
rect 62081 149147 62109 149175
rect 62019 149085 62047 149113
rect 62081 149085 62109 149113
rect 62019 149023 62047 149051
rect 62081 149023 62109 149051
rect 62019 148961 62047 148989
rect 62081 148961 62109 148989
rect 54339 146147 54367 146175
rect 54401 146147 54429 146175
rect 54339 146085 54367 146113
rect 54401 146085 54429 146113
rect 54339 146023 54367 146051
rect 54401 146023 54429 146051
rect 54339 145961 54367 145989
rect 54401 145961 54429 145989
rect 64197 146147 64225 146175
rect 64259 146147 64287 146175
rect 64321 146147 64349 146175
rect 64383 146147 64411 146175
rect 64197 146085 64225 146113
rect 64259 146085 64287 146113
rect 64321 146085 64349 146113
rect 64383 146085 64411 146113
rect 64197 146023 64225 146051
rect 64259 146023 64287 146051
rect 64321 146023 64349 146051
rect 64383 146023 64411 146051
rect 64197 145961 64225 145989
rect 64259 145961 64287 145989
rect 64321 145961 64349 145989
rect 64383 145961 64411 145989
rect 50697 140147 50725 140175
rect 50759 140147 50787 140175
rect 50821 140147 50849 140175
rect 50883 140147 50911 140175
rect 50697 140085 50725 140113
rect 50759 140085 50787 140113
rect 50821 140085 50849 140113
rect 50883 140085 50911 140113
rect 50697 140023 50725 140051
rect 50759 140023 50787 140051
rect 50821 140023 50849 140051
rect 50883 140023 50911 140051
rect 50697 139961 50725 139989
rect 50759 139961 50787 139989
rect 50821 139961 50849 139989
rect 50883 139961 50911 139989
rect 62019 140147 62047 140175
rect 62081 140147 62109 140175
rect 62019 140085 62047 140113
rect 62081 140085 62109 140113
rect 62019 140023 62047 140051
rect 62081 140023 62109 140051
rect 62019 139961 62047 139989
rect 62081 139961 62109 139989
rect 54339 137147 54367 137175
rect 54401 137147 54429 137175
rect 54339 137085 54367 137113
rect 54401 137085 54429 137113
rect 54339 137023 54367 137051
rect 54401 137023 54429 137051
rect 54339 136961 54367 136989
rect 54401 136961 54429 136989
rect 64197 137147 64225 137175
rect 64259 137147 64287 137175
rect 64321 137147 64349 137175
rect 64383 137147 64411 137175
rect 64197 137085 64225 137113
rect 64259 137085 64287 137113
rect 64321 137085 64349 137113
rect 64383 137085 64411 137113
rect 64197 137023 64225 137051
rect 64259 137023 64287 137051
rect 64321 137023 64349 137051
rect 64383 137023 64411 137051
rect 64197 136961 64225 136989
rect 64259 136961 64287 136989
rect 64321 136961 64349 136989
rect 64383 136961 64411 136989
rect 50697 131147 50725 131175
rect 50759 131147 50787 131175
rect 50821 131147 50849 131175
rect 50883 131147 50911 131175
rect 50697 131085 50725 131113
rect 50759 131085 50787 131113
rect 50821 131085 50849 131113
rect 50883 131085 50911 131113
rect 50697 131023 50725 131051
rect 50759 131023 50787 131051
rect 50821 131023 50849 131051
rect 50883 131023 50911 131051
rect 50697 130961 50725 130989
rect 50759 130961 50787 130989
rect 50821 130961 50849 130989
rect 50883 130961 50911 130989
rect 62019 131147 62047 131175
rect 62081 131147 62109 131175
rect 62019 131085 62047 131113
rect 62081 131085 62109 131113
rect 62019 131023 62047 131051
rect 62081 131023 62109 131051
rect 62019 130961 62047 130989
rect 62081 130961 62109 130989
rect 54339 128147 54367 128175
rect 54401 128147 54429 128175
rect 54339 128085 54367 128113
rect 54401 128085 54429 128113
rect 54339 128023 54367 128051
rect 54401 128023 54429 128051
rect 54339 127961 54367 127989
rect 54401 127961 54429 127989
rect 64197 128147 64225 128175
rect 64259 128147 64287 128175
rect 64321 128147 64349 128175
rect 64383 128147 64411 128175
rect 64197 128085 64225 128113
rect 64259 128085 64287 128113
rect 64321 128085 64349 128113
rect 64383 128085 64411 128113
rect 64197 128023 64225 128051
rect 64259 128023 64287 128051
rect 64321 128023 64349 128051
rect 64383 128023 64411 128051
rect 64197 127961 64225 127989
rect 64259 127961 64287 127989
rect 64321 127961 64349 127989
rect 64383 127961 64411 127989
rect 50697 122147 50725 122175
rect 50759 122147 50787 122175
rect 50821 122147 50849 122175
rect 50883 122147 50911 122175
rect 50697 122085 50725 122113
rect 50759 122085 50787 122113
rect 50821 122085 50849 122113
rect 50883 122085 50911 122113
rect 50697 122023 50725 122051
rect 50759 122023 50787 122051
rect 50821 122023 50849 122051
rect 50883 122023 50911 122051
rect 50697 121961 50725 121989
rect 50759 121961 50787 121989
rect 50821 121961 50849 121989
rect 50883 121961 50911 121989
rect 62019 122147 62047 122175
rect 62081 122147 62109 122175
rect 62019 122085 62047 122113
rect 62081 122085 62109 122113
rect 62019 122023 62047 122051
rect 62081 122023 62109 122051
rect 62019 121961 62047 121989
rect 62081 121961 62109 121989
rect 54339 119147 54367 119175
rect 54401 119147 54429 119175
rect 54339 119085 54367 119113
rect 54401 119085 54429 119113
rect 54339 119023 54367 119051
rect 54401 119023 54429 119051
rect 54339 118961 54367 118989
rect 54401 118961 54429 118989
rect 64197 119147 64225 119175
rect 64259 119147 64287 119175
rect 64321 119147 64349 119175
rect 64383 119147 64411 119175
rect 64197 119085 64225 119113
rect 64259 119085 64287 119113
rect 64321 119085 64349 119113
rect 64383 119085 64411 119113
rect 64197 119023 64225 119051
rect 64259 119023 64287 119051
rect 64321 119023 64349 119051
rect 64383 119023 64411 119051
rect 64197 118961 64225 118989
rect 64259 118961 64287 118989
rect 64321 118961 64349 118989
rect 64383 118961 64411 118989
rect 50697 113147 50725 113175
rect 50759 113147 50787 113175
rect 50821 113147 50849 113175
rect 50883 113147 50911 113175
rect 50697 113085 50725 113113
rect 50759 113085 50787 113113
rect 50821 113085 50849 113113
rect 50883 113085 50911 113113
rect 50697 113023 50725 113051
rect 50759 113023 50787 113051
rect 50821 113023 50849 113051
rect 50883 113023 50911 113051
rect 50697 112961 50725 112989
rect 50759 112961 50787 112989
rect 50821 112961 50849 112989
rect 50883 112961 50911 112989
rect 62019 113147 62047 113175
rect 62081 113147 62109 113175
rect 62019 113085 62047 113113
rect 62081 113085 62109 113113
rect 62019 113023 62047 113051
rect 62081 113023 62109 113051
rect 62019 112961 62047 112989
rect 62081 112961 62109 112989
rect 54339 110147 54367 110175
rect 54401 110147 54429 110175
rect 54339 110085 54367 110113
rect 54401 110085 54429 110113
rect 54339 110023 54367 110051
rect 54401 110023 54429 110051
rect 54339 109961 54367 109989
rect 54401 109961 54429 109989
rect 64197 110147 64225 110175
rect 64259 110147 64287 110175
rect 64321 110147 64349 110175
rect 64383 110147 64411 110175
rect 64197 110085 64225 110113
rect 64259 110085 64287 110113
rect 64321 110085 64349 110113
rect 64383 110085 64411 110113
rect 64197 110023 64225 110051
rect 64259 110023 64287 110051
rect 64321 110023 64349 110051
rect 64383 110023 64411 110051
rect 64197 109961 64225 109989
rect 64259 109961 64287 109989
rect 64321 109961 64349 109989
rect 64383 109961 64411 109989
rect 50697 104147 50725 104175
rect 50759 104147 50787 104175
rect 50821 104147 50849 104175
rect 50883 104147 50911 104175
rect 50697 104085 50725 104113
rect 50759 104085 50787 104113
rect 50821 104085 50849 104113
rect 50883 104085 50911 104113
rect 50697 104023 50725 104051
rect 50759 104023 50787 104051
rect 50821 104023 50849 104051
rect 50883 104023 50911 104051
rect 50697 103961 50725 103989
rect 50759 103961 50787 103989
rect 50821 103961 50849 103989
rect 50883 103961 50911 103989
rect 62019 104147 62047 104175
rect 62081 104147 62109 104175
rect 62019 104085 62047 104113
rect 62081 104085 62109 104113
rect 62019 104023 62047 104051
rect 62081 104023 62109 104051
rect 62019 103961 62047 103989
rect 62081 103961 62109 103989
rect 54339 101147 54367 101175
rect 54401 101147 54429 101175
rect 54339 101085 54367 101113
rect 54401 101085 54429 101113
rect 54339 101023 54367 101051
rect 54401 101023 54429 101051
rect 54339 100961 54367 100989
rect 54401 100961 54429 100989
rect 64197 101147 64225 101175
rect 64259 101147 64287 101175
rect 64321 101147 64349 101175
rect 64383 101147 64411 101175
rect 64197 101085 64225 101113
rect 64259 101085 64287 101113
rect 64321 101085 64349 101113
rect 64383 101085 64411 101113
rect 64197 101023 64225 101051
rect 64259 101023 64287 101051
rect 64321 101023 64349 101051
rect 64383 101023 64411 101051
rect 64197 100961 64225 100989
rect 64259 100961 64287 100989
rect 64321 100961 64349 100989
rect 64383 100961 64411 100989
rect 50697 95147 50725 95175
rect 50759 95147 50787 95175
rect 50821 95147 50849 95175
rect 50883 95147 50911 95175
rect 50697 95085 50725 95113
rect 50759 95085 50787 95113
rect 50821 95085 50849 95113
rect 50883 95085 50911 95113
rect 50697 95023 50725 95051
rect 50759 95023 50787 95051
rect 50821 95023 50849 95051
rect 50883 95023 50911 95051
rect 50697 94961 50725 94989
rect 50759 94961 50787 94989
rect 50821 94961 50849 94989
rect 50883 94961 50911 94989
rect 62019 95147 62047 95175
rect 62081 95147 62109 95175
rect 62019 95085 62047 95113
rect 62081 95085 62109 95113
rect 62019 95023 62047 95051
rect 62081 95023 62109 95051
rect 62019 94961 62047 94989
rect 62081 94961 62109 94989
rect 54339 92147 54367 92175
rect 54401 92147 54429 92175
rect 54339 92085 54367 92113
rect 54401 92085 54429 92113
rect 54339 92023 54367 92051
rect 54401 92023 54429 92051
rect 54339 91961 54367 91989
rect 54401 91961 54429 91989
rect 64197 92147 64225 92175
rect 64259 92147 64287 92175
rect 64321 92147 64349 92175
rect 64383 92147 64411 92175
rect 64197 92085 64225 92113
rect 64259 92085 64287 92113
rect 64321 92085 64349 92113
rect 64383 92085 64411 92113
rect 64197 92023 64225 92051
rect 64259 92023 64287 92051
rect 64321 92023 64349 92051
rect 64383 92023 64411 92051
rect 64197 91961 64225 91989
rect 64259 91961 64287 91989
rect 64321 91961 64349 91989
rect 64383 91961 64411 91989
rect 50697 86147 50725 86175
rect 50759 86147 50787 86175
rect 50821 86147 50849 86175
rect 50883 86147 50911 86175
rect 50697 86085 50725 86113
rect 50759 86085 50787 86113
rect 50821 86085 50849 86113
rect 50883 86085 50911 86113
rect 50697 86023 50725 86051
rect 50759 86023 50787 86051
rect 50821 86023 50849 86051
rect 50883 86023 50911 86051
rect 50697 85961 50725 85989
rect 50759 85961 50787 85989
rect 50821 85961 50849 85989
rect 50883 85961 50911 85989
rect 62019 86147 62047 86175
rect 62081 86147 62109 86175
rect 62019 86085 62047 86113
rect 62081 86085 62109 86113
rect 62019 86023 62047 86051
rect 62081 86023 62109 86051
rect 62019 85961 62047 85989
rect 62081 85961 62109 85989
rect 54339 83147 54367 83175
rect 54401 83147 54429 83175
rect 54339 83085 54367 83113
rect 54401 83085 54429 83113
rect 54339 83023 54367 83051
rect 54401 83023 54429 83051
rect 54339 82961 54367 82989
rect 54401 82961 54429 82989
rect 64197 83147 64225 83175
rect 64259 83147 64287 83175
rect 64321 83147 64349 83175
rect 64383 83147 64411 83175
rect 64197 83085 64225 83113
rect 64259 83085 64287 83113
rect 64321 83085 64349 83113
rect 64383 83085 64411 83113
rect 64197 83023 64225 83051
rect 64259 83023 64287 83051
rect 64321 83023 64349 83051
rect 64383 83023 64411 83051
rect 64197 82961 64225 82989
rect 64259 82961 64287 82989
rect 64321 82961 64349 82989
rect 64383 82961 64411 82989
rect 50697 77147 50725 77175
rect 50759 77147 50787 77175
rect 50821 77147 50849 77175
rect 50883 77147 50911 77175
rect 50697 77085 50725 77113
rect 50759 77085 50787 77113
rect 50821 77085 50849 77113
rect 50883 77085 50911 77113
rect 50697 77023 50725 77051
rect 50759 77023 50787 77051
rect 50821 77023 50849 77051
rect 50883 77023 50911 77051
rect 50697 76961 50725 76989
rect 50759 76961 50787 76989
rect 50821 76961 50849 76989
rect 50883 76961 50911 76989
rect 62019 77147 62047 77175
rect 62081 77147 62109 77175
rect 62019 77085 62047 77113
rect 62081 77085 62109 77113
rect 62019 77023 62047 77051
rect 62081 77023 62109 77051
rect 62019 76961 62047 76989
rect 62081 76961 62109 76989
rect 54339 74147 54367 74175
rect 54401 74147 54429 74175
rect 54339 74085 54367 74113
rect 54401 74085 54429 74113
rect 54339 74023 54367 74051
rect 54401 74023 54429 74051
rect 54339 73961 54367 73989
rect 54401 73961 54429 73989
rect 64197 74147 64225 74175
rect 64259 74147 64287 74175
rect 64321 74147 64349 74175
rect 64383 74147 64411 74175
rect 64197 74085 64225 74113
rect 64259 74085 64287 74113
rect 64321 74085 64349 74113
rect 64383 74085 64411 74113
rect 64197 74023 64225 74051
rect 64259 74023 64287 74051
rect 64321 74023 64349 74051
rect 64383 74023 64411 74051
rect 64197 73961 64225 73989
rect 64259 73961 64287 73989
rect 64321 73961 64349 73989
rect 64383 73961 64411 73989
rect 50697 68147 50725 68175
rect 50759 68147 50787 68175
rect 50821 68147 50849 68175
rect 50883 68147 50911 68175
rect 50697 68085 50725 68113
rect 50759 68085 50787 68113
rect 50821 68085 50849 68113
rect 50883 68085 50911 68113
rect 50697 68023 50725 68051
rect 50759 68023 50787 68051
rect 50821 68023 50849 68051
rect 50883 68023 50911 68051
rect 50697 67961 50725 67989
rect 50759 67961 50787 67989
rect 50821 67961 50849 67989
rect 50883 67961 50911 67989
rect 62019 68147 62047 68175
rect 62081 68147 62109 68175
rect 62019 68085 62047 68113
rect 62081 68085 62109 68113
rect 62019 68023 62047 68051
rect 62081 68023 62109 68051
rect 62019 67961 62047 67989
rect 62081 67961 62109 67989
rect 54339 65147 54367 65175
rect 54401 65147 54429 65175
rect 54339 65085 54367 65113
rect 54401 65085 54429 65113
rect 54339 65023 54367 65051
rect 54401 65023 54429 65051
rect 54339 64961 54367 64989
rect 54401 64961 54429 64989
rect 64197 65147 64225 65175
rect 64259 65147 64287 65175
rect 64321 65147 64349 65175
rect 64383 65147 64411 65175
rect 64197 65085 64225 65113
rect 64259 65085 64287 65113
rect 64321 65085 64349 65113
rect 64383 65085 64411 65113
rect 64197 65023 64225 65051
rect 64259 65023 64287 65051
rect 64321 65023 64349 65051
rect 64383 65023 64411 65051
rect 64197 64961 64225 64989
rect 64259 64961 64287 64989
rect 64321 64961 64349 64989
rect 64383 64961 64411 64989
rect 50697 59147 50725 59175
rect 50759 59147 50787 59175
rect 50821 59147 50849 59175
rect 50883 59147 50911 59175
rect 50697 59085 50725 59113
rect 50759 59085 50787 59113
rect 50821 59085 50849 59113
rect 50883 59085 50911 59113
rect 50697 59023 50725 59051
rect 50759 59023 50787 59051
rect 50821 59023 50849 59051
rect 50883 59023 50911 59051
rect 50697 58961 50725 58989
rect 50759 58961 50787 58989
rect 50821 58961 50849 58989
rect 50883 58961 50911 58989
rect 62019 59147 62047 59175
rect 62081 59147 62109 59175
rect 62019 59085 62047 59113
rect 62081 59085 62109 59113
rect 62019 59023 62047 59051
rect 62081 59023 62109 59051
rect 62019 58961 62047 58989
rect 62081 58961 62109 58989
rect 54339 56147 54367 56175
rect 54401 56147 54429 56175
rect 54339 56085 54367 56113
rect 54401 56085 54429 56113
rect 54339 56023 54367 56051
rect 54401 56023 54429 56051
rect 54339 55961 54367 55989
rect 54401 55961 54429 55989
rect 64197 56147 64225 56175
rect 64259 56147 64287 56175
rect 64321 56147 64349 56175
rect 64383 56147 64411 56175
rect 64197 56085 64225 56113
rect 64259 56085 64287 56113
rect 64321 56085 64349 56113
rect 64383 56085 64411 56113
rect 64197 56023 64225 56051
rect 64259 56023 64287 56051
rect 64321 56023 64349 56051
rect 64383 56023 64411 56051
rect 64197 55961 64225 55989
rect 64259 55961 64287 55989
rect 64321 55961 64349 55989
rect 64383 55961 64411 55989
rect 50697 50147 50725 50175
rect 50759 50147 50787 50175
rect 50821 50147 50849 50175
rect 50883 50147 50911 50175
rect 50697 50085 50725 50113
rect 50759 50085 50787 50113
rect 50821 50085 50849 50113
rect 50883 50085 50911 50113
rect 50697 50023 50725 50051
rect 50759 50023 50787 50051
rect 50821 50023 50849 50051
rect 50883 50023 50911 50051
rect 50697 49961 50725 49989
rect 50759 49961 50787 49989
rect 50821 49961 50849 49989
rect 50883 49961 50911 49989
rect 62019 50147 62047 50175
rect 62081 50147 62109 50175
rect 62019 50085 62047 50113
rect 62081 50085 62109 50113
rect 62019 50023 62047 50051
rect 62081 50023 62109 50051
rect 62019 49961 62047 49989
rect 62081 49961 62109 49989
rect 54339 47147 54367 47175
rect 54401 47147 54429 47175
rect 54339 47085 54367 47113
rect 54401 47085 54429 47113
rect 54339 47023 54367 47051
rect 54401 47023 54429 47051
rect 54339 46961 54367 46989
rect 54401 46961 54429 46989
rect 64197 47147 64225 47175
rect 64259 47147 64287 47175
rect 64321 47147 64349 47175
rect 64383 47147 64411 47175
rect 64197 47085 64225 47113
rect 64259 47085 64287 47113
rect 64321 47085 64349 47113
rect 64383 47085 64411 47113
rect 64197 47023 64225 47051
rect 64259 47023 64287 47051
rect 64321 47023 64349 47051
rect 64383 47023 64411 47051
rect 64197 46961 64225 46989
rect 64259 46961 64287 46989
rect 64321 46961 64349 46989
rect 64383 46961 64411 46989
rect 50697 41147 50725 41175
rect 50759 41147 50787 41175
rect 50821 41147 50849 41175
rect 50883 41147 50911 41175
rect 50697 41085 50725 41113
rect 50759 41085 50787 41113
rect 50821 41085 50849 41113
rect 50883 41085 50911 41113
rect 50697 41023 50725 41051
rect 50759 41023 50787 41051
rect 50821 41023 50849 41051
rect 50883 41023 50911 41051
rect 50697 40961 50725 40989
rect 50759 40961 50787 40989
rect 50821 40961 50849 40989
rect 50883 40961 50911 40989
rect 62019 41147 62047 41175
rect 62081 41147 62109 41175
rect 62019 41085 62047 41113
rect 62081 41085 62109 41113
rect 62019 41023 62047 41051
rect 62081 41023 62109 41051
rect 62019 40961 62047 40989
rect 62081 40961 62109 40989
rect 54339 38147 54367 38175
rect 54401 38147 54429 38175
rect 54339 38085 54367 38113
rect 54401 38085 54429 38113
rect 54339 38023 54367 38051
rect 54401 38023 54429 38051
rect 54339 37961 54367 37989
rect 54401 37961 54429 37989
rect 64197 38147 64225 38175
rect 64259 38147 64287 38175
rect 64321 38147 64349 38175
rect 64383 38147 64411 38175
rect 64197 38085 64225 38113
rect 64259 38085 64287 38113
rect 64321 38085 64349 38113
rect 64383 38085 64411 38113
rect 64197 38023 64225 38051
rect 64259 38023 64287 38051
rect 64321 38023 64349 38051
rect 64383 38023 64411 38051
rect 64197 37961 64225 37989
rect 64259 37961 64287 37989
rect 64321 37961 64349 37989
rect 64383 37961 64411 37989
rect 50697 32147 50725 32175
rect 50759 32147 50787 32175
rect 50821 32147 50849 32175
rect 50883 32147 50911 32175
rect 50697 32085 50725 32113
rect 50759 32085 50787 32113
rect 50821 32085 50849 32113
rect 50883 32085 50911 32113
rect 50697 32023 50725 32051
rect 50759 32023 50787 32051
rect 50821 32023 50849 32051
rect 50883 32023 50911 32051
rect 50697 31961 50725 31989
rect 50759 31961 50787 31989
rect 50821 31961 50849 31989
rect 50883 31961 50911 31989
rect 62019 32147 62047 32175
rect 62081 32147 62109 32175
rect 62019 32085 62047 32113
rect 62081 32085 62109 32113
rect 62019 32023 62047 32051
rect 62081 32023 62109 32051
rect 62019 31961 62047 31989
rect 62081 31961 62109 31989
rect 54339 29147 54367 29175
rect 54401 29147 54429 29175
rect 54339 29085 54367 29113
rect 54401 29085 54429 29113
rect 54339 29023 54367 29051
rect 54401 29023 54429 29051
rect 54339 28961 54367 28989
rect 54401 28961 54429 28989
rect 64197 29147 64225 29175
rect 64259 29147 64287 29175
rect 64321 29147 64349 29175
rect 64383 29147 64411 29175
rect 64197 29085 64225 29113
rect 64259 29085 64287 29113
rect 64321 29085 64349 29113
rect 64383 29085 64411 29113
rect 64197 29023 64225 29051
rect 64259 29023 64287 29051
rect 64321 29023 64349 29051
rect 64383 29023 64411 29051
rect 64197 28961 64225 28989
rect 64259 28961 64287 28989
rect 64321 28961 64349 28989
rect 64383 28961 64411 28989
rect 50697 23147 50725 23175
rect 50759 23147 50787 23175
rect 50821 23147 50849 23175
rect 50883 23147 50911 23175
rect 50697 23085 50725 23113
rect 50759 23085 50787 23113
rect 50821 23085 50849 23113
rect 50883 23085 50911 23113
rect 50697 23023 50725 23051
rect 50759 23023 50787 23051
rect 50821 23023 50849 23051
rect 50883 23023 50911 23051
rect 50697 22961 50725 22989
rect 50759 22961 50787 22989
rect 50821 22961 50849 22989
rect 50883 22961 50911 22989
rect 62019 23147 62047 23175
rect 62081 23147 62109 23175
rect 62019 23085 62047 23113
rect 62081 23085 62109 23113
rect 62019 23023 62047 23051
rect 62081 23023 62109 23051
rect 62019 22961 62047 22989
rect 62081 22961 62109 22989
rect 54339 20147 54367 20175
rect 54401 20147 54429 20175
rect 54339 20085 54367 20113
rect 54401 20085 54429 20113
rect 54339 20023 54367 20051
rect 54401 20023 54429 20051
rect 54339 19961 54367 19989
rect 54401 19961 54429 19989
rect 64197 20147 64225 20175
rect 64259 20147 64287 20175
rect 64321 20147 64349 20175
rect 64383 20147 64411 20175
rect 64197 20085 64225 20113
rect 64259 20085 64287 20113
rect 64321 20085 64349 20113
rect 64383 20085 64411 20113
rect 64197 20023 64225 20051
rect 64259 20023 64287 20051
rect 64321 20023 64349 20051
rect 64383 20023 64411 20051
rect 64197 19961 64225 19989
rect 64259 19961 64287 19989
rect 64321 19961 64349 19989
rect 64383 19961 64411 19989
rect 50697 14147 50725 14175
rect 50759 14147 50787 14175
rect 50821 14147 50849 14175
rect 50883 14147 50911 14175
rect 50697 14085 50725 14113
rect 50759 14085 50787 14113
rect 50821 14085 50849 14113
rect 50883 14085 50911 14113
rect 50697 14023 50725 14051
rect 50759 14023 50787 14051
rect 50821 14023 50849 14051
rect 50883 14023 50911 14051
rect 50697 13961 50725 13989
rect 50759 13961 50787 13989
rect 50821 13961 50849 13989
rect 50883 13961 50911 13989
rect 62019 14147 62047 14175
rect 62081 14147 62109 14175
rect 62019 14085 62047 14113
rect 62081 14085 62109 14113
rect 62019 14023 62047 14051
rect 62081 14023 62109 14051
rect 62019 13961 62047 13989
rect 62081 13961 62109 13989
rect 54339 11147 54367 11175
rect 54401 11147 54429 11175
rect 54339 11085 54367 11113
rect 54401 11085 54429 11113
rect 54339 11023 54367 11051
rect 54401 11023 54429 11051
rect 54339 10961 54367 10989
rect 54401 10961 54429 10989
rect 64197 11147 64225 11175
rect 64259 11147 64287 11175
rect 64321 11147 64349 11175
rect 64383 11147 64411 11175
rect 64197 11085 64225 11113
rect 64259 11085 64287 11113
rect 64321 11085 64349 11113
rect 64383 11085 64411 11113
rect 64197 11023 64225 11051
rect 64259 11023 64287 11051
rect 64321 11023 64349 11051
rect 64383 11023 64411 11051
rect 64197 10961 64225 10989
rect 64259 10961 64287 10989
rect 64321 10961 64349 10989
rect 64383 10961 64411 10989
rect 50697 5147 50725 5175
rect 50759 5147 50787 5175
rect 50821 5147 50849 5175
rect 50883 5147 50911 5175
rect 50697 5085 50725 5113
rect 50759 5085 50787 5113
rect 50821 5085 50849 5113
rect 50883 5085 50911 5113
rect 50697 5023 50725 5051
rect 50759 5023 50787 5051
rect 50821 5023 50849 5051
rect 50883 5023 50911 5051
rect 50697 4961 50725 4989
rect 50759 4961 50787 4989
rect 50821 4961 50849 4989
rect 50883 4961 50911 4989
rect 62019 5147 62047 5175
rect 62081 5147 62109 5175
rect 62019 5085 62047 5113
rect 62081 5085 62109 5113
rect 62019 5023 62047 5051
rect 62081 5023 62109 5051
rect 62019 4961 62047 4989
rect 62081 4961 62109 4989
rect 50697 -588 50725 -560
rect 50759 -588 50787 -560
rect 50821 -588 50849 -560
rect 50883 -588 50911 -560
rect 50697 -650 50725 -622
rect 50759 -650 50787 -622
rect 50821 -650 50849 -622
rect 50883 -650 50911 -622
rect 50697 -712 50725 -684
rect 50759 -712 50787 -684
rect 50821 -712 50849 -684
rect 50883 -712 50911 -684
rect 50697 -774 50725 -746
rect 50759 -774 50787 -746
rect 50821 -774 50849 -746
rect 50883 -774 50911 -746
rect 64197 2147 64225 2175
rect 64259 2147 64287 2175
rect 64321 2147 64349 2175
rect 64383 2147 64411 2175
rect 64197 2085 64225 2113
rect 64259 2085 64287 2113
rect 64321 2085 64349 2113
rect 64383 2085 64411 2113
rect 64197 2023 64225 2051
rect 64259 2023 64287 2051
rect 64321 2023 64349 2051
rect 64383 2023 64411 2051
rect 64197 1961 64225 1989
rect 64259 1961 64287 1989
rect 64321 1961 64349 1989
rect 64383 1961 64411 1989
rect 64197 -108 64225 -80
rect 64259 -108 64287 -80
rect 64321 -108 64349 -80
rect 64383 -108 64411 -80
rect 64197 -170 64225 -142
rect 64259 -170 64287 -142
rect 64321 -170 64349 -142
rect 64383 -170 64411 -142
rect 64197 -232 64225 -204
rect 64259 -232 64287 -204
rect 64321 -232 64349 -204
rect 64383 -232 64411 -204
rect 64197 -294 64225 -266
rect 64259 -294 64287 -266
rect 64321 -294 64349 -266
rect 64383 -294 64411 -266
rect 66057 299058 66085 299086
rect 66119 299058 66147 299086
rect 66181 299058 66209 299086
rect 66243 299058 66271 299086
rect 66057 298996 66085 299024
rect 66119 298996 66147 299024
rect 66181 298996 66209 299024
rect 66243 298996 66271 299024
rect 66057 298934 66085 298962
rect 66119 298934 66147 298962
rect 66181 298934 66209 298962
rect 66243 298934 66271 298962
rect 66057 298872 66085 298900
rect 66119 298872 66147 298900
rect 66181 298872 66209 298900
rect 66243 298872 66271 298900
rect 66057 293147 66085 293175
rect 66119 293147 66147 293175
rect 66181 293147 66209 293175
rect 66243 293147 66271 293175
rect 66057 293085 66085 293113
rect 66119 293085 66147 293113
rect 66181 293085 66209 293113
rect 66243 293085 66271 293113
rect 66057 293023 66085 293051
rect 66119 293023 66147 293051
rect 66181 293023 66209 293051
rect 66243 293023 66271 293051
rect 66057 292961 66085 292989
rect 66119 292961 66147 292989
rect 66181 292961 66209 292989
rect 66243 292961 66271 292989
rect 66057 284147 66085 284175
rect 66119 284147 66147 284175
rect 66181 284147 66209 284175
rect 66243 284147 66271 284175
rect 66057 284085 66085 284113
rect 66119 284085 66147 284113
rect 66181 284085 66209 284113
rect 66243 284085 66271 284113
rect 66057 284023 66085 284051
rect 66119 284023 66147 284051
rect 66181 284023 66209 284051
rect 66243 284023 66271 284051
rect 66057 283961 66085 283989
rect 66119 283961 66147 283989
rect 66181 283961 66209 283989
rect 66243 283961 66271 283989
rect 66057 275147 66085 275175
rect 66119 275147 66147 275175
rect 66181 275147 66209 275175
rect 66243 275147 66271 275175
rect 66057 275085 66085 275113
rect 66119 275085 66147 275113
rect 66181 275085 66209 275113
rect 66243 275085 66271 275113
rect 66057 275023 66085 275051
rect 66119 275023 66147 275051
rect 66181 275023 66209 275051
rect 66243 275023 66271 275051
rect 66057 274961 66085 274989
rect 66119 274961 66147 274989
rect 66181 274961 66209 274989
rect 66243 274961 66271 274989
rect 66057 266147 66085 266175
rect 66119 266147 66147 266175
rect 66181 266147 66209 266175
rect 66243 266147 66271 266175
rect 66057 266085 66085 266113
rect 66119 266085 66147 266113
rect 66181 266085 66209 266113
rect 66243 266085 66271 266113
rect 66057 266023 66085 266051
rect 66119 266023 66147 266051
rect 66181 266023 66209 266051
rect 66243 266023 66271 266051
rect 66057 265961 66085 265989
rect 66119 265961 66147 265989
rect 66181 265961 66209 265989
rect 66243 265961 66271 265989
rect 66057 257147 66085 257175
rect 66119 257147 66147 257175
rect 66181 257147 66209 257175
rect 66243 257147 66271 257175
rect 66057 257085 66085 257113
rect 66119 257085 66147 257113
rect 66181 257085 66209 257113
rect 66243 257085 66271 257113
rect 66057 257023 66085 257051
rect 66119 257023 66147 257051
rect 66181 257023 66209 257051
rect 66243 257023 66271 257051
rect 66057 256961 66085 256989
rect 66119 256961 66147 256989
rect 66181 256961 66209 256989
rect 66243 256961 66271 256989
rect 66057 248147 66085 248175
rect 66119 248147 66147 248175
rect 66181 248147 66209 248175
rect 66243 248147 66271 248175
rect 66057 248085 66085 248113
rect 66119 248085 66147 248113
rect 66181 248085 66209 248113
rect 66243 248085 66271 248113
rect 66057 248023 66085 248051
rect 66119 248023 66147 248051
rect 66181 248023 66209 248051
rect 66243 248023 66271 248051
rect 66057 247961 66085 247989
rect 66119 247961 66147 247989
rect 66181 247961 66209 247989
rect 66243 247961 66271 247989
rect 66057 239147 66085 239175
rect 66119 239147 66147 239175
rect 66181 239147 66209 239175
rect 66243 239147 66271 239175
rect 66057 239085 66085 239113
rect 66119 239085 66147 239113
rect 66181 239085 66209 239113
rect 66243 239085 66271 239113
rect 66057 239023 66085 239051
rect 66119 239023 66147 239051
rect 66181 239023 66209 239051
rect 66243 239023 66271 239051
rect 66057 238961 66085 238989
rect 66119 238961 66147 238989
rect 66181 238961 66209 238989
rect 66243 238961 66271 238989
rect 66057 230147 66085 230175
rect 66119 230147 66147 230175
rect 66181 230147 66209 230175
rect 66243 230147 66271 230175
rect 66057 230085 66085 230113
rect 66119 230085 66147 230113
rect 66181 230085 66209 230113
rect 66243 230085 66271 230113
rect 66057 230023 66085 230051
rect 66119 230023 66147 230051
rect 66181 230023 66209 230051
rect 66243 230023 66271 230051
rect 66057 229961 66085 229989
rect 66119 229961 66147 229989
rect 66181 229961 66209 229989
rect 66243 229961 66271 229989
rect 66057 221147 66085 221175
rect 66119 221147 66147 221175
rect 66181 221147 66209 221175
rect 66243 221147 66271 221175
rect 66057 221085 66085 221113
rect 66119 221085 66147 221113
rect 66181 221085 66209 221113
rect 66243 221085 66271 221113
rect 66057 221023 66085 221051
rect 66119 221023 66147 221051
rect 66181 221023 66209 221051
rect 66243 221023 66271 221051
rect 66057 220961 66085 220989
rect 66119 220961 66147 220989
rect 66181 220961 66209 220989
rect 66243 220961 66271 220989
rect 66057 212147 66085 212175
rect 66119 212147 66147 212175
rect 66181 212147 66209 212175
rect 66243 212147 66271 212175
rect 66057 212085 66085 212113
rect 66119 212085 66147 212113
rect 66181 212085 66209 212113
rect 66243 212085 66271 212113
rect 66057 212023 66085 212051
rect 66119 212023 66147 212051
rect 66181 212023 66209 212051
rect 66243 212023 66271 212051
rect 66057 211961 66085 211989
rect 66119 211961 66147 211989
rect 66181 211961 66209 211989
rect 66243 211961 66271 211989
rect 66057 203147 66085 203175
rect 66119 203147 66147 203175
rect 66181 203147 66209 203175
rect 66243 203147 66271 203175
rect 66057 203085 66085 203113
rect 66119 203085 66147 203113
rect 66181 203085 66209 203113
rect 66243 203085 66271 203113
rect 66057 203023 66085 203051
rect 66119 203023 66147 203051
rect 66181 203023 66209 203051
rect 66243 203023 66271 203051
rect 66057 202961 66085 202989
rect 66119 202961 66147 202989
rect 66181 202961 66209 202989
rect 66243 202961 66271 202989
rect 66057 194147 66085 194175
rect 66119 194147 66147 194175
rect 66181 194147 66209 194175
rect 66243 194147 66271 194175
rect 66057 194085 66085 194113
rect 66119 194085 66147 194113
rect 66181 194085 66209 194113
rect 66243 194085 66271 194113
rect 66057 194023 66085 194051
rect 66119 194023 66147 194051
rect 66181 194023 66209 194051
rect 66243 194023 66271 194051
rect 66057 193961 66085 193989
rect 66119 193961 66147 193989
rect 66181 193961 66209 193989
rect 66243 193961 66271 193989
rect 66057 185147 66085 185175
rect 66119 185147 66147 185175
rect 66181 185147 66209 185175
rect 66243 185147 66271 185175
rect 66057 185085 66085 185113
rect 66119 185085 66147 185113
rect 66181 185085 66209 185113
rect 66243 185085 66271 185113
rect 66057 185023 66085 185051
rect 66119 185023 66147 185051
rect 66181 185023 66209 185051
rect 66243 185023 66271 185051
rect 66057 184961 66085 184989
rect 66119 184961 66147 184989
rect 66181 184961 66209 184989
rect 66243 184961 66271 184989
rect 66057 176147 66085 176175
rect 66119 176147 66147 176175
rect 66181 176147 66209 176175
rect 66243 176147 66271 176175
rect 66057 176085 66085 176113
rect 66119 176085 66147 176113
rect 66181 176085 66209 176113
rect 66243 176085 66271 176113
rect 66057 176023 66085 176051
rect 66119 176023 66147 176051
rect 66181 176023 66209 176051
rect 66243 176023 66271 176051
rect 66057 175961 66085 175989
rect 66119 175961 66147 175989
rect 66181 175961 66209 175989
rect 66243 175961 66271 175989
rect 79557 298578 79585 298606
rect 79619 298578 79647 298606
rect 79681 298578 79709 298606
rect 79743 298578 79771 298606
rect 79557 298516 79585 298544
rect 79619 298516 79647 298544
rect 79681 298516 79709 298544
rect 79743 298516 79771 298544
rect 79557 298454 79585 298482
rect 79619 298454 79647 298482
rect 79681 298454 79709 298482
rect 79743 298454 79771 298482
rect 79557 298392 79585 298420
rect 79619 298392 79647 298420
rect 79681 298392 79709 298420
rect 79743 298392 79771 298420
rect 79557 290147 79585 290175
rect 79619 290147 79647 290175
rect 79681 290147 79709 290175
rect 79743 290147 79771 290175
rect 79557 290085 79585 290113
rect 79619 290085 79647 290113
rect 79681 290085 79709 290113
rect 79743 290085 79771 290113
rect 79557 290023 79585 290051
rect 79619 290023 79647 290051
rect 79681 290023 79709 290051
rect 79743 290023 79771 290051
rect 79557 289961 79585 289989
rect 79619 289961 79647 289989
rect 79681 289961 79709 289989
rect 79743 289961 79771 289989
rect 79557 281147 79585 281175
rect 79619 281147 79647 281175
rect 79681 281147 79709 281175
rect 79743 281147 79771 281175
rect 79557 281085 79585 281113
rect 79619 281085 79647 281113
rect 79681 281085 79709 281113
rect 79743 281085 79771 281113
rect 79557 281023 79585 281051
rect 79619 281023 79647 281051
rect 79681 281023 79709 281051
rect 79743 281023 79771 281051
rect 79557 280961 79585 280989
rect 79619 280961 79647 280989
rect 79681 280961 79709 280989
rect 79743 280961 79771 280989
rect 79557 272147 79585 272175
rect 79619 272147 79647 272175
rect 79681 272147 79709 272175
rect 79743 272147 79771 272175
rect 79557 272085 79585 272113
rect 79619 272085 79647 272113
rect 79681 272085 79709 272113
rect 79743 272085 79771 272113
rect 79557 272023 79585 272051
rect 79619 272023 79647 272051
rect 79681 272023 79709 272051
rect 79743 272023 79771 272051
rect 79557 271961 79585 271989
rect 79619 271961 79647 271989
rect 79681 271961 79709 271989
rect 79743 271961 79771 271989
rect 79557 263147 79585 263175
rect 79619 263147 79647 263175
rect 79681 263147 79709 263175
rect 79743 263147 79771 263175
rect 79557 263085 79585 263113
rect 79619 263085 79647 263113
rect 79681 263085 79709 263113
rect 79743 263085 79771 263113
rect 79557 263023 79585 263051
rect 79619 263023 79647 263051
rect 79681 263023 79709 263051
rect 79743 263023 79771 263051
rect 79557 262961 79585 262989
rect 79619 262961 79647 262989
rect 79681 262961 79709 262989
rect 79743 262961 79771 262989
rect 79557 254147 79585 254175
rect 79619 254147 79647 254175
rect 79681 254147 79709 254175
rect 79743 254147 79771 254175
rect 79557 254085 79585 254113
rect 79619 254085 79647 254113
rect 79681 254085 79709 254113
rect 79743 254085 79771 254113
rect 79557 254023 79585 254051
rect 79619 254023 79647 254051
rect 79681 254023 79709 254051
rect 79743 254023 79771 254051
rect 79557 253961 79585 253989
rect 79619 253961 79647 253989
rect 79681 253961 79709 253989
rect 79743 253961 79771 253989
rect 79557 245147 79585 245175
rect 79619 245147 79647 245175
rect 79681 245147 79709 245175
rect 79743 245147 79771 245175
rect 79557 245085 79585 245113
rect 79619 245085 79647 245113
rect 79681 245085 79709 245113
rect 79743 245085 79771 245113
rect 79557 245023 79585 245051
rect 79619 245023 79647 245051
rect 79681 245023 79709 245051
rect 79743 245023 79771 245051
rect 79557 244961 79585 244989
rect 79619 244961 79647 244989
rect 79681 244961 79709 244989
rect 79743 244961 79771 244989
rect 79557 236147 79585 236175
rect 79619 236147 79647 236175
rect 79681 236147 79709 236175
rect 79743 236147 79771 236175
rect 79557 236085 79585 236113
rect 79619 236085 79647 236113
rect 79681 236085 79709 236113
rect 79743 236085 79771 236113
rect 79557 236023 79585 236051
rect 79619 236023 79647 236051
rect 79681 236023 79709 236051
rect 79743 236023 79771 236051
rect 79557 235961 79585 235989
rect 79619 235961 79647 235989
rect 79681 235961 79709 235989
rect 79743 235961 79771 235989
rect 79557 227147 79585 227175
rect 79619 227147 79647 227175
rect 79681 227147 79709 227175
rect 79743 227147 79771 227175
rect 79557 227085 79585 227113
rect 79619 227085 79647 227113
rect 79681 227085 79709 227113
rect 79743 227085 79771 227113
rect 79557 227023 79585 227051
rect 79619 227023 79647 227051
rect 79681 227023 79709 227051
rect 79743 227023 79771 227051
rect 79557 226961 79585 226989
rect 79619 226961 79647 226989
rect 79681 226961 79709 226989
rect 79743 226961 79771 226989
rect 79557 218147 79585 218175
rect 79619 218147 79647 218175
rect 79681 218147 79709 218175
rect 79743 218147 79771 218175
rect 79557 218085 79585 218113
rect 79619 218085 79647 218113
rect 79681 218085 79709 218113
rect 79743 218085 79771 218113
rect 79557 218023 79585 218051
rect 79619 218023 79647 218051
rect 79681 218023 79709 218051
rect 79743 218023 79771 218051
rect 79557 217961 79585 217989
rect 79619 217961 79647 217989
rect 79681 217961 79709 217989
rect 79743 217961 79771 217989
rect 79557 209147 79585 209175
rect 79619 209147 79647 209175
rect 79681 209147 79709 209175
rect 79743 209147 79771 209175
rect 79557 209085 79585 209113
rect 79619 209085 79647 209113
rect 79681 209085 79709 209113
rect 79743 209085 79771 209113
rect 79557 209023 79585 209051
rect 79619 209023 79647 209051
rect 79681 209023 79709 209051
rect 79743 209023 79771 209051
rect 79557 208961 79585 208989
rect 79619 208961 79647 208989
rect 79681 208961 79709 208989
rect 79743 208961 79771 208989
rect 79557 200147 79585 200175
rect 79619 200147 79647 200175
rect 79681 200147 79709 200175
rect 79743 200147 79771 200175
rect 79557 200085 79585 200113
rect 79619 200085 79647 200113
rect 79681 200085 79709 200113
rect 79743 200085 79771 200113
rect 79557 200023 79585 200051
rect 79619 200023 79647 200051
rect 79681 200023 79709 200051
rect 79743 200023 79771 200051
rect 79557 199961 79585 199989
rect 79619 199961 79647 199989
rect 79681 199961 79709 199989
rect 79743 199961 79771 199989
rect 79557 191147 79585 191175
rect 79619 191147 79647 191175
rect 79681 191147 79709 191175
rect 79743 191147 79771 191175
rect 79557 191085 79585 191113
rect 79619 191085 79647 191113
rect 79681 191085 79709 191113
rect 79743 191085 79771 191113
rect 79557 191023 79585 191051
rect 79619 191023 79647 191051
rect 79681 191023 79709 191051
rect 79743 191023 79771 191051
rect 79557 190961 79585 190989
rect 79619 190961 79647 190989
rect 79681 190961 79709 190989
rect 79743 190961 79771 190989
rect 79557 182147 79585 182175
rect 79619 182147 79647 182175
rect 79681 182147 79709 182175
rect 79743 182147 79771 182175
rect 79557 182085 79585 182113
rect 79619 182085 79647 182113
rect 79681 182085 79709 182113
rect 79743 182085 79771 182113
rect 79557 182023 79585 182051
rect 79619 182023 79647 182051
rect 79681 182023 79709 182051
rect 79743 182023 79771 182051
rect 79557 181961 79585 181989
rect 79619 181961 79647 181989
rect 79681 181961 79709 181989
rect 79743 181961 79771 181989
rect 69699 173147 69727 173175
rect 69761 173147 69789 173175
rect 69699 173085 69727 173113
rect 69761 173085 69789 173113
rect 69699 173023 69727 173051
rect 69761 173023 69789 173051
rect 69699 172961 69727 172989
rect 69761 172961 69789 172989
rect 79557 173147 79585 173175
rect 79619 173147 79647 173175
rect 79681 173147 79709 173175
rect 79743 173147 79771 173175
rect 79557 173085 79585 173113
rect 79619 173085 79647 173113
rect 79681 173085 79709 173113
rect 79743 173085 79771 173113
rect 79557 173023 79585 173051
rect 79619 173023 79647 173051
rect 79681 173023 79709 173051
rect 79743 173023 79771 173051
rect 79557 172961 79585 172989
rect 79619 172961 79647 172989
rect 79681 172961 79709 172989
rect 79743 172961 79771 172989
rect 66057 167147 66085 167175
rect 66119 167147 66147 167175
rect 66181 167147 66209 167175
rect 66243 167147 66271 167175
rect 66057 167085 66085 167113
rect 66119 167085 66147 167113
rect 66181 167085 66209 167113
rect 66243 167085 66271 167113
rect 66057 167023 66085 167051
rect 66119 167023 66147 167051
rect 66181 167023 66209 167051
rect 66243 167023 66271 167051
rect 66057 166961 66085 166989
rect 66119 166961 66147 166989
rect 66181 166961 66209 166989
rect 66243 166961 66271 166989
rect 77379 167147 77407 167175
rect 77441 167147 77469 167175
rect 77379 167085 77407 167113
rect 77441 167085 77469 167113
rect 77379 167023 77407 167051
rect 77441 167023 77469 167051
rect 77379 166961 77407 166989
rect 77441 166961 77469 166989
rect 69699 164147 69727 164175
rect 69761 164147 69789 164175
rect 69699 164085 69727 164113
rect 69761 164085 69789 164113
rect 69699 164023 69727 164051
rect 69761 164023 69789 164051
rect 69699 163961 69727 163989
rect 69761 163961 69789 163989
rect 79557 164147 79585 164175
rect 79619 164147 79647 164175
rect 79681 164147 79709 164175
rect 79743 164147 79771 164175
rect 79557 164085 79585 164113
rect 79619 164085 79647 164113
rect 79681 164085 79709 164113
rect 79743 164085 79771 164113
rect 79557 164023 79585 164051
rect 79619 164023 79647 164051
rect 79681 164023 79709 164051
rect 79743 164023 79771 164051
rect 79557 163961 79585 163989
rect 79619 163961 79647 163989
rect 79681 163961 79709 163989
rect 79743 163961 79771 163989
rect 66057 158147 66085 158175
rect 66119 158147 66147 158175
rect 66181 158147 66209 158175
rect 66243 158147 66271 158175
rect 66057 158085 66085 158113
rect 66119 158085 66147 158113
rect 66181 158085 66209 158113
rect 66243 158085 66271 158113
rect 66057 158023 66085 158051
rect 66119 158023 66147 158051
rect 66181 158023 66209 158051
rect 66243 158023 66271 158051
rect 66057 157961 66085 157989
rect 66119 157961 66147 157989
rect 66181 157961 66209 157989
rect 66243 157961 66271 157989
rect 77379 158147 77407 158175
rect 77441 158147 77469 158175
rect 77379 158085 77407 158113
rect 77441 158085 77469 158113
rect 77379 158023 77407 158051
rect 77441 158023 77469 158051
rect 77379 157961 77407 157989
rect 77441 157961 77469 157989
rect 69699 155147 69727 155175
rect 69761 155147 69789 155175
rect 69699 155085 69727 155113
rect 69761 155085 69789 155113
rect 69699 155023 69727 155051
rect 69761 155023 69789 155051
rect 69699 154961 69727 154989
rect 69761 154961 69789 154989
rect 79557 155147 79585 155175
rect 79619 155147 79647 155175
rect 79681 155147 79709 155175
rect 79743 155147 79771 155175
rect 79557 155085 79585 155113
rect 79619 155085 79647 155113
rect 79681 155085 79709 155113
rect 79743 155085 79771 155113
rect 79557 155023 79585 155051
rect 79619 155023 79647 155051
rect 79681 155023 79709 155051
rect 79743 155023 79771 155051
rect 79557 154961 79585 154989
rect 79619 154961 79647 154989
rect 79681 154961 79709 154989
rect 79743 154961 79771 154989
rect 66057 149147 66085 149175
rect 66119 149147 66147 149175
rect 66181 149147 66209 149175
rect 66243 149147 66271 149175
rect 66057 149085 66085 149113
rect 66119 149085 66147 149113
rect 66181 149085 66209 149113
rect 66243 149085 66271 149113
rect 66057 149023 66085 149051
rect 66119 149023 66147 149051
rect 66181 149023 66209 149051
rect 66243 149023 66271 149051
rect 66057 148961 66085 148989
rect 66119 148961 66147 148989
rect 66181 148961 66209 148989
rect 66243 148961 66271 148989
rect 77379 149147 77407 149175
rect 77441 149147 77469 149175
rect 77379 149085 77407 149113
rect 77441 149085 77469 149113
rect 77379 149023 77407 149051
rect 77441 149023 77469 149051
rect 77379 148961 77407 148989
rect 77441 148961 77469 148989
rect 69699 146147 69727 146175
rect 69761 146147 69789 146175
rect 69699 146085 69727 146113
rect 69761 146085 69789 146113
rect 69699 146023 69727 146051
rect 69761 146023 69789 146051
rect 69699 145961 69727 145989
rect 69761 145961 69789 145989
rect 79557 146147 79585 146175
rect 79619 146147 79647 146175
rect 79681 146147 79709 146175
rect 79743 146147 79771 146175
rect 79557 146085 79585 146113
rect 79619 146085 79647 146113
rect 79681 146085 79709 146113
rect 79743 146085 79771 146113
rect 79557 146023 79585 146051
rect 79619 146023 79647 146051
rect 79681 146023 79709 146051
rect 79743 146023 79771 146051
rect 79557 145961 79585 145989
rect 79619 145961 79647 145989
rect 79681 145961 79709 145989
rect 79743 145961 79771 145989
rect 66057 140147 66085 140175
rect 66119 140147 66147 140175
rect 66181 140147 66209 140175
rect 66243 140147 66271 140175
rect 66057 140085 66085 140113
rect 66119 140085 66147 140113
rect 66181 140085 66209 140113
rect 66243 140085 66271 140113
rect 66057 140023 66085 140051
rect 66119 140023 66147 140051
rect 66181 140023 66209 140051
rect 66243 140023 66271 140051
rect 66057 139961 66085 139989
rect 66119 139961 66147 139989
rect 66181 139961 66209 139989
rect 66243 139961 66271 139989
rect 77379 140147 77407 140175
rect 77441 140147 77469 140175
rect 77379 140085 77407 140113
rect 77441 140085 77469 140113
rect 77379 140023 77407 140051
rect 77441 140023 77469 140051
rect 77379 139961 77407 139989
rect 77441 139961 77469 139989
rect 69699 137147 69727 137175
rect 69761 137147 69789 137175
rect 69699 137085 69727 137113
rect 69761 137085 69789 137113
rect 69699 137023 69727 137051
rect 69761 137023 69789 137051
rect 69699 136961 69727 136989
rect 69761 136961 69789 136989
rect 79557 137147 79585 137175
rect 79619 137147 79647 137175
rect 79681 137147 79709 137175
rect 79743 137147 79771 137175
rect 79557 137085 79585 137113
rect 79619 137085 79647 137113
rect 79681 137085 79709 137113
rect 79743 137085 79771 137113
rect 79557 137023 79585 137051
rect 79619 137023 79647 137051
rect 79681 137023 79709 137051
rect 79743 137023 79771 137051
rect 79557 136961 79585 136989
rect 79619 136961 79647 136989
rect 79681 136961 79709 136989
rect 79743 136961 79771 136989
rect 66057 131147 66085 131175
rect 66119 131147 66147 131175
rect 66181 131147 66209 131175
rect 66243 131147 66271 131175
rect 66057 131085 66085 131113
rect 66119 131085 66147 131113
rect 66181 131085 66209 131113
rect 66243 131085 66271 131113
rect 66057 131023 66085 131051
rect 66119 131023 66147 131051
rect 66181 131023 66209 131051
rect 66243 131023 66271 131051
rect 66057 130961 66085 130989
rect 66119 130961 66147 130989
rect 66181 130961 66209 130989
rect 66243 130961 66271 130989
rect 77379 131147 77407 131175
rect 77441 131147 77469 131175
rect 77379 131085 77407 131113
rect 77441 131085 77469 131113
rect 77379 131023 77407 131051
rect 77441 131023 77469 131051
rect 77379 130961 77407 130989
rect 77441 130961 77469 130989
rect 69699 128147 69727 128175
rect 69761 128147 69789 128175
rect 69699 128085 69727 128113
rect 69761 128085 69789 128113
rect 69699 128023 69727 128051
rect 69761 128023 69789 128051
rect 69699 127961 69727 127989
rect 69761 127961 69789 127989
rect 79557 128147 79585 128175
rect 79619 128147 79647 128175
rect 79681 128147 79709 128175
rect 79743 128147 79771 128175
rect 79557 128085 79585 128113
rect 79619 128085 79647 128113
rect 79681 128085 79709 128113
rect 79743 128085 79771 128113
rect 79557 128023 79585 128051
rect 79619 128023 79647 128051
rect 79681 128023 79709 128051
rect 79743 128023 79771 128051
rect 79557 127961 79585 127989
rect 79619 127961 79647 127989
rect 79681 127961 79709 127989
rect 79743 127961 79771 127989
rect 66057 122147 66085 122175
rect 66119 122147 66147 122175
rect 66181 122147 66209 122175
rect 66243 122147 66271 122175
rect 66057 122085 66085 122113
rect 66119 122085 66147 122113
rect 66181 122085 66209 122113
rect 66243 122085 66271 122113
rect 66057 122023 66085 122051
rect 66119 122023 66147 122051
rect 66181 122023 66209 122051
rect 66243 122023 66271 122051
rect 66057 121961 66085 121989
rect 66119 121961 66147 121989
rect 66181 121961 66209 121989
rect 66243 121961 66271 121989
rect 77379 122147 77407 122175
rect 77441 122147 77469 122175
rect 77379 122085 77407 122113
rect 77441 122085 77469 122113
rect 77379 122023 77407 122051
rect 77441 122023 77469 122051
rect 77379 121961 77407 121989
rect 77441 121961 77469 121989
rect 69699 119147 69727 119175
rect 69761 119147 69789 119175
rect 69699 119085 69727 119113
rect 69761 119085 69789 119113
rect 69699 119023 69727 119051
rect 69761 119023 69789 119051
rect 69699 118961 69727 118989
rect 69761 118961 69789 118989
rect 79557 119147 79585 119175
rect 79619 119147 79647 119175
rect 79681 119147 79709 119175
rect 79743 119147 79771 119175
rect 79557 119085 79585 119113
rect 79619 119085 79647 119113
rect 79681 119085 79709 119113
rect 79743 119085 79771 119113
rect 79557 119023 79585 119051
rect 79619 119023 79647 119051
rect 79681 119023 79709 119051
rect 79743 119023 79771 119051
rect 79557 118961 79585 118989
rect 79619 118961 79647 118989
rect 79681 118961 79709 118989
rect 79743 118961 79771 118989
rect 66057 113147 66085 113175
rect 66119 113147 66147 113175
rect 66181 113147 66209 113175
rect 66243 113147 66271 113175
rect 66057 113085 66085 113113
rect 66119 113085 66147 113113
rect 66181 113085 66209 113113
rect 66243 113085 66271 113113
rect 66057 113023 66085 113051
rect 66119 113023 66147 113051
rect 66181 113023 66209 113051
rect 66243 113023 66271 113051
rect 66057 112961 66085 112989
rect 66119 112961 66147 112989
rect 66181 112961 66209 112989
rect 66243 112961 66271 112989
rect 77379 113147 77407 113175
rect 77441 113147 77469 113175
rect 77379 113085 77407 113113
rect 77441 113085 77469 113113
rect 77379 113023 77407 113051
rect 77441 113023 77469 113051
rect 77379 112961 77407 112989
rect 77441 112961 77469 112989
rect 69699 110147 69727 110175
rect 69761 110147 69789 110175
rect 69699 110085 69727 110113
rect 69761 110085 69789 110113
rect 69699 110023 69727 110051
rect 69761 110023 69789 110051
rect 69699 109961 69727 109989
rect 69761 109961 69789 109989
rect 79557 110147 79585 110175
rect 79619 110147 79647 110175
rect 79681 110147 79709 110175
rect 79743 110147 79771 110175
rect 79557 110085 79585 110113
rect 79619 110085 79647 110113
rect 79681 110085 79709 110113
rect 79743 110085 79771 110113
rect 79557 110023 79585 110051
rect 79619 110023 79647 110051
rect 79681 110023 79709 110051
rect 79743 110023 79771 110051
rect 79557 109961 79585 109989
rect 79619 109961 79647 109989
rect 79681 109961 79709 109989
rect 79743 109961 79771 109989
rect 66057 104147 66085 104175
rect 66119 104147 66147 104175
rect 66181 104147 66209 104175
rect 66243 104147 66271 104175
rect 66057 104085 66085 104113
rect 66119 104085 66147 104113
rect 66181 104085 66209 104113
rect 66243 104085 66271 104113
rect 66057 104023 66085 104051
rect 66119 104023 66147 104051
rect 66181 104023 66209 104051
rect 66243 104023 66271 104051
rect 66057 103961 66085 103989
rect 66119 103961 66147 103989
rect 66181 103961 66209 103989
rect 66243 103961 66271 103989
rect 77379 104147 77407 104175
rect 77441 104147 77469 104175
rect 77379 104085 77407 104113
rect 77441 104085 77469 104113
rect 77379 104023 77407 104051
rect 77441 104023 77469 104051
rect 77379 103961 77407 103989
rect 77441 103961 77469 103989
rect 69699 101147 69727 101175
rect 69761 101147 69789 101175
rect 69699 101085 69727 101113
rect 69761 101085 69789 101113
rect 69699 101023 69727 101051
rect 69761 101023 69789 101051
rect 69699 100961 69727 100989
rect 69761 100961 69789 100989
rect 79557 101147 79585 101175
rect 79619 101147 79647 101175
rect 79681 101147 79709 101175
rect 79743 101147 79771 101175
rect 79557 101085 79585 101113
rect 79619 101085 79647 101113
rect 79681 101085 79709 101113
rect 79743 101085 79771 101113
rect 79557 101023 79585 101051
rect 79619 101023 79647 101051
rect 79681 101023 79709 101051
rect 79743 101023 79771 101051
rect 79557 100961 79585 100989
rect 79619 100961 79647 100989
rect 79681 100961 79709 100989
rect 79743 100961 79771 100989
rect 66057 95147 66085 95175
rect 66119 95147 66147 95175
rect 66181 95147 66209 95175
rect 66243 95147 66271 95175
rect 66057 95085 66085 95113
rect 66119 95085 66147 95113
rect 66181 95085 66209 95113
rect 66243 95085 66271 95113
rect 66057 95023 66085 95051
rect 66119 95023 66147 95051
rect 66181 95023 66209 95051
rect 66243 95023 66271 95051
rect 66057 94961 66085 94989
rect 66119 94961 66147 94989
rect 66181 94961 66209 94989
rect 66243 94961 66271 94989
rect 77379 95147 77407 95175
rect 77441 95147 77469 95175
rect 77379 95085 77407 95113
rect 77441 95085 77469 95113
rect 77379 95023 77407 95051
rect 77441 95023 77469 95051
rect 77379 94961 77407 94989
rect 77441 94961 77469 94989
rect 69699 92147 69727 92175
rect 69761 92147 69789 92175
rect 69699 92085 69727 92113
rect 69761 92085 69789 92113
rect 69699 92023 69727 92051
rect 69761 92023 69789 92051
rect 69699 91961 69727 91989
rect 69761 91961 69789 91989
rect 79557 92147 79585 92175
rect 79619 92147 79647 92175
rect 79681 92147 79709 92175
rect 79743 92147 79771 92175
rect 79557 92085 79585 92113
rect 79619 92085 79647 92113
rect 79681 92085 79709 92113
rect 79743 92085 79771 92113
rect 79557 92023 79585 92051
rect 79619 92023 79647 92051
rect 79681 92023 79709 92051
rect 79743 92023 79771 92051
rect 79557 91961 79585 91989
rect 79619 91961 79647 91989
rect 79681 91961 79709 91989
rect 79743 91961 79771 91989
rect 66057 86147 66085 86175
rect 66119 86147 66147 86175
rect 66181 86147 66209 86175
rect 66243 86147 66271 86175
rect 66057 86085 66085 86113
rect 66119 86085 66147 86113
rect 66181 86085 66209 86113
rect 66243 86085 66271 86113
rect 66057 86023 66085 86051
rect 66119 86023 66147 86051
rect 66181 86023 66209 86051
rect 66243 86023 66271 86051
rect 66057 85961 66085 85989
rect 66119 85961 66147 85989
rect 66181 85961 66209 85989
rect 66243 85961 66271 85989
rect 77379 86147 77407 86175
rect 77441 86147 77469 86175
rect 77379 86085 77407 86113
rect 77441 86085 77469 86113
rect 77379 86023 77407 86051
rect 77441 86023 77469 86051
rect 77379 85961 77407 85989
rect 77441 85961 77469 85989
rect 69699 83147 69727 83175
rect 69761 83147 69789 83175
rect 69699 83085 69727 83113
rect 69761 83085 69789 83113
rect 69699 83023 69727 83051
rect 69761 83023 69789 83051
rect 69699 82961 69727 82989
rect 69761 82961 69789 82989
rect 79557 83147 79585 83175
rect 79619 83147 79647 83175
rect 79681 83147 79709 83175
rect 79743 83147 79771 83175
rect 79557 83085 79585 83113
rect 79619 83085 79647 83113
rect 79681 83085 79709 83113
rect 79743 83085 79771 83113
rect 79557 83023 79585 83051
rect 79619 83023 79647 83051
rect 79681 83023 79709 83051
rect 79743 83023 79771 83051
rect 79557 82961 79585 82989
rect 79619 82961 79647 82989
rect 79681 82961 79709 82989
rect 79743 82961 79771 82989
rect 66057 77147 66085 77175
rect 66119 77147 66147 77175
rect 66181 77147 66209 77175
rect 66243 77147 66271 77175
rect 66057 77085 66085 77113
rect 66119 77085 66147 77113
rect 66181 77085 66209 77113
rect 66243 77085 66271 77113
rect 66057 77023 66085 77051
rect 66119 77023 66147 77051
rect 66181 77023 66209 77051
rect 66243 77023 66271 77051
rect 66057 76961 66085 76989
rect 66119 76961 66147 76989
rect 66181 76961 66209 76989
rect 66243 76961 66271 76989
rect 77379 77147 77407 77175
rect 77441 77147 77469 77175
rect 77379 77085 77407 77113
rect 77441 77085 77469 77113
rect 77379 77023 77407 77051
rect 77441 77023 77469 77051
rect 77379 76961 77407 76989
rect 77441 76961 77469 76989
rect 69699 74147 69727 74175
rect 69761 74147 69789 74175
rect 69699 74085 69727 74113
rect 69761 74085 69789 74113
rect 69699 74023 69727 74051
rect 69761 74023 69789 74051
rect 69699 73961 69727 73989
rect 69761 73961 69789 73989
rect 79557 74147 79585 74175
rect 79619 74147 79647 74175
rect 79681 74147 79709 74175
rect 79743 74147 79771 74175
rect 79557 74085 79585 74113
rect 79619 74085 79647 74113
rect 79681 74085 79709 74113
rect 79743 74085 79771 74113
rect 79557 74023 79585 74051
rect 79619 74023 79647 74051
rect 79681 74023 79709 74051
rect 79743 74023 79771 74051
rect 79557 73961 79585 73989
rect 79619 73961 79647 73989
rect 79681 73961 79709 73989
rect 79743 73961 79771 73989
rect 66057 68147 66085 68175
rect 66119 68147 66147 68175
rect 66181 68147 66209 68175
rect 66243 68147 66271 68175
rect 66057 68085 66085 68113
rect 66119 68085 66147 68113
rect 66181 68085 66209 68113
rect 66243 68085 66271 68113
rect 66057 68023 66085 68051
rect 66119 68023 66147 68051
rect 66181 68023 66209 68051
rect 66243 68023 66271 68051
rect 66057 67961 66085 67989
rect 66119 67961 66147 67989
rect 66181 67961 66209 67989
rect 66243 67961 66271 67989
rect 77379 68147 77407 68175
rect 77441 68147 77469 68175
rect 77379 68085 77407 68113
rect 77441 68085 77469 68113
rect 77379 68023 77407 68051
rect 77441 68023 77469 68051
rect 77379 67961 77407 67989
rect 77441 67961 77469 67989
rect 69699 65147 69727 65175
rect 69761 65147 69789 65175
rect 69699 65085 69727 65113
rect 69761 65085 69789 65113
rect 69699 65023 69727 65051
rect 69761 65023 69789 65051
rect 69699 64961 69727 64989
rect 69761 64961 69789 64989
rect 79557 65147 79585 65175
rect 79619 65147 79647 65175
rect 79681 65147 79709 65175
rect 79743 65147 79771 65175
rect 79557 65085 79585 65113
rect 79619 65085 79647 65113
rect 79681 65085 79709 65113
rect 79743 65085 79771 65113
rect 79557 65023 79585 65051
rect 79619 65023 79647 65051
rect 79681 65023 79709 65051
rect 79743 65023 79771 65051
rect 79557 64961 79585 64989
rect 79619 64961 79647 64989
rect 79681 64961 79709 64989
rect 79743 64961 79771 64989
rect 66057 59147 66085 59175
rect 66119 59147 66147 59175
rect 66181 59147 66209 59175
rect 66243 59147 66271 59175
rect 66057 59085 66085 59113
rect 66119 59085 66147 59113
rect 66181 59085 66209 59113
rect 66243 59085 66271 59113
rect 66057 59023 66085 59051
rect 66119 59023 66147 59051
rect 66181 59023 66209 59051
rect 66243 59023 66271 59051
rect 66057 58961 66085 58989
rect 66119 58961 66147 58989
rect 66181 58961 66209 58989
rect 66243 58961 66271 58989
rect 77379 59147 77407 59175
rect 77441 59147 77469 59175
rect 77379 59085 77407 59113
rect 77441 59085 77469 59113
rect 77379 59023 77407 59051
rect 77441 59023 77469 59051
rect 77379 58961 77407 58989
rect 77441 58961 77469 58989
rect 69699 56147 69727 56175
rect 69761 56147 69789 56175
rect 69699 56085 69727 56113
rect 69761 56085 69789 56113
rect 69699 56023 69727 56051
rect 69761 56023 69789 56051
rect 69699 55961 69727 55989
rect 69761 55961 69789 55989
rect 79557 56147 79585 56175
rect 79619 56147 79647 56175
rect 79681 56147 79709 56175
rect 79743 56147 79771 56175
rect 79557 56085 79585 56113
rect 79619 56085 79647 56113
rect 79681 56085 79709 56113
rect 79743 56085 79771 56113
rect 79557 56023 79585 56051
rect 79619 56023 79647 56051
rect 79681 56023 79709 56051
rect 79743 56023 79771 56051
rect 79557 55961 79585 55989
rect 79619 55961 79647 55989
rect 79681 55961 79709 55989
rect 79743 55961 79771 55989
rect 66057 50147 66085 50175
rect 66119 50147 66147 50175
rect 66181 50147 66209 50175
rect 66243 50147 66271 50175
rect 66057 50085 66085 50113
rect 66119 50085 66147 50113
rect 66181 50085 66209 50113
rect 66243 50085 66271 50113
rect 66057 50023 66085 50051
rect 66119 50023 66147 50051
rect 66181 50023 66209 50051
rect 66243 50023 66271 50051
rect 66057 49961 66085 49989
rect 66119 49961 66147 49989
rect 66181 49961 66209 49989
rect 66243 49961 66271 49989
rect 77379 50147 77407 50175
rect 77441 50147 77469 50175
rect 77379 50085 77407 50113
rect 77441 50085 77469 50113
rect 77379 50023 77407 50051
rect 77441 50023 77469 50051
rect 77379 49961 77407 49989
rect 77441 49961 77469 49989
rect 69699 47147 69727 47175
rect 69761 47147 69789 47175
rect 69699 47085 69727 47113
rect 69761 47085 69789 47113
rect 69699 47023 69727 47051
rect 69761 47023 69789 47051
rect 69699 46961 69727 46989
rect 69761 46961 69789 46989
rect 79557 47147 79585 47175
rect 79619 47147 79647 47175
rect 79681 47147 79709 47175
rect 79743 47147 79771 47175
rect 79557 47085 79585 47113
rect 79619 47085 79647 47113
rect 79681 47085 79709 47113
rect 79743 47085 79771 47113
rect 79557 47023 79585 47051
rect 79619 47023 79647 47051
rect 79681 47023 79709 47051
rect 79743 47023 79771 47051
rect 79557 46961 79585 46989
rect 79619 46961 79647 46989
rect 79681 46961 79709 46989
rect 79743 46961 79771 46989
rect 66057 41147 66085 41175
rect 66119 41147 66147 41175
rect 66181 41147 66209 41175
rect 66243 41147 66271 41175
rect 66057 41085 66085 41113
rect 66119 41085 66147 41113
rect 66181 41085 66209 41113
rect 66243 41085 66271 41113
rect 66057 41023 66085 41051
rect 66119 41023 66147 41051
rect 66181 41023 66209 41051
rect 66243 41023 66271 41051
rect 66057 40961 66085 40989
rect 66119 40961 66147 40989
rect 66181 40961 66209 40989
rect 66243 40961 66271 40989
rect 77379 41147 77407 41175
rect 77441 41147 77469 41175
rect 77379 41085 77407 41113
rect 77441 41085 77469 41113
rect 77379 41023 77407 41051
rect 77441 41023 77469 41051
rect 77379 40961 77407 40989
rect 77441 40961 77469 40989
rect 69699 38147 69727 38175
rect 69761 38147 69789 38175
rect 69699 38085 69727 38113
rect 69761 38085 69789 38113
rect 69699 38023 69727 38051
rect 69761 38023 69789 38051
rect 69699 37961 69727 37989
rect 69761 37961 69789 37989
rect 79557 38147 79585 38175
rect 79619 38147 79647 38175
rect 79681 38147 79709 38175
rect 79743 38147 79771 38175
rect 79557 38085 79585 38113
rect 79619 38085 79647 38113
rect 79681 38085 79709 38113
rect 79743 38085 79771 38113
rect 79557 38023 79585 38051
rect 79619 38023 79647 38051
rect 79681 38023 79709 38051
rect 79743 38023 79771 38051
rect 79557 37961 79585 37989
rect 79619 37961 79647 37989
rect 79681 37961 79709 37989
rect 79743 37961 79771 37989
rect 66057 32147 66085 32175
rect 66119 32147 66147 32175
rect 66181 32147 66209 32175
rect 66243 32147 66271 32175
rect 66057 32085 66085 32113
rect 66119 32085 66147 32113
rect 66181 32085 66209 32113
rect 66243 32085 66271 32113
rect 66057 32023 66085 32051
rect 66119 32023 66147 32051
rect 66181 32023 66209 32051
rect 66243 32023 66271 32051
rect 66057 31961 66085 31989
rect 66119 31961 66147 31989
rect 66181 31961 66209 31989
rect 66243 31961 66271 31989
rect 77379 32147 77407 32175
rect 77441 32147 77469 32175
rect 77379 32085 77407 32113
rect 77441 32085 77469 32113
rect 77379 32023 77407 32051
rect 77441 32023 77469 32051
rect 77379 31961 77407 31989
rect 77441 31961 77469 31989
rect 69699 29147 69727 29175
rect 69761 29147 69789 29175
rect 69699 29085 69727 29113
rect 69761 29085 69789 29113
rect 69699 29023 69727 29051
rect 69761 29023 69789 29051
rect 69699 28961 69727 28989
rect 69761 28961 69789 28989
rect 79557 29147 79585 29175
rect 79619 29147 79647 29175
rect 79681 29147 79709 29175
rect 79743 29147 79771 29175
rect 79557 29085 79585 29113
rect 79619 29085 79647 29113
rect 79681 29085 79709 29113
rect 79743 29085 79771 29113
rect 79557 29023 79585 29051
rect 79619 29023 79647 29051
rect 79681 29023 79709 29051
rect 79743 29023 79771 29051
rect 79557 28961 79585 28989
rect 79619 28961 79647 28989
rect 79681 28961 79709 28989
rect 79743 28961 79771 28989
rect 66057 23147 66085 23175
rect 66119 23147 66147 23175
rect 66181 23147 66209 23175
rect 66243 23147 66271 23175
rect 66057 23085 66085 23113
rect 66119 23085 66147 23113
rect 66181 23085 66209 23113
rect 66243 23085 66271 23113
rect 66057 23023 66085 23051
rect 66119 23023 66147 23051
rect 66181 23023 66209 23051
rect 66243 23023 66271 23051
rect 66057 22961 66085 22989
rect 66119 22961 66147 22989
rect 66181 22961 66209 22989
rect 66243 22961 66271 22989
rect 77379 23147 77407 23175
rect 77441 23147 77469 23175
rect 77379 23085 77407 23113
rect 77441 23085 77469 23113
rect 77379 23023 77407 23051
rect 77441 23023 77469 23051
rect 77379 22961 77407 22989
rect 77441 22961 77469 22989
rect 69699 20147 69727 20175
rect 69761 20147 69789 20175
rect 69699 20085 69727 20113
rect 69761 20085 69789 20113
rect 69699 20023 69727 20051
rect 69761 20023 69789 20051
rect 69699 19961 69727 19989
rect 69761 19961 69789 19989
rect 79557 20147 79585 20175
rect 79619 20147 79647 20175
rect 79681 20147 79709 20175
rect 79743 20147 79771 20175
rect 79557 20085 79585 20113
rect 79619 20085 79647 20113
rect 79681 20085 79709 20113
rect 79743 20085 79771 20113
rect 79557 20023 79585 20051
rect 79619 20023 79647 20051
rect 79681 20023 79709 20051
rect 79743 20023 79771 20051
rect 79557 19961 79585 19989
rect 79619 19961 79647 19989
rect 79681 19961 79709 19989
rect 79743 19961 79771 19989
rect 66057 14147 66085 14175
rect 66119 14147 66147 14175
rect 66181 14147 66209 14175
rect 66243 14147 66271 14175
rect 66057 14085 66085 14113
rect 66119 14085 66147 14113
rect 66181 14085 66209 14113
rect 66243 14085 66271 14113
rect 66057 14023 66085 14051
rect 66119 14023 66147 14051
rect 66181 14023 66209 14051
rect 66243 14023 66271 14051
rect 66057 13961 66085 13989
rect 66119 13961 66147 13989
rect 66181 13961 66209 13989
rect 66243 13961 66271 13989
rect 77379 14147 77407 14175
rect 77441 14147 77469 14175
rect 77379 14085 77407 14113
rect 77441 14085 77469 14113
rect 77379 14023 77407 14051
rect 77441 14023 77469 14051
rect 77379 13961 77407 13989
rect 77441 13961 77469 13989
rect 69699 11147 69727 11175
rect 69761 11147 69789 11175
rect 69699 11085 69727 11113
rect 69761 11085 69789 11113
rect 69699 11023 69727 11051
rect 69761 11023 69789 11051
rect 69699 10961 69727 10989
rect 69761 10961 69789 10989
rect 79557 11147 79585 11175
rect 79619 11147 79647 11175
rect 79681 11147 79709 11175
rect 79743 11147 79771 11175
rect 79557 11085 79585 11113
rect 79619 11085 79647 11113
rect 79681 11085 79709 11113
rect 79743 11085 79771 11113
rect 79557 11023 79585 11051
rect 79619 11023 79647 11051
rect 79681 11023 79709 11051
rect 79743 11023 79771 11051
rect 79557 10961 79585 10989
rect 79619 10961 79647 10989
rect 79681 10961 79709 10989
rect 79743 10961 79771 10989
rect 66057 5147 66085 5175
rect 66119 5147 66147 5175
rect 66181 5147 66209 5175
rect 66243 5147 66271 5175
rect 66057 5085 66085 5113
rect 66119 5085 66147 5113
rect 66181 5085 66209 5113
rect 66243 5085 66271 5113
rect 66057 5023 66085 5051
rect 66119 5023 66147 5051
rect 66181 5023 66209 5051
rect 66243 5023 66271 5051
rect 66057 4961 66085 4989
rect 66119 4961 66147 4989
rect 66181 4961 66209 4989
rect 66243 4961 66271 4989
rect 77379 5147 77407 5175
rect 77441 5147 77469 5175
rect 77379 5085 77407 5113
rect 77441 5085 77469 5113
rect 77379 5023 77407 5051
rect 77441 5023 77469 5051
rect 77379 4961 77407 4989
rect 77441 4961 77469 4989
rect 66057 -588 66085 -560
rect 66119 -588 66147 -560
rect 66181 -588 66209 -560
rect 66243 -588 66271 -560
rect 66057 -650 66085 -622
rect 66119 -650 66147 -622
rect 66181 -650 66209 -622
rect 66243 -650 66271 -622
rect 66057 -712 66085 -684
rect 66119 -712 66147 -684
rect 66181 -712 66209 -684
rect 66243 -712 66271 -684
rect 66057 -774 66085 -746
rect 66119 -774 66147 -746
rect 66181 -774 66209 -746
rect 66243 -774 66271 -746
rect 79557 2147 79585 2175
rect 79619 2147 79647 2175
rect 79681 2147 79709 2175
rect 79743 2147 79771 2175
rect 79557 2085 79585 2113
rect 79619 2085 79647 2113
rect 79681 2085 79709 2113
rect 79743 2085 79771 2113
rect 79557 2023 79585 2051
rect 79619 2023 79647 2051
rect 79681 2023 79709 2051
rect 79743 2023 79771 2051
rect 79557 1961 79585 1989
rect 79619 1961 79647 1989
rect 79681 1961 79709 1989
rect 79743 1961 79771 1989
rect 79557 -108 79585 -80
rect 79619 -108 79647 -80
rect 79681 -108 79709 -80
rect 79743 -108 79771 -80
rect 79557 -170 79585 -142
rect 79619 -170 79647 -142
rect 79681 -170 79709 -142
rect 79743 -170 79771 -142
rect 79557 -232 79585 -204
rect 79619 -232 79647 -204
rect 79681 -232 79709 -204
rect 79743 -232 79771 -204
rect 79557 -294 79585 -266
rect 79619 -294 79647 -266
rect 79681 -294 79709 -266
rect 79743 -294 79771 -266
rect 81417 299058 81445 299086
rect 81479 299058 81507 299086
rect 81541 299058 81569 299086
rect 81603 299058 81631 299086
rect 81417 298996 81445 299024
rect 81479 298996 81507 299024
rect 81541 298996 81569 299024
rect 81603 298996 81631 299024
rect 81417 298934 81445 298962
rect 81479 298934 81507 298962
rect 81541 298934 81569 298962
rect 81603 298934 81631 298962
rect 81417 298872 81445 298900
rect 81479 298872 81507 298900
rect 81541 298872 81569 298900
rect 81603 298872 81631 298900
rect 81417 293147 81445 293175
rect 81479 293147 81507 293175
rect 81541 293147 81569 293175
rect 81603 293147 81631 293175
rect 81417 293085 81445 293113
rect 81479 293085 81507 293113
rect 81541 293085 81569 293113
rect 81603 293085 81631 293113
rect 81417 293023 81445 293051
rect 81479 293023 81507 293051
rect 81541 293023 81569 293051
rect 81603 293023 81631 293051
rect 81417 292961 81445 292989
rect 81479 292961 81507 292989
rect 81541 292961 81569 292989
rect 81603 292961 81631 292989
rect 81417 284147 81445 284175
rect 81479 284147 81507 284175
rect 81541 284147 81569 284175
rect 81603 284147 81631 284175
rect 81417 284085 81445 284113
rect 81479 284085 81507 284113
rect 81541 284085 81569 284113
rect 81603 284085 81631 284113
rect 81417 284023 81445 284051
rect 81479 284023 81507 284051
rect 81541 284023 81569 284051
rect 81603 284023 81631 284051
rect 81417 283961 81445 283989
rect 81479 283961 81507 283989
rect 81541 283961 81569 283989
rect 81603 283961 81631 283989
rect 81417 275147 81445 275175
rect 81479 275147 81507 275175
rect 81541 275147 81569 275175
rect 81603 275147 81631 275175
rect 81417 275085 81445 275113
rect 81479 275085 81507 275113
rect 81541 275085 81569 275113
rect 81603 275085 81631 275113
rect 81417 275023 81445 275051
rect 81479 275023 81507 275051
rect 81541 275023 81569 275051
rect 81603 275023 81631 275051
rect 81417 274961 81445 274989
rect 81479 274961 81507 274989
rect 81541 274961 81569 274989
rect 81603 274961 81631 274989
rect 81417 266147 81445 266175
rect 81479 266147 81507 266175
rect 81541 266147 81569 266175
rect 81603 266147 81631 266175
rect 81417 266085 81445 266113
rect 81479 266085 81507 266113
rect 81541 266085 81569 266113
rect 81603 266085 81631 266113
rect 81417 266023 81445 266051
rect 81479 266023 81507 266051
rect 81541 266023 81569 266051
rect 81603 266023 81631 266051
rect 81417 265961 81445 265989
rect 81479 265961 81507 265989
rect 81541 265961 81569 265989
rect 81603 265961 81631 265989
rect 81417 257147 81445 257175
rect 81479 257147 81507 257175
rect 81541 257147 81569 257175
rect 81603 257147 81631 257175
rect 81417 257085 81445 257113
rect 81479 257085 81507 257113
rect 81541 257085 81569 257113
rect 81603 257085 81631 257113
rect 81417 257023 81445 257051
rect 81479 257023 81507 257051
rect 81541 257023 81569 257051
rect 81603 257023 81631 257051
rect 81417 256961 81445 256989
rect 81479 256961 81507 256989
rect 81541 256961 81569 256989
rect 81603 256961 81631 256989
rect 81417 248147 81445 248175
rect 81479 248147 81507 248175
rect 81541 248147 81569 248175
rect 81603 248147 81631 248175
rect 81417 248085 81445 248113
rect 81479 248085 81507 248113
rect 81541 248085 81569 248113
rect 81603 248085 81631 248113
rect 81417 248023 81445 248051
rect 81479 248023 81507 248051
rect 81541 248023 81569 248051
rect 81603 248023 81631 248051
rect 81417 247961 81445 247989
rect 81479 247961 81507 247989
rect 81541 247961 81569 247989
rect 81603 247961 81631 247989
rect 81417 239147 81445 239175
rect 81479 239147 81507 239175
rect 81541 239147 81569 239175
rect 81603 239147 81631 239175
rect 81417 239085 81445 239113
rect 81479 239085 81507 239113
rect 81541 239085 81569 239113
rect 81603 239085 81631 239113
rect 81417 239023 81445 239051
rect 81479 239023 81507 239051
rect 81541 239023 81569 239051
rect 81603 239023 81631 239051
rect 81417 238961 81445 238989
rect 81479 238961 81507 238989
rect 81541 238961 81569 238989
rect 81603 238961 81631 238989
rect 81417 230147 81445 230175
rect 81479 230147 81507 230175
rect 81541 230147 81569 230175
rect 81603 230147 81631 230175
rect 81417 230085 81445 230113
rect 81479 230085 81507 230113
rect 81541 230085 81569 230113
rect 81603 230085 81631 230113
rect 81417 230023 81445 230051
rect 81479 230023 81507 230051
rect 81541 230023 81569 230051
rect 81603 230023 81631 230051
rect 81417 229961 81445 229989
rect 81479 229961 81507 229989
rect 81541 229961 81569 229989
rect 81603 229961 81631 229989
rect 81417 221147 81445 221175
rect 81479 221147 81507 221175
rect 81541 221147 81569 221175
rect 81603 221147 81631 221175
rect 81417 221085 81445 221113
rect 81479 221085 81507 221113
rect 81541 221085 81569 221113
rect 81603 221085 81631 221113
rect 81417 221023 81445 221051
rect 81479 221023 81507 221051
rect 81541 221023 81569 221051
rect 81603 221023 81631 221051
rect 81417 220961 81445 220989
rect 81479 220961 81507 220989
rect 81541 220961 81569 220989
rect 81603 220961 81631 220989
rect 81417 212147 81445 212175
rect 81479 212147 81507 212175
rect 81541 212147 81569 212175
rect 81603 212147 81631 212175
rect 81417 212085 81445 212113
rect 81479 212085 81507 212113
rect 81541 212085 81569 212113
rect 81603 212085 81631 212113
rect 81417 212023 81445 212051
rect 81479 212023 81507 212051
rect 81541 212023 81569 212051
rect 81603 212023 81631 212051
rect 81417 211961 81445 211989
rect 81479 211961 81507 211989
rect 81541 211961 81569 211989
rect 81603 211961 81631 211989
rect 81417 203147 81445 203175
rect 81479 203147 81507 203175
rect 81541 203147 81569 203175
rect 81603 203147 81631 203175
rect 81417 203085 81445 203113
rect 81479 203085 81507 203113
rect 81541 203085 81569 203113
rect 81603 203085 81631 203113
rect 81417 203023 81445 203051
rect 81479 203023 81507 203051
rect 81541 203023 81569 203051
rect 81603 203023 81631 203051
rect 81417 202961 81445 202989
rect 81479 202961 81507 202989
rect 81541 202961 81569 202989
rect 81603 202961 81631 202989
rect 81417 194147 81445 194175
rect 81479 194147 81507 194175
rect 81541 194147 81569 194175
rect 81603 194147 81631 194175
rect 81417 194085 81445 194113
rect 81479 194085 81507 194113
rect 81541 194085 81569 194113
rect 81603 194085 81631 194113
rect 81417 194023 81445 194051
rect 81479 194023 81507 194051
rect 81541 194023 81569 194051
rect 81603 194023 81631 194051
rect 81417 193961 81445 193989
rect 81479 193961 81507 193989
rect 81541 193961 81569 193989
rect 81603 193961 81631 193989
rect 81417 185147 81445 185175
rect 81479 185147 81507 185175
rect 81541 185147 81569 185175
rect 81603 185147 81631 185175
rect 81417 185085 81445 185113
rect 81479 185085 81507 185113
rect 81541 185085 81569 185113
rect 81603 185085 81631 185113
rect 81417 185023 81445 185051
rect 81479 185023 81507 185051
rect 81541 185023 81569 185051
rect 81603 185023 81631 185051
rect 81417 184961 81445 184989
rect 81479 184961 81507 184989
rect 81541 184961 81569 184989
rect 81603 184961 81631 184989
rect 81417 176147 81445 176175
rect 81479 176147 81507 176175
rect 81541 176147 81569 176175
rect 81603 176147 81631 176175
rect 81417 176085 81445 176113
rect 81479 176085 81507 176113
rect 81541 176085 81569 176113
rect 81603 176085 81631 176113
rect 81417 176023 81445 176051
rect 81479 176023 81507 176051
rect 81541 176023 81569 176051
rect 81603 176023 81631 176051
rect 81417 175961 81445 175989
rect 81479 175961 81507 175989
rect 81541 175961 81569 175989
rect 81603 175961 81631 175989
rect 94917 298578 94945 298606
rect 94979 298578 95007 298606
rect 95041 298578 95069 298606
rect 95103 298578 95131 298606
rect 94917 298516 94945 298544
rect 94979 298516 95007 298544
rect 95041 298516 95069 298544
rect 95103 298516 95131 298544
rect 94917 298454 94945 298482
rect 94979 298454 95007 298482
rect 95041 298454 95069 298482
rect 95103 298454 95131 298482
rect 94917 298392 94945 298420
rect 94979 298392 95007 298420
rect 95041 298392 95069 298420
rect 95103 298392 95131 298420
rect 94917 290147 94945 290175
rect 94979 290147 95007 290175
rect 95041 290147 95069 290175
rect 95103 290147 95131 290175
rect 94917 290085 94945 290113
rect 94979 290085 95007 290113
rect 95041 290085 95069 290113
rect 95103 290085 95131 290113
rect 94917 290023 94945 290051
rect 94979 290023 95007 290051
rect 95041 290023 95069 290051
rect 95103 290023 95131 290051
rect 94917 289961 94945 289989
rect 94979 289961 95007 289989
rect 95041 289961 95069 289989
rect 95103 289961 95131 289989
rect 94917 281147 94945 281175
rect 94979 281147 95007 281175
rect 95041 281147 95069 281175
rect 95103 281147 95131 281175
rect 94917 281085 94945 281113
rect 94979 281085 95007 281113
rect 95041 281085 95069 281113
rect 95103 281085 95131 281113
rect 94917 281023 94945 281051
rect 94979 281023 95007 281051
rect 95041 281023 95069 281051
rect 95103 281023 95131 281051
rect 94917 280961 94945 280989
rect 94979 280961 95007 280989
rect 95041 280961 95069 280989
rect 95103 280961 95131 280989
rect 94917 272147 94945 272175
rect 94979 272147 95007 272175
rect 95041 272147 95069 272175
rect 95103 272147 95131 272175
rect 94917 272085 94945 272113
rect 94979 272085 95007 272113
rect 95041 272085 95069 272113
rect 95103 272085 95131 272113
rect 94917 272023 94945 272051
rect 94979 272023 95007 272051
rect 95041 272023 95069 272051
rect 95103 272023 95131 272051
rect 94917 271961 94945 271989
rect 94979 271961 95007 271989
rect 95041 271961 95069 271989
rect 95103 271961 95131 271989
rect 94917 263147 94945 263175
rect 94979 263147 95007 263175
rect 95041 263147 95069 263175
rect 95103 263147 95131 263175
rect 94917 263085 94945 263113
rect 94979 263085 95007 263113
rect 95041 263085 95069 263113
rect 95103 263085 95131 263113
rect 94917 263023 94945 263051
rect 94979 263023 95007 263051
rect 95041 263023 95069 263051
rect 95103 263023 95131 263051
rect 94917 262961 94945 262989
rect 94979 262961 95007 262989
rect 95041 262961 95069 262989
rect 95103 262961 95131 262989
rect 94917 254147 94945 254175
rect 94979 254147 95007 254175
rect 95041 254147 95069 254175
rect 95103 254147 95131 254175
rect 94917 254085 94945 254113
rect 94979 254085 95007 254113
rect 95041 254085 95069 254113
rect 95103 254085 95131 254113
rect 94917 254023 94945 254051
rect 94979 254023 95007 254051
rect 95041 254023 95069 254051
rect 95103 254023 95131 254051
rect 94917 253961 94945 253989
rect 94979 253961 95007 253989
rect 95041 253961 95069 253989
rect 95103 253961 95131 253989
rect 94917 245147 94945 245175
rect 94979 245147 95007 245175
rect 95041 245147 95069 245175
rect 95103 245147 95131 245175
rect 94917 245085 94945 245113
rect 94979 245085 95007 245113
rect 95041 245085 95069 245113
rect 95103 245085 95131 245113
rect 94917 245023 94945 245051
rect 94979 245023 95007 245051
rect 95041 245023 95069 245051
rect 95103 245023 95131 245051
rect 94917 244961 94945 244989
rect 94979 244961 95007 244989
rect 95041 244961 95069 244989
rect 95103 244961 95131 244989
rect 94917 236147 94945 236175
rect 94979 236147 95007 236175
rect 95041 236147 95069 236175
rect 95103 236147 95131 236175
rect 94917 236085 94945 236113
rect 94979 236085 95007 236113
rect 95041 236085 95069 236113
rect 95103 236085 95131 236113
rect 94917 236023 94945 236051
rect 94979 236023 95007 236051
rect 95041 236023 95069 236051
rect 95103 236023 95131 236051
rect 94917 235961 94945 235989
rect 94979 235961 95007 235989
rect 95041 235961 95069 235989
rect 95103 235961 95131 235989
rect 94917 227147 94945 227175
rect 94979 227147 95007 227175
rect 95041 227147 95069 227175
rect 95103 227147 95131 227175
rect 94917 227085 94945 227113
rect 94979 227085 95007 227113
rect 95041 227085 95069 227113
rect 95103 227085 95131 227113
rect 94917 227023 94945 227051
rect 94979 227023 95007 227051
rect 95041 227023 95069 227051
rect 95103 227023 95131 227051
rect 94917 226961 94945 226989
rect 94979 226961 95007 226989
rect 95041 226961 95069 226989
rect 95103 226961 95131 226989
rect 94917 218147 94945 218175
rect 94979 218147 95007 218175
rect 95041 218147 95069 218175
rect 95103 218147 95131 218175
rect 94917 218085 94945 218113
rect 94979 218085 95007 218113
rect 95041 218085 95069 218113
rect 95103 218085 95131 218113
rect 94917 218023 94945 218051
rect 94979 218023 95007 218051
rect 95041 218023 95069 218051
rect 95103 218023 95131 218051
rect 94917 217961 94945 217989
rect 94979 217961 95007 217989
rect 95041 217961 95069 217989
rect 95103 217961 95131 217989
rect 94917 209147 94945 209175
rect 94979 209147 95007 209175
rect 95041 209147 95069 209175
rect 95103 209147 95131 209175
rect 94917 209085 94945 209113
rect 94979 209085 95007 209113
rect 95041 209085 95069 209113
rect 95103 209085 95131 209113
rect 94917 209023 94945 209051
rect 94979 209023 95007 209051
rect 95041 209023 95069 209051
rect 95103 209023 95131 209051
rect 94917 208961 94945 208989
rect 94979 208961 95007 208989
rect 95041 208961 95069 208989
rect 95103 208961 95131 208989
rect 94917 200147 94945 200175
rect 94979 200147 95007 200175
rect 95041 200147 95069 200175
rect 95103 200147 95131 200175
rect 94917 200085 94945 200113
rect 94979 200085 95007 200113
rect 95041 200085 95069 200113
rect 95103 200085 95131 200113
rect 94917 200023 94945 200051
rect 94979 200023 95007 200051
rect 95041 200023 95069 200051
rect 95103 200023 95131 200051
rect 94917 199961 94945 199989
rect 94979 199961 95007 199989
rect 95041 199961 95069 199989
rect 95103 199961 95131 199989
rect 94917 191147 94945 191175
rect 94979 191147 95007 191175
rect 95041 191147 95069 191175
rect 95103 191147 95131 191175
rect 94917 191085 94945 191113
rect 94979 191085 95007 191113
rect 95041 191085 95069 191113
rect 95103 191085 95131 191113
rect 94917 191023 94945 191051
rect 94979 191023 95007 191051
rect 95041 191023 95069 191051
rect 95103 191023 95131 191051
rect 94917 190961 94945 190989
rect 94979 190961 95007 190989
rect 95041 190961 95069 190989
rect 95103 190961 95131 190989
rect 94917 182147 94945 182175
rect 94979 182147 95007 182175
rect 95041 182147 95069 182175
rect 95103 182147 95131 182175
rect 94917 182085 94945 182113
rect 94979 182085 95007 182113
rect 95041 182085 95069 182113
rect 95103 182085 95131 182113
rect 94917 182023 94945 182051
rect 94979 182023 95007 182051
rect 95041 182023 95069 182051
rect 95103 182023 95131 182051
rect 94917 181961 94945 181989
rect 94979 181961 95007 181989
rect 95041 181961 95069 181989
rect 95103 181961 95131 181989
rect 85059 173147 85087 173175
rect 85121 173147 85149 173175
rect 85059 173085 85087 173113
rect 85121 173085 85149 173113
rect 85059 173023 85087 173051
rect 85121 173023 85149 173051
rect 85059 172961 85087 172989
rect 85121 172961 85149 172989
rect 94917 173147 94945 173175
rect 94979 173147 95007 173175
rect 95041 173147 95069 173175
rect 95103 173147 95131 173175
rect 94917 173085 94945 173113
rect 94979 173085 95007 173113
rect 95041 173085 95069 173113
rect 95103 173085 95131 173113
rect 94917 173023 94945 173051
rect 94979 173023 95007 173051
rect 95041 173023 95069 173051
rect 95103 173023 95131 173051
rect 94917 172961 94945 172989
rect 94979 172961 95007 172989
rect 95041 172961 95069 172989
rect 95103 172961 95131 172989
rect 81417 167147 81445 167175
rect 81479 167147 81507 167175
rect 81541 167147 81569 167175
rect 81603 167147 81631 167175
rect 81417 167085 81445 167113
rect 81479 167085 81507 167113
rect 81541 167085 81569 167113
rect 81603 167085 81631 167113
rect 81417 167023 81445 167051
rect 81479 167023 81507 167051
rect 81541 167023 81569 167051
rect 81603 167023 81631 167051
rect 81417 166961 81445 166989
rect 81479 166961 81507 166989
rect 81541 166961 81569 166989
rect 81603 166961 81631 166989
rect 92739 167147 92767 167175
rect 92801 167147 92829 167175
rect 92739 167085 92767 167113
rect 92801 167085 92829 167113
rect 92739 167023 92767 167051
rect 92801 167023 92829 167051
rect 92739 166961 92767 166989
rect 92801 166961 92829 166989
rect 85059 164147 85087 164175
rect 85121 164147 85149 164175
rect 85059 164085 85087 164113
rect 85121 164085 85149 164113
rect 85059 164023 85087 164051
rect 85121 164023 85149 164051
rect 85059 163961 85087 163989
rect 85121 163961 85149 163989
rect 94917 164147 94945 164175
rect 94979 164147 95007 164175
rect 95041 164147 95069 164175
rect 95103 164147 95131 164175
rect 94917 164085 94945 164113
rect 94979 164085 95007 164113
rect 95041 164085 95069 164113
rect 95103 164085 95131 164113
rect 94917 164023 94945 164051
rect 94979 164023 95007 164051
rect 95041 164023 95069 164051
rect 95103 164023 95131 164051
rect 94917 163961 94945 163989
rect 94979 163961 95007 163989
rect 95041 163961 95069 163989
rect 95103 163961 95131 163989
rect 81417 158147 81445 158175
rect 81479 158147 81507 158175
rect 81541 158147 81569 158175
rect 81603 158147 81631 158175
rect 81417 158085 81445 158113
rect 81479 158085 81507 158113
rect 81541 158085 81569 158113
rect 81603 158085 81631 158113
rect 81417 158023 81445 158051
rect 81479 158023 81507 158051
rect 81541 158023 81569 158051
rect 81603 158023 81631 158051
rect 81417 157961 81445 157989
rect 81479 157961 81507 157989
rect 81541 157961 81569 157989
rect 81603 157961 81631 157989
rect 92739 158147 92767 158175
rect 92801 158147 92829 158175
rect 92739 158085 92767 158113
rect 92801 158085 92829 158113
rect 92739 158023 92767 158051
rect 92801 158023 92829 158051
rect 92739 157961 92767 157989
rect 92801 157961 92829 157989
rect 85059 155147 85087 155175
rect 85121 155147 85149 155175
rect 85059 155085 85087 155113
rect 85121 155085 85149 155113
rect 85059 155023 85087 155051
rect 85121 155023 85149 155051
rect 85059 154961 85087 154989
rect 85121 154961 85149 154989
rect 94917 155147 94945 155175
rect 94979 155147 95007 155175
rect 95041 155147 95069 155175
rect 95103 155147 95131 155175
rect 94917 155085 94945 155113
rect 94979 155085 95007 155113
rect 95041 155085 95069 155113
rect 95103 155085 95131 155113
rect 94917 155023 94945 155051
rect 94979 155023 95007 155051
rect 95041 155023 95069 155051
rect 95103 155023 95131 155051
rect 94917 154961 94945 154989
rect 94979 154961 95007 154989
rect 95041 154961 95069 154989
rect 95103 154961 95131 154989
rect 81417 149147 81445 149175
rect 81479 149147 81507 149175
rect 81541 149147 81569 149175
rect 81603 149147 81631 149175
rect 81417 149085 81445 149113
rect 81479 149085 81507 149113
rect 81541 149085 81569 149113
rect 81603 149085 81631 149113
rect 81417 149023 81445 149051
rect 81479 149023 81507 149051
rect 81541 149023 81569 149051
rect 81603 149023 81631 149051
rect 81417 148961 81445 148989
rect 81479 148961 81507 148989
rect 81541 148961 81569 148989
rect 81603 148961 81631 148989
rect 92739 149147 92767 149175
rect 92801 149147 92829 149175
rect 92739 149085 92767 149113
rect 92801 149085 92829 149113
rect 92739 149023 92767 149051
rect 92801 149023 92829 149051
rect 92739 148961 92767 148989
rect 92801 148961 92829 148989
rect 85059 146147 85087 146175
rect 85121 146147 85149 146175
rect 85059 146085 85087 146113
rect 85121 146085 85149 146113
rect 85059 146023 85087 146051
rect 85121 146023 85149 146051
rect 85059 145961 85087 145989
rect 85121 145961 85149 145989
rect 94917 146147 94945 146175
rect 94979 146147 95007 146175
rect 95041 146147 95069 146175
rect 95103 146147 95131 146175
rect 94917 146085 94945 146113
rect 94979 146085 95007 146113
rect 95041 146085 95069 146113
rect 95103 146085 95131 146113
rect 94917 146023 94945 146051
rect 94979 146023 95007 146051
rect 95041 146023 95069 146051
rect 95103 146023 95131 146051
rect 94917 145961 94945 145989
rect 94979 145961 95007 145989
rect 95041 145961 95069 145989
rect 95103 145961 95131 145989
rect 81417 140147 81445 140175
rect 81479 140147 81507 140175
rect 81541 140147 81569 140175
rect 81603 140147 81631 140175
rect 81417 140085 81445 140113
rect 81479 140085 81507 140113
rect 81541 140085 81569 140113
rect 81603 140085 81631 140113
rect 81417 140023 81445 140051
rect 81479 140023 81507 140051
rect 81541 140023 81569 140051
rect 81603 140023 81631 140051
rect 81417 139961 81445 139989
rect 81479 139961 81507 139989
rect 81541 139961 81569 139989
rect 81603 139961 81631 139989
rect 92739 140147 92767 140175
rect 92801 140147 92829 140175
rect 92739 140085 92767 140113
rect 92801 140085 92829 140113
rect 92739 140023 92767 140051
rect 92801 140023 92829 140051
rect 92739 139961 92767 139989
rect 92801 139961 92829 139989
rect 85059 137147 85087 137175
rect 85121 137147 85149 137175
rect 85059 137085 85087 137113
rect 85121 137085 85149 137113
rect 85059 137023 85087 137051
rect 85121 137023 85149 137051
rect 85059 136961 85087 136989
rect 85121 136961 85149 136989
rect 94917 137147 94945 137175
rect 94979 137147 95007 137175
rect 95041 137147 95069 137175
rect 95103 137147 95131 137175
rect 94917 137085 94945 137113
rect 94979 137085 95007 137113
rect 95041 137085 95069 137113
rect 95103 137085 95131 137113
rect 94917 137023 94945 137051
rect 94979 137023 95007 137051
rect 95041 137023 95069 137051
rect 95103 137023 95131 137051
rect 94917 136961 94945 136989
rect 94979 136961 95007 136989
rect 95041 136961 95069 136989
rect 95103 136961 95131 136989
rect 81417 131147 81445 131175
rect 81479 131147 81507 131175
rect 81541 131147 81569 131175
rect 81603 131147 81631 131175
rect 81417 131085 81445 131113
rect 81479 131085 81507 131113
rect 81541 131085 81569 131113
rect 81603 131085 81631 131113
rect 81417 131023 81445 131051
rect 81479 131023 81507 131051
rect 81541 131023 81569 131051
rect 81603 131023 81631 131051
rect 81417 130961 81445 130989
rect 81479 130961 81507 130989
rect 81541 130961 81569 130989
rect 81603 130961 81631 130989
rect 92739 131147 92767 131175
rect 92801 131147 92829 131175
rect 92739 131085 92767 131113
rect 92801 131085 92829 131113
rect 92739 131023 92767 131051
rect 92801 131023 92829 131051
rect 92739 130961 92767 130989
rect 92801 130961 92829 130989
rect 85059 128147 85087 128175
rect 85121 128147 85149 128175
rect 85059 128085 85087 128113
rect 85121 128085 85149 128113
rect 85059 128023 85087 128051
rect 85121 128023 85149 128051
rect 85059 127961 85087 127989
rect 85121 127961 85149 127989
rect 94917 128147 94945 128175
rect 94979 128147 95007 128175
rect 95041 128147 95069 128175
rect 95103 128147 95131 128175
rect 94917 128085 94945 128113
rect 94979 128085 95007 128113
rect 95041 128085 95069 128113
rect 95103 128085 95131 128113
rect 94917 128023 94945 128051
rect 94979 128023 95007 128051
rect 95041 128023 95069 128051
rect 95103 128023 95131 128051
rect 94917 127961 94945 127989
rect 94979 127961 95007 127989
rect 95041 127961 95069 127989
rect 95103 127961 95131 127989
rect 81417 122147 81445 122175
rect 81479 122147 81507 122175
rect 81541 122147 81569 122175
rect 81603 122147 81631 122175
rect 81417 122085 81445 122113
rect 81479 122085 81507 122113
rect 81541 122085 81569 122113
rect 81603 122085 81631 122113
rect 81417 122023 81445 122051
rect 81479 122023 81507 122051
rect 81541 122023 81569 122051
rect 81603 122023 81631 122051
rect 81417 121961 81445 121989
rect 81479 121961 81507 121989
rect 81541 121961 81569 121989
rect 81603 121961 81631 121989
rect 92739 122147 92767 122175
rect 92801 122147 92829 122175
rect 92739 122085 92767 122113
rect 92801 122085 92829 122113
rect 92739 122023 92767 122051
rect 92801 122023 92829 122051
rect 92739 121961 92767 121989
rect 92801 121961 92829 121989
rect 85059 119147 85087 119175
rect 85121 119147 85149 119175
rect 85059 119085 85087 119113
rect 85121 119085 85149 119113
rect 85059 119023 85087 119051
rect 85121 119023 85149 119051
rect 85059 118961 85087 118989
rect 85121 118961 85149 118989
rect 94917 119147 94945 119175
rect 94979 119147 95007 119175
rect 95041 119147 95069 119175
rect 95103 119147 95131 119175
rect 94917 119085 94945 119113
rect 94979 119085 95007 119113
rect 95041 119085 95069 119113
rect 95103 119085 95131 119113
rect 94917 119023 94945 119051
rect 94979 119023 95007 119051
rect 95041 119023 95069 119051
rect 95103 119023 95131 119051
rect 94917 118961 94945 118989
rect 94979 118961 95007 118989
rect 95041 118961 95069 118989
rect 95103 118961 95131 118989
rect 81417 113147 81445 113175
rect 81479 113147 81507 113175
rect 81541 113147 81569 113175
rect 81603 113147 81631 113175
rect 81417 113085 81445 113113
rect 81479 113085 81507 113113
rect 81541 113085 81569 113113
rect 81603 113085 81631 113113
rect 81417 113023 81445 113051
rect 81479 113023 81507 113051
rect 81541 113023 81569 113051
rect 81603 113023 81631 113051
rect 81417 112961 81445 112989
rect 81479 112961 81507 112989
rect 81541 112961 81569 112989
rect 81603 112961 81631 112989
rect 92739 113147 92767 113175
rect 92801 113147 92829 113175
rect 92739 113085 92767 113113
rect 92801 113085 92829 113113
rect 92739 113023 92767 113051
rect 92801 113023 92829 113051
rect 92739 112961 92767 112989
rect 92801 112961 92829 112989
rect 85059 110147 85087 110175
rect 85121 110147 85149 110175
rect 85059 110085 85087 110113
rect 85121 110085 85149 110113
rect 85059 110023 85087 110051
rect 85121 110023 85149 110051
rect 85059 109961 85087 109989
rect 85121 109961 85149 109989
rect 94917 110147 94945 110175
rect 94979 110147 95007 110175
rect 95041 110147 95069 110175
rect 95103 110147 95131 110175
rect 94917 110085 94945 110113
rect 94979 110085 95007 110113
rect 95041 110085 95069 110113
rect 95103 110085 95131 110113
rect 94917 110023 94945 110051
rect 94979 110023 95007 110051
rect 95041 110023 95069 110051
rect 95103 110023 95131 110051
rect 94917 109961 94945 109989
rect 94979 109961 95007 109989
rect 95041 109961 95069 109989
rect 95103 109961 95131 109989
rect 81417 104147 81445 104175
rect 81479 104147 81507 104175
rect 81541 104147 81569 104175
rect 81603 104147 81631 104175
rect 81417 104085 81445 104113
rect 81479 104085 81507 104113
rect 81541 104085 81569 104113
rect 81603 104085 81631 104113
rect 81417 104023 81445 104051
rect 81479 104023 81507 104051
rect 81541 104023 81569 104051
rect 81603 104023 81631 104051
rect 81417 103961 81445 103989
rect 81479 103961 81507 103989
rect 81541 103961 81569 103989
rect 81603 103961 81631 103989
rect 92739 104147 92767 104175
rect 92801 104147 92829 104175
rect 92739 104085 92767 104113
rect 92801 104085 92829 104113
rect 92739 104023 92767 104051
rect 92801 104023 92829 104051
rect 92739 103961 92767 103989
rect 92801 103961 92829 103989
rect 85059 101147 85087 101175
rect 85121 101147 85149 101175
rect 85059 101085 85087 101113
rect 85121 101085 85149 101113
rect 85059 101023 85087 101051
rect 85121 101023 85149 101051
rect 85059 100961 85087 100989
rect 85121 100961 85149 100989
rect 94917 101147 94945 101175
rect 94979 101147 95007 101175
rect 95041 101147 95069 101175
rect 95103 101147 95131 101175
rect 94917 101085 94945 101113
rect 94979 101085 95007 101113
rect 95041 101085 95069 101113
rect 95103 101085 95131 101113
rect 94917 101023 94945 101051
rect 94979 101023 95007 101051
rect 95041 101023 95069 101051
rect 95103 101023 95131 101051
rect 94917 100961 94945 100989
rect 94979 100961 95007 100989
rect 95041 100961 95069 100989
rect 95103 100961 95131 100989
rect 81417 95147 81445 95175
rect 81479 95147 81507 95175
rect 81541 95147 81569 95175
rect 81603 95147 81631 95175
rect 81417 95085 81445 95113
rect 81479 95085 81507 95113
rect 81541 95085 81569 95113
rect 81603 95085 81631 95113
rect 81417 95023 81445 95051
rect 81479 95023 81507 95051
rect 81541 95023 81569 95051
rect 81603 95023 81631 95051
rect 81417 94961 81445 94989
rect 81479 94961 81507 94989
rect 81541 94961 81569 94989
rect 81603 94961 81631 94989
rect 92739 95147 92767 95175
rect 92801 95147 92829 95175
rect 92739 95085 92767 95113
rect 92801 95085 92829 95113
rect 92739 95023 92767 95051
rect 92801 95023 92829 95051
rect 92739 94961 92767 94989
rect 92801 94961 92829 94989
rect 85059 92147 85087 92175
rect 85121 92147 85149 92175
rect 85059 92085 85087 92113
rect 85121 92085 85149 92113
rect 85059 92023 85087 92051
rect 85121 92023 85149 92051
rect 85059 91961 85087 91989
rect 85121 91961 85149 91989
rect 94917 92147 94945 92175
rect 94979 92147 95007 92175
rect 95041 92147 95069 92175
rect 95103 92147 95131 92175
rect 94917 92085 94945 92113
rect 94979 92085 95007 92113
rect 95041 92085 95069 92113
rect 95103 92085 95131 92113
rect 94917 92023 94945 92051
rect 94979 92023 95007 92051
rect 95041 92023 95069 92051
rect 95103 92023 95131 92051
rect 94917 91961 94945 91989
rect 94979 91961 95007 91989
rect 95041 91961 95069 91989
rect 95103 91961 95131 91989
rect 81417 86147 81445 86175
rect 81479 86147 81507 86175
rect 81541 86147 81569 86175
rect 81603 86147 81631 86175
rect 81417 86085 81445 86113
rect 81479 86085 81507 86113
rect 81541 86085 81569 86113
rect 81603 86085 81631 86113
rect 81417 86023 81445 86051
rect 81479 86023 81507 86051
rect 81541 86023 81569 86051
rect 81603 86023 81631 86051
rect 81417 85961 81445 85989
rect 81479 85961 81507 85989
rect 81541 85961 81569 85989
rect 81603 85961 81631 85989
rect 92739 86147 92767 86175
rect 92801 86147 92829 86175
rect 92739 86085 92767 86113
rect 92801 86085 92829 86113
rect 92739 86023 92767 86051
rect 92801 86023 92829 86051
rect 92739 85961 92767 85989
rect 92801 85961 92829 85989
rect 85059 83147 85087 83175
rect 85121 83147 85149 83175
rect 85059 83085 85087 83113
rect 85121 83085 85149 83113
rect 85059 83023 85087 83051
rect 85121 83023 85149 83051
rect 85059 82961 85087 82989
rect 85121 82961 85149 82989
rect 94917 83147 94945 83175
rect 94979 83147 95007 83175
rect 95041 83147 95069 83175
rect 95103 83147 95131 83175
rect 94917 83085 94945 83113
rect 94979 83085 95007 83113
rect 95041 83085 95069 83113
rect 95103 83085 95131 83113
rect 94917 83023 94945 83051
rect 94979 83023 95007 83051
rect 95041 83023 95069 83051
rect 95103 83023 95131 83051
rect 94917 82961 94945 82989
rect 94979 82961 95007 82989
rect 95041 82961 95069 82989
rect 95103 82961 95131 82989
rect 81417 77147 81445 77175
rect 81479 77147 81507 77175
rect 81541 77147 81569 77175
rect 81603 77147 81631 77175
rect 81417 77085 81445 77113
rect 81479 77085 81507 77113
rect 81541 77085 81569 77113
rect 81603 77085 81631 77113
rect 81417 77023 81445 77051
rect 81479 77023 81507 77051
rect 81541 77023 81569 77051
rect 81603 77023 81631 77051
rect 81417 76961 81445 76989
rect 81479 76961 81507 76989
rect 81541 76961 81569 76989
rect 81603 76961 81631 76989
rect 92739 77147 92767 77175
rect 92801 77147 92829 77175
rect 92739 77085 92767 77113
rect 92801 77085 92829 77113
rect 92739 77023 92767 77051
rect 92801 77023 92829 77051
rect 92739 76961 92767 76989
rect 92801 76961 92829 76989
rect 85059 74147 85087 74175
rect 85121 74147 85149 74175
rect 85059 74085 85087 74113
rect 85121 74085 85149 74113
rect 85059 74023 85087 74051
rect 85121 74023 85149 74051
rect 85059 73961 85087 73989
rect 85121 73961 85149 73989
rect 94917 74147 94945 74175
rect 94979 74147 95007 74175
rect 95041 74147 95069 74175
rect 95103 74147 95131 74175
rect 94917 74085 94945 74113
rect 94979 74085 95007 74113
rect 95041 74085 95069 74113
rect 95103 74085 95131 74113
rect 94917 74023 94945 74051
rect 94979 74023 95007 74051
rect 95041 74023 95069 74051
rect 95103 74023 95131 74051
rect 94917 73961 94945 73989
rect 94979 73961 95007 73989
rect 95041 73961 95069 73989
rect 95103 73961 95131 73989
rect 81417 68147 81445 68175
rect 81479 68147 81507 68175
rect 81541 68147 81569 68175
rect 81603 68147 81631 68175
rect 81417 68085 81445 68113
rect 81479 68085 81507 68113
rect 81541 68085 81569 68113
rect 81603 68085 81631 68113
rect 81417 68023 81445 68051
rect 81479 68023 81507 68051
rect 81541 68023 81569 68051
rect 81603 68023 81631 68051
rect 81417 67961 81445 67989
rect 81479 67961 81507 67989
rect 81541 67961 81569 67989
rect 81603 67961 81631 67989
rect 92739 68147 92767 68175
rect 92801 68147 92829 68175
rect 92739 68085 92767 68113
rect 92801 68085 92829 68113
rect 92739 68023 92767 68051
rect 92801 68023 92829 68051
rect 92739 67961 92767 67989
rect 92801 67961 92829 67989
rect 85059 65147 85087 65175
rect 85121 65147 85149 65175
rect 85059 65085 85087 65113
rect 85121 65085 85149 65113
rect 85059 65023 85087 65051
rect 85121 65023 85149 65051
rect 85059 64961 85087 64989
rect 85121 64961 85149 64989
rect 94917 65147 94945 65175
rect 94979 65147 95007 65175
rect 95041 65147 95069 65175
rect 95103 65147 95131 65175
rect 94917 65085 94945 65113
rect 94979 65085 95007 65113
rect 95041 65085 95069 65113
rect 95103 65085 95131 65113
rect 94917 65023 94945 65051
rect 94979 65023 95007 65051
rect 95041 65023 95069 65051
rect 95103 65023 95131 65051
rect 94917 64961 94945 64989
rect 94979 64961 95007 64989
rect 95041 64961 95069 64989
rect 95103 64961 95131 64989
rect 81417 59147 81445 59175
rect 81479 59147 81507 59175
rect 81541 59147 81569 59175
rect 81603 59147 81631 59175
rect 81417 59085 81445 59113
rect 81479 59085 81507 59113
rect 81541 59085 81569 59113
rect 81603 59085 81631 59113
rect 81417 59023 81445 59051
rect 81479 59023 81507 59051
rect 81541 59023 81569 59051
rect 81603 59023 81631 59051
rect 81417 58961 81445 58989
rect 81479 58961 81507 58989
rect 81541 58961 81569 58989
rect 81603 58961 81631 58989
rect 92739 59147 92767 59175
rect 92801 59147 92829 59175
rect 92739 59085 92767 59113
rect 92801 59085 92829 59113
rect 92739 59023 92767 59051
rect 92801 59023 92829 59051
rect 92739 58961 92767 58989
rect 92801 58961 92829 58989
rect 85059 56147 85087 56175
rect 85121 56147 85149 56175
rect 85059 56085 85087 56113
rect 85121 56085 85149 56113
rect 85059 56023 85087 56051
rect 85121 56023 85149 56051
rect 85059 55961 85087 55989
rect 85121 55961 85149 55989
rect 94917 56147 94945 56175
rect 94979 56147 95007 56175
rect 95041 56147 95069 56175
rect 95103 56147 95131 56175
rect 94917 56085 94945 56113
rect 94979 56085 95007 56113
rect 95041 56085 95069 56113
rect 95103 56085 95131 56113
rect 94917 56023 94945 56051
rect 94979 56023 95007 56051
rect 95041 56023 95069 56051
rect 95103 56023 95131 56051
rect 94917 55961 94945 55989
rect 94979 55961 95007 55989
rect 95041 55961 95069 55989
rect 95103 55961 95131 55989
rect 81417 50147 81445 50175
rect 81479 50147 81507 50175
rect 81541 50147 81569 50175
rect 81603 50147 81631 50175
rect 81417 50085 81445 50113
rect 81479 50085 81507 50113
rect 81541 50085 81569 50113
rect 81603 50085 81631 50113
rect 81417 50023 81445 50051
rect 81479 50023 81507 50051
rect 81541 50023 81569 50051
rect 81603 50023 81631 50051
rect 81417 49961 81445 49989
rect 81479 49961 81507 49989
rect 81541 49961 81569 49989
rect 81603 49961 81631 49989
rect 92739 50147 92767 50175
rect 92801 50147 92829 50175
rect 92739 50085 92767 50113
rect 92801 50085 92829 50113
rect 92739 50023 92767 50051
rect 92801 50023 92829 50051
rect 92739 49961 92767 49989
rect 92801 49961 92829 49989
rect 85059 47147 85087 47175
rect 85121 47147 85149 47175
rect 85059 47085 85087 47113
rect 85121 47085 85149 47113
rect 85059 47023 85087 47051
rect 85121 47023 85149 47051
rect 85059 46961 85087 46989
rect 85121 46961 85149 46989
rect 94917 47147 94945 47175
rect 94979 47147 95007 47175
rect 95041 47147 95069 47175
rect 95103 47147 95131 47175
rect 94917 47085 94945 47113
rect 94979 47085 95007 47113
rect 95041 47085 95069 47113
rect 95103 47085 95131 47113
rect 94917 47023 94945 47051
rect 94979 47023 95007 47051
rect 95041 47023 95069 47051
rect 95103 47023 95131 47051
rect 94917 46961 94945 46989
rect 94979 46961 95007 46989
rect 95041 46961 95069 46989
rect 95103 46961 95131 46989
rect 81417 41147 81445 41175
rect 81479 41147 81507 41175
rect 81541 41147 81569 41175
rect 81603 41147 81631 41175
rect 81417 41085 81445 41113
rect 81479 41085 81507 41113
rect 81541 41085 81569 41113
rect 81603 41085 81631 41113
rect 81417 41023 81445 41051
rect 81479 41023 81507 41051
rect 81541 41023 81569 41051
rect 81603 41023 81631 41051
rect 81417 40961 81445 40989
rect 81479 40961 81507 40989
rect 81541 40961 81569 40989
rect 81603 40961 81631 40989
rect 92739 41147 92767 41175
rect 92801 41147 92829 41175
rect 92739 41085 92767 41113
rect 92801 41085 92829 41113
rect 92739 41023 92767 41051
rect 92801 41023 92829 41051
rect 92739 40961 92767 40989
rect 92801 40961 92829 40989
rect 85059 38147 85087 38175
rect 85121 38147 85149 38175
rect 85059 38085 85087 38113
rect 85121 38085 85149 38113
rect 85059 38023 85087 38051
rect 85121 38023 85149 38051
rect 85059 37961 85087 37989
rect 85121 37961 85149 37989
rect 94917 38147 94945 38175
rect 94979 38147 95007 38175
rect 95041 38147 95069 38175
rect 95103 38147 95131 38175
rect 94917 38085 94945 38113
rect 94979 38085 95007 38113
rect 95041 38085 95069 38113
rect 95103 38085 95131 38113
rect 94917 38023 94945 38051
rect 94979 38023 95007 38051
rect 95041 38023 95069 38051
rect 95103 38023 95131 38051
rect 94917 37961 94945 37989
rect 94979 37961 95007 37989
rect 95041 37961 95069 37989
rect 95103 37961 95131 37989
rect 81417 32147 81445 32175
rect 81479 32147 81507 32175
rect 81541 32147 81569 32175
rect 81603 32147 81631 32175
rect 81417 32085 81445 32113
rect 81479 32085 81507 32113
rect 81541 32085 81569 32113
rect 81603 32085 81631 32113
rect 81417 32023 81445 32051
rect 81479 32023 81507 32051
rect 81541 32023 81569 32051
rect 81603 32023 81631 32051
rect 81417 31961 81445 31989
rect 81479 31961 81507 31989
rect 81541 31961 81569 31989
rect 81603 31961 81631 31989
rect 92739 32147 92767 32175
rect 92801 32147 92829 32175
rect 92739 32085 92767 32113
rect 92801 32085 92829 32113
rect 92739 32023 92767 32051
rect 92801 32023 92829 32051
rect 92739 31961 92767 31989
rect 92801 31961 92829 31989
rect 85059 29147 85087 29175
rect 85121 29147 85149 29175
rect 85059 29085 85087 29113
rect 85121 29085 85149 29113
rect 85059 29023 85087 29051
rect 85121 29023 85149 29051
rect 85059 28961 85087 28989
rect 85121 28961 85149 28989
rect 94917 29147 94945 29175
rect 94979 29147 95007 29175
rect 95041 29147 95069 29175
rect 95103 29147 95131 29175
rect 94917 29085 94945 29113
rect 94979 29085 95007 29113
rect 95041 29085 95069 29113
rect 95103 29085 95131 29113
rect 94917 29023 94945 29051
rect 94979 29023 95007 29051
rect 95041 29023 95069 29051
rect 95103 29023 95131 29051
rect 94917 28961 94945 28989
rect 94979 28961 95007 28989
rect 95041 28961 95069 28989
rect 95103 28961 95131 28989
rect 81417 23147 81445 23175
rect 81479 23147 81507 23175
rect 81541 23147 81569 23175
rect 81603 23147 81631 23175
rect 81417 23085 81445 23113
rect 81479 23085 81507 23113
rect 81541 23085 81569 23113
rect 81603 23085 81631 23113
rect 81417 23023 81445 23051
rect 81479 23023 81507 23051
rect 81541 23023 81569 23051
rect 81603 23023 81631 23051
rect 81417 22961 81445 22989
rect 81479 22961 81507 22989
rect 81541 22961 81569 22989
rect 81603 22961 81631 22989
rect 92739 23147 92767 23175
rect 92801 23147 92829 23175
rect 92739 23085 92767 23113
rect 92801 23085 92829 23113
rect 92739 23023 92767 23051
rect 92801 23023 92829 23051
rect 92739 22961 92767 22989
rect 92801 22961 92829 22989
rect 85059 20147 85087 20175
rect 85121 20147 85149 20175
rect 85059 20085 85087 20113
rect 85121 20085 85149 20113
rect 85059 20023 85087 20051
rect 85121 20023 85149 20051
rect 85059 19961 85087 19989
rect 85121 19961 85149 19989
rect 94917 20147 94945 20175
rect 94979 20147 95007 20175
rect 95041 20147 95069 20175
rect 95103 20147 95131 20175
rect 94917 20085 94945 20113
rect 94979 20085 95007 20113
rect 95041 20085 95069 20113
rect 95103 20085 95131 20113
rect 94917 20023 94945 20051
rect 94979 20023 95007 20051
rect 95041 20023 95069 20051
rect 95103 20023 95131 20051
rect 94917 19961 94945 19989
rect 94979 19961 95007 19989
rect 95041 19961 95069 19989
rect 95103 19961 95131 19989
rect 81417 14147 81445 14175
rect 81479 14147 81507 14175
rect 81541 14147 81569 14175
rect 81603 14147 81631 14175
rect 81417 14085 81445 14113
rect 81479 14085 81507 14113
rect 81541 14085 81569 14113
rect 81603 14085 81631 14113
rect 81417 14023 81445 14051
rect 81479 14023 81507 14051
rect 81541 14023 81569 14051
rect 81603 14023 81631 14051
rect 81417 13961 81445 13989
rect 81479 13961 81507 13989
rect 81541 13961 81569 13989
rect 81603 13961 81631 13989
rect 92739 14147 92767 14175
rect 92801 14147 92829 14175
rect 92739 14085 92767 14113
rect 92801 14085 92829 14113
rect 92739 14023 92767 14051
rect 92801 14023 92829 14051
rect 92739 13961 92767 13989
rect 92801 13961 92829 13989
rect 85059 11147 85087 11175
rect 85121 11147 85149 11175
rect 85059 11085 85087 11113
rect 85121 11085 85149 11113
rect 85059 11023 85087 11051
rect 85121 11023 85149 11051
rect 85059 10961 85087 10989
rect 85121 10961 85149 10989
rect 94917 11147 94945 11175
rect 94979 11147 95007 11175
rect 95041 11147 95069 11175
rect 95103 11147 95131 11175
rect 94917 11085 94945 11113
rect 94979 11085 95007 11113
rect 95041 11085 95069 11113
rect 95103 11085 95131 11113
rect 94917 11023 94945 11051
rect 94979 11023 95007 11051
rect 95041 11023 95069 11051
rect 95103 11023 95131 11051
rect 94917 10961 94945 10989
rect 94979 10961 95007 10989
rect 95041 10961 95069 10989
rect 95103 10961 95131 10989
rect 81417 5147 81445 5175
rect 81479 5147 81507 5175
rect 81541 5147 81569 5175
rect 81603 5147 81631 5175
rect 81417 5085 81445 5113
rect 81479 5085 81507 5113
rect 81541 5085 81569 5113
rect 81603 5085 81631 5113
rect 81417 5023 81445 5051
rect 81479 5023 81507 5051
rect 81541 5023 81569 5051
rect 81603 5023 81631 5051
rect 81417 4961 81445 4989
rect 81479 4961 81507 4989
rect 81541 4961 81569 4989
rect 81603 4961 81631 4989
rect 92739 5147 92767 5175
rect 92801 5147 92829 5175
rect 92739 5085 92767 5113
rect 92801 5085 92829 5113
rect 92739 5023 92767 5051
rect 92801 5023 92829 5051
rect 92739 4961 92767 4989
rect 92801 4961 92829 4989
rect 81417 -588 81445 -560
rect 81479 -588 81507 -560
rect 81541 -588 81569 -560
rect 81603 -588 81631 -560
rect 81417 -650 81445 -622
rect 81479 -650 81507 -622
rect 81541 -650 81569 -622
rect 81603 -650 81631 -622
rect 81417 -712 81445 -684
rect 81479 -712 81507 -684
rect 81541 -712 81569 -684
rect 81603 -712 81631 -684
rect 81417 -774 81445 -746
rect 81479 -774 81507 -746
rect 81541 -774 81569 -746
rect 81603 -774 81631 -746
rect 94917 2147 94945 2175
rect 94979 2147 95007 2175
rect 95041 2147 95069 2175
rect 95103 2147 95131 2175
rect 94917 2085 94945 2113
rect 94979 2085 95007 2113
rect 95041 2085 95069 2113
rect 95103 2085 95131 2113
rect 94917 2023 94945 2051
rect 94979 2023 95007 2051
rect 95041 2023 95069 2051
rect 95103 2023 95131 2051
rect 94917 1961 94945 1989
rect 94979 1961 95007 1989
rect 95041 1961 95069 1989
rect 95103 1961 95131 1989
rect 94917 -108 94945 -80
rect 94979 -108 95007 -80
rect 95041 -108 95069 -80
rect 95103 -108 95131 -80
rect 94917 -170 94945 -142
rect 94979 -170 95007 -142
rect 95041 -170 95069 -142
rect 95103 -170 95131 -142
rect 94917 -232 94945 -204
rect 94979 -232 95007 -204
rect 95041 -232 95069 -204
rect 95103 -232 95131 -204
rect 94917 -294 94945 -266
rect 94979 -294 95007 -266
rect 95041 -294 95069 -266
rect 95103 -294 95131 -266
rect 96777 299058 96805 299086
rect 96839 299058 96867 299086
rect 96901 299058 96929 299086
rect 96963 299058 96991 299086
rect 96777 298996 96805 299024
rect 96839 298996 96867 299024
rect 96901 298996 96929 299024
rect 96963 298996 96991 299024
rect 96777 298934 96805 298962
rect 96839 298934 96867 298962
rect 96901 298934 96929 298962
rect 96963 298934 96991 298962
rect 96777 298872 96805 298900
rect 96839 298872 96867 298900
rect 96901 298872 96929 298900
rect 96963 298872 96991 298900
rect 96777 293147 96805 293175
rect 96839 293147 96867 293175
rect 96901 293147 96929 293175
rect 96963 293147 96991 293175
rect 96777 293085 96805 293113
rect 96839 293085 96867 293113
rect 96901 293085 96929 293113
rect 96963 293085 96991 293113
rect 96777 293023 96805 293051
rect 96839 293023 96867 293051
rect 96901 293023 96929 293051
rect 96963 293023 96991 293051
rect 96777 292961 96805 292989
rect 96839 292961 96867 292989
rect 96901 292961 96929 292989
rect 96963 292961 96991 292989
rect 96777 284147 96805 284175
rect 96839 284147 96867 284175
rect 96901 284147 96929 284175
rect 96963 284147 96991 284175
rect 96777 284085 96805 284113
rect 96839 284085 96867 284113
rect 96901 284085 96929 284113
rect 96963 284085 96991 284113
rect 96777 284023 96805 284051
rect 96839 284023 96867 284051
rect 96901 284023 96929 284051
rect 96963 284023 96991 284051
rect 96777 283961 96805 283989
rect 96839 283961 96867 283989
rect 96901 283961 96929 283989
rect 96963 283961 96991 283989
rect 96777 275147 96805 275175
rect 96839 275147 96867 275175
rect 96901 275147 96929 275175
rect 96963 275147 96991 275175
rect 96777 275085 96805 275113
rect 96839 275085 96867 275113
rect 96901 275085 96929 275113
rect 96963 275085 96991 275113
rect 96777 275023 96805 275051
rect 96839 275023 96867 275051
rect 96901 275023 96929 275051
rect 96963 275023 96991 275051
rect 96777 274961 96805 274989
rect 96839 274961 96867 274989
rect 96901 274961 96929 274989
rect 96963 274961 96991 274989
rect 96777 266147 96805 266175
rect 96839 266147 96867 266175
rect 96901 266147 96929 266175
rect 96963 266147 96991 266175
rect 96777 266085 96805 266113
rect 96839 266085 96867 266113
rect 96901 266085 96929 266113
rect 96963 266085 96991 266113
rect 96777 266023 96805 266051
rect 96839 266023 96867 266051
rect 96901 266023 96929 266051
rect 96963 266023 96991 266051
rect 96777 265961 96805 265989
rect 96839 265961 96867 265989
rect 96901 265961 96929 265989
rect 96963 265961 96991 265989
rect 96777 257147 96805 257175
rect 96839 257147 96867 257175
rect 96901 257147 96929 257175
rect 96963 257147 96991 257175
rect 96777 257085 96805 257113
rect 96839 257085 96867 257113
rect 96901 257085 96929 257113
rect 96963 257085 96991 257113
rect 96777 257023 96805 257051
rect 96839 257023 96867 257051
rect 96901 257023 96929 257051
rect 96963 257023 96991 257051
rect 96777 256961 96805 256989
rect 96839 256961 96867 256989
rect 96901 256961 96929 256989
rect 96963 256961 96991 256989
rect 96777 248147 96805 248175
rect 96839 248147 96867 248175
rect 96901 248147 96929 248175
rect 96963 248147 96991 248175
rect 96777 248085 96805 248113
rect 96839 248085 96867 248113
rect 96901 248085 96929 248113
rect 96963 248085 96991 248113
rect 96777 248023 96805 248051
rect 96839 248023 96867 248051
rect 96901 248023 96929 248051
rect 96963 248023 96991 248051
rect 96777 247961 96805 247989
rect 96839 247961 96867 247989
rect 96901 247961 96929 247989
rect 96963 247961 96991 247989
rect 96777 239147 96805 239175
rect 96839 239147 96867 239175
rect 96901 239147 96929 239175
rect 96963 239147 96991 239175
rect 96777 239085 96805 239113
rect 96839 239085 96867 239113
rect 96901 239085 96929 239113
rect 96963 239085 96991 239113
rect 96777 239023 96805 239051
rect 96839 239023 96867 239051
rect 96901 239023 96929 239051
rect 96963 239023 96991 239051
rect 96777 238961 96805 238989
rect 96839 238961 96867 238989
rect 96901 238961 96929 238989
rect 96963 238961 96991 238989
rect 96777 230147 96805 230175
rect 96839 230147 96867 230175
rect 96901 230147 96929 230175
rect 96963 230147 96991 230175
rect 96777 230085 96805 230113
rect 96839 230085 96867 230113
rect 96901 230085 96929 230113
rect 96963 230085 96991 230113
rect 96777 230023 96805 230051
rect 96839 230023 96867 230051
rect 96901 230023 96929 230051
rect 96963 230023 96991 230051
rect 96777 229961 96805 229989
rect 96839 229961 96867 229989
rect 96901 229961 96929 229989
rect 96963 229961 96991 229989
rect 96777 221147 96805 221175
rect 96839 221147 96867 221175
rect 96901 221147 96929 221175
rect 96963 221147 96991 221175
rect 96777 221085 96805 221113
rect 96839 221085 96867 221113
rect 96901 221085 96929 221113
rect 96963 221085 96991 221113
rect 96777 221023 96805 221051
rect 96839 221023 96867 221051
rect 96901 221023 96929 221051
rect 96963 221023 96991 221051
rect 96777 220961 96805 220989
rect 96839 220961 96867 220989
rect 96901 220961 96929 220989
rect 96963 220961 96991 220989
rect 96777 212147 96805 212175
rect 96839 212147 96867 212175
rect 96901 212147 96929 212175
rect 96963 212147 96991 212175
rect 96777 212085 96805 212113
rect 96839 212085 96867 212113
rect 96901 212085 96929 212113
rect 96963 212085 96991 212113
rect 96777 212023 96805 212051
rect 96839 212023 96867 212051
rect 96901 212023 96929 212051
rect 96963 212023 96991 212051
rect 96777 211961 96805 211989
rect 96839 211961 96867 211989
rect 96901 211961 96929 211989
rect 96963 211961 96991 211989
rect 96777 203147 96805 203175
rect 96839 203147 96867 203175
rect 96901 203147 96929 203175
rect 96963 203147 96991 203175
rect 96777 203085 96805 203113
rect 96839 203085 96867 203113
rect 96901 203085 96929 203113
rect 96963 203085 96991 203113
rect 96777 203023 96805 203051
rect 96839 203023 96867 203051
rect 96901 203023 96929 203051
rect 96963 203023 96991 203051
rect 96777 202961 96805 202989
rect 96839 202961 96867 202989
rect 96901 202961 96929 202989
rect 96963 202961 96991 202989
rect 96777 194147 96805 194175
rect 96839 194147 96867 194175
rect 96901 194147 96929 194175
rect 96963 194147 96991 194175
rect 96777 194085 96805 194113
rect 96839 194085 96867 194113
rect 96901 194085 96929 194113
rect 96963 194085 96991 194113
rect 96777 194023 96805 194051
rect 96839 194023 96867 194051
rect 96901 194023 96929 194051
rect 96963 194023 96991 194051
rect 96777 193961 96805 193989
rect 96839 193961 96867 193989
rect 96901 193961 96929 193989
rect 96963 193961 96991 193989
rect 96777 185147 96805 185175
rect 96839 185147 96867 185175
rect 96901 185147 96929 185175
rect 96963 185147 96991 185175
rect 96777 185085 96805 185113
rect 96839 185085 96867 185113
rect 96901 185085 96929 185113
rect 96963 185085 96991 185113
rect 96777 185023 96805 185051
rect 96839 185023 96867 185051
rect 96901 185023 96929 185051
rect 96963 185023 96991 185051
rect 96777 184961 96805 184989
rect 96839 184961 96867 184989
rect 96901 184961 96929 184989
rect 96963 184961 96991 184989
rect 96777 176147 96805 176175
rect 96839 176147 96867 176175
rect 96901 176147 96929 176175
rect 96963 176147 96991 176175
rect 96777 176085 96805 176113
rect 96839 176085 96867 176113
rect 96901 176085 96929 176113
rect 96963 176085 96991 176113
rect 96777 176023 96805 176051
rect 96839 176023 96867 176051
rect 96901 176023 96929 176051
rect 96963 176023 96991 176051
rect 96777 175961 96805 175989
rect 96839 175961 96867 175989
rect 96901 175961 96929 175989
rect 96963 175961 96991 175989
rect 110277 298578 110305 298606
rect 110339 298578 110367 298606
rect 110401 298578 110429 298606
rect 110463 298578 110491 298606
rect 110277 298516 110305 298544
rect 110339 298516 110367 298544
rect 110401 298516 110429 298544
rect 110463 298516 110491 298544
rect 110277 298454 110305 298482
rect 110339 298454 110367 298482
rect 110401 298454 110429 298482
rect 110463 298454 110491 298482
rect 110277 298392 110305 298420
rect 110339 298392 110367 298420
rect 110401 298392 110429 298420
rect 110463 298392 110491 298420
rect 110277 290147 110305 290175
rect 110339 290147 110367 290175
rect 110401 290147 110429 290175
rect 110463 290147 110491 290175
rect 110277 290085 110305 290113
rect 110339 290085 110367 290113
rect 110401 290085 110429 290113
rect 110463 290085 110491 290113
rect 110277 290023 110305 290051
rect 110339 290023 110367 290051
rect 110401 290023 110429 290051
rect 110463 290023 110491 290051
rect 110277 289961 110305 289989
rect 110339 289961 110367 289989
rect 110401 289961 110429 289989
rect 110463 289961 110491 289989
rect 110277 281147 110305 281175
rect 110339 281147 110367 281175
rect 110401 281147 110429 281175
rect 110463 281147 110491 281175
rect 110277 281085 110305 281113
rect 110339 281085 110367 281113
rect 110401 281085 110429 281113
rect 110463 281085 110491 281113
rect 110277 281023 110305 281051
rect 110339 281023 110367 281051
rect 110401 281023 110429 281051
rect 110463 281023 110491 281051
rect 110277 280961 110305 280989
rect 110339 280961 110367 280989
rect 110401 280961 110429 280989
rect 110463 280961 110491 280989
rect 110277 272147 110305 272175
rect 110339 272147 110367 272175
rect 110401 272147 110429 272175
rect 110463 272147 110491 272175
rect 110277 272085 110305 272113
rect 110339 272085 110367 272113
rect 110401 272085 110429 272113
rect 110463 272085 110491 272113
rect 110277 272023 110305 272051
rect 110339 272023 110367 272051
rect 110401 272023 110429 272051
rect 110463 272023 110491 272051
rect 110277 271961 110305 271989
rect 110339 271961 110367 271989
rect 110401 271961 110429 271989
rect 110463 271961 110491 271989
rect 110277 263147 110305 263175
rect 110339 263147 110367 263175
rect 110401 263147 110429 263175
rect 110463 263147 110491 263175
rect 110277 263085 110305 263113
rect 110339 263085 110367 263113
rect 110401 263085 110429 263113
rect 110463 263085 110491 263113
rect 110277 263023 110305 263051
rect 110339 263023 110367 263051
rect 110401 263023 110429 263051
rect 110463 263023 110491 263051
rect 110277 262961 110305 262989
rect 110339 262961 110367 262989
rect 110401 262961 110429 262989
rect 110463 262961 110491 262989
rect 110277 254147 110305 254175
rect 110339 254147 110367 254175
rect 110401 254147 110429 254175
rect 110463 254147 110491 254175
rect 110277 254085 110305 254113
rect 110339 254085 110367 254113
rect 110401 254085 110429 254113
rect 110463 254085 110491 254113
rect 110277 254023 110305 254051
rect 110339 254023 110367 254051
rect 110401 254023 110429 254051
rect 110463 254023 110491 254051
rect 110277 253961 110305 253989
rect 110339 253961 110367 253989
rect 110401 253961 110429 253989
rect 110463 253961 110491 253989
rect 110277 245147 110305 245175
rect 110339 245147 110367 245175
rect 110401 245147 110429 245175
rect 110463 245147 110491 245175
rect 110277 245085 110305 245113
rect 110339 245085 110367 245113
rect 110401 245085 110429 245113
rect 110463 245085 110491 245113
rect 110277 245023 110305 245051
rect 110339 245023 110367 245051
rect 110401 245023 110429 245051
rect 110463 245023 110491 245051
rect 110277 244961 110305 244989
rect 110339 244961 110367 244989
rect 110401 244961 110429 244989
rect 110463 244961 110491 244989
rect 110277 236147 110305 236175
rect 110339 236147 110367 236175
rect 110401 236147 110429 236175
rect 110463 236147 110491 236175
rect 110277 236085 110305 236113
rect 110339 236085 110367 236113
rect 110401 236085 110429 236113
rect 110463 236085 110491 236113
rect 110277 236023 110305 236051
rect 110339 236023 110367 236051
rect 110401 236023 110429 236051
rect 110463 236023 110491 236051
rect 110277 235961 110305 235989
rect 110339 235961 110367 235989
rect 110401 235961 110429 235989
rect 110463 235961 110491 235989
rect 110277 227147 110305 227175
rect 110339 227147 110367 227175
rect 110401 227147 110429 227175
rect 110463 227147 110491 227175
rect 110277 227085 110305 227113
rect 110339 227085 110367 227113
rect 110401 227085 110429 227113
rect 110463 227085 110491 227113
rect 110277 227023 110305 227051
rect 110339 227023 110367 227051
rect 110401 227023 110429 227051
rect 110463 227023 110491 227051
rect 110277 226961 110305 226989
rect 110339 226961 110367 226989
rect 110401 226961 110429 226989
rect 110463 226961 110491 226989
rect 110277 218147 110305 218175
rect 110339 218147 110367 218175
rect 110401 218147 110429 218175
rect 110463 218147 110491 218175
rect 110277 218085 110305 218113
rect 110339 218085 110367 218113
rect 110401 218085 110429 218113
rect 110463 218085 110491 218113
rect 110277 218023 110305 218051
rect 110339 218023 110367 218051
rect 110401 218023 110429 218051
rect 110463 218023 110491 218051
rect 110277 217961 110305 217989
rect 110339 217961 110367 217989
rect 110401 217961 110429 217989
rect 110463 217961 110491 217989
rect 110277 209147 110305 209175
rect 110339 209147 110367 209175
rect 110401 209147 110429 209175
rect 110463 209147 110491 209175
rect 110277 209085 110305 209113
rect 110339 209085 110367 209113
rect 110401 209085 110429 209113
rect 110463 209085 110491 209113
rect 110277 209023 110305 209051
rect 110339 209023 110367 209051
rect 110401 209023 110429 209051
rect 110463 209023 110491 209051
rect 110277 208961 110305 208989
rect 110339 208961 110367 208989
rect 110401 208961 110429 208989
rect 110463 208961 110491 208989
rect 110277 200147 110305 200175
rect 110339 200147 110367 200175
rect 110401 200147 110429 200175
rect 110463 200147 110491 200175
rect 110277 200085 110305 200113
rect 110339 200085 110367 200113
rect 110401 200085 110429 200113
rect 110463 200085 110491 200113
rect 110277 200023 110305 200051
rect 110339 200023 110367 200051
rect 110401 200023 110429 200051
rect 110463 200023 110491 200051
rect 110277 199961 110305 199989
rect 110339 199961 110367 199989
rect 110401 199961 110429 199989
rect 110463 199961 110491 199989
rect 110277 191147 110305 191175
rect 110339 191147 110367 191175
rect 110401 191147 110429 191175
rect 110463 191147 110491 191175
rect 110277 191085 110305 191113
rect 110339 191085 110367 191113
rect 110401 191085 110429 191113
rect 110463 191085 110491 191113
rect 110277 191023 110305 191051
rect 110339 191023 110367 191051
rect 110401 191023 110429 191051
rect 110463 191023 110491 191051
rect 110277 190961 110305 190989
rect 110339 190961 110367 190989
rect 110401 190961 110429 190989
rect 110463 190961 110491 190989
rect 110277 182147 110305 182175
rect 110339 182147 110367 182175
rect 110401 182147 110429 182175
rect 110463 182147 110491 182175
rect 110277 182085 110305 182113
rect 110339 182085 110367 182113
rect 110401 182085 110429 182113
rect 110463 182085 110491 182113
rect 110277 182023 110305 182051
rect 110339 182023 110367 182051
rect 110401 182023 110429 182051
rect 110463 182023 110491 182051
rect 110277 181961 110305 181989
rect 110339 181961 110367 181989
rect 110401 181961 110429 181989
rect 110463 181961 110491 181989
rect 100419 173147 100447 173175
rect 100481 173147 100509 173175
rect 100419 173085 100447 173113
rect 100481 173085 100509 173113
rect 100419 173023 100447 173051
rect 100481 173023 100509 173051
rect 100419 172961 100447 172989
rect 100481 172961 100509 172989
rect 110277 173147 110305 173175
rect 110339 173147 110367 173175
rect 110401 173147 110429 173175
rect 110463 173147 110491 173175
rect 110277 173085 110305 173113
rect 110339 173085 110367 173113
rect 110401 173085 110429 173113
rect 110463 173085 110491 173113
rect 110277 173023 110305 173051
rect 110339 173023 110367 173051
rect 110401 173023 110429 173051
rect 110463 173023 110491 173051
rect 110277 172961 110305 172989
rect 110339 172961 110367 172989
rect 110401 172961 110429 172989
rect 110463 172961 110491 172989
rect 96777 167147 96805 167175
rect 96839 167147 96867 167175
rect 96901 167147 96929 167175
rect 96963 167147 96991 167175
rect 96777 167085 96805 167113
rect 96839 167085 96867 167113
rect 96901 167085 96929 167113
rect 96963 167085 96991 167113
rect 96777 167023 96805 167051
rect 96839 167023 96867 167051
rect 96901 167023 96929 167051
rect 96963 167023 96991 167051
rect 96777 166961 96805 166989
rect 96839 166961 96867 166989
rect 96901 166961 96929 166989
rect 96963 166961 96991 166989
rect 108099 167147 108127 167175
rect 108161 167147 108189 167175
rect 108099 167085 108127 167113
rect 108161 167085 108189 167113
rect 108099 167023 108127 167051
rect 108161 167023 108189 167051
rect 108099 166961 108127 166989
rect 108161 166961 108189 166989
rect 100419 164147 100447 164175
rect 100481 164147 100509 164175
rect 100419 164085 100447 164113
rect 100481 164085 100509 164113
rect 100419 164023 100447 164051
rect 100481 164023 100509 164051
rect 100419 163961 100447 163989
rect 100481 163961 100509 163989
rect 110277 164147 110305 164175
rect 110339 164147 110367 164175
rect 110401 164147 110429 164175
rect 110463 164147 110491 164175
rect 110277 164085 110305 164113
rect 110339 164085 110367 164113
rect 110401 164085 110429 164113
rect 110463 164085 110491 164113
rect 110277 164023 110305 164051
rect 110339 164023 110367 164051
rect 110401 164023 110429 164051
rect 110463 164023 110491 164051
rect 110277 163961 110305 163989
rect 110339 163961 110367 163989
rect 110401 163961 110429 163989
rect 110463 163961 110491 163989
rect 96777 158147 96805 158175
rect 96839 158147 96867 158175
rect 96901 158147 96929 158175
rect 96963 158147 96991 158175
rect 96777 158085 96805 158113
rect 96839 158085 96867 158113
rect 96901 158085 96929 158113
rect 96963 158085 96991 158113
rect 96777 158023 96805 158051
rect 96839 158023 96867 158051
rect 96901 158023 96929 158051
rect 96963 158023 96991 158051
rect 96777 157961 96805 157989
rect 96839 157961 96867 157989
rect 96901 157961 96929 157989
rect 96963 157961 96991 157989
rect 108099 158147 108127 158175
rect 108161 158147 108189 158175
rect 108099 158085 108127 158113
rect 108161 158085 108189 158113
rect 108099 158023 108127 158051
rect 108161 158023 108189 158051
rect 108099 157961 108127 157989
rect 108161 157961 108189 157989
rect 100419 155147 100447 155175
rect 100481 155147 100509 155175
rect 100419 155085 100447 155113
rect 100481 155085 100509 155113
rect 100419 155023 100447 155051
rect 100481 155023 100509 155051
rect 100419 154961 100447 154989
rect 100481 154961 100509 154989
rect 110277 155147 110305 155175
rect 110339 155147 110367 155175
rect 110401 155147 110429 155175
rect 110463 155147 110491 155175
rect 110277 155085 110305 155113
rect 110339 155085 110367 155113
rect 110401 155085 110429 155113
rect 110463 155085 110491 155113
rect 110277 155023 110305 155051
rect 110339 155023 110367 155051
rect 110401 155023 110429 155051
rect 110463 155023 110491 155051
rect 110277 154961 110305 154989
rect 110339 154961 110367 154989
rect 110401 154961 110429 154989
rect 110463 154961 110491 154989
rect 96777 149147 96805 149175
rect 96839 149147 96867 149175
rect 96901 149147 96929 149175
rect 96963 149147 96991 149175
rect 96777 149085 96805 149113
rect 96839 149085 96867 149113
rect 96901 149085 96929 149113
rect 96963 149085 96991 149113
rect 96777 149023 96805 149051
rect 96839 149023 96867 149051
rect 96901 149023 96929 149051
rect 96963 149023 96991 149051
rect 96777 148961 96805 148989
rect 96839 148961 96867 148989
rect 96901 148961 96929 148989
rect 96963 148961 96991 148989
rect 108099 149147 108127 149175
rect 108161 149147 108189 149175
rect 108099 149085 108127 149113
rect 108161 149085 108189 149113
rect 108099 149023 108127 149051
rect 108161 149023 108189 149051
rect 108099 148961 108127 148989
rect 108161 148961 108189 148989
rect 100419 146147 100447 146175
rect 100481 146147 100509 146175
rect 100419 146085 100447 146113
rect 100481 146085 100509 146113
rect 100419 146023 100447 146051
rect 100481 146023 100509 146051
rect 100419 145961 100447 145989
rect 100481 145961 100509 145989
rect 110277 146147 110305 146175
rect 110339 146147 110367 146175
rect 110401 146147 110429 146175
rect 110463 146147 110491 146175
rect 110277 146085 110305 146113
rect 110339 146085 110367 146113
rect 110401 146085 110429 146113
rect 110463 146085 110491 146113
rect 110277 146023 110305 146051
rect 110339 146023 110367 146051
rect 110401 146023 110429 146051
rect 110463 146023 110491 146051
rect 110277 145961 110305 145989
rect 110339 145961 110367 145989
rect 110401 145961 110429 145989
rect 110463 145961 110491 145989
rect 96777 140147 96805 140175
rect 96839 140147 96867 140175
rect 96901 140147 96929 140175
rect 96963 140147 96991 140175
rect 96777 140085 96805 140113
rect 96839 140085 96867 140113
rect 96901 140085 96929 140113
rect 96963 140085 96991 140113
rect 96777 140023 96805 140051
rect 96839 140023 96867 140051
rect 96901 140023 96929 140051
rect 96963 140023 96991 140051
rect 96777 139961 96805 139989
rect 96839 139961 96867 139989
rect 96901 139961 96929 139989
rect 96963 139961 96991 139989
rect 108099 140147 108127 140175
rect 108161 140147 108189 140175
rect 108099 140085 108127 140113
rect 108161 140085 108189 140113
rect 108099 140023 108127 140051
rect 108161 140023 108189 140051
rect 108099 139961 108127 139989
rect 108161 139961 108189 139989
rect 100419 137147 100447 137175
rect 100481 137147 100509 137175
rect 100419 137085 100447 137113
rect 100481 137085 100509 137113
rect 100419 137023 100447 137051
rect 100481 137023 100509 137051
rect 100419 136961 100447 136989
rect 100481 136961 100509 136989
rect 110277 137147 110305 137175
rect 110339 137147 110367 137175
rect 110401 137147 110429 137175
rect 110463 137147 110491 137175
rect 110277 137085 110305 137113
rect 110339 137085 110367 137113
rect 110401 137085 110429 137113
rect 110463 137085 110491 137113
rect 110277 137023 110305 137051
rect 110339 137023 110367 137051
rect 110401 137023 110429 137051
rect 110463 137023 110491 137051
rect 110277 136961 110305 136989
rect 110339 136961 110367 136989
rect 110401 136961 110429 136989
rect 110463 136961 110491 136989
rect 96777 131147 96805 131175
rect 96839 131147 96867 131175
rect 96901 131147 96929 131175
rect 96963 131147 96991 131175
rect 96777 131085 96805 131113
rect 96839 131085 96867 131113
rect 96901 131085 96929 131113
rect 96963 131085 96991 131113
rect 96777 131023 96805 131051
rect 96839 131023 96867 131051
rect 96901 131023 96929 131051
rect 96963 131023 96991 131051
rect 96777 130961 96805 130989
rect 96839 130961 96867 130989
rect 96901 130961 96929 130989
rect 96963 130961 96991 130989
rect 108099 131147 108127 131175
rect 108161 131147 108189 131175
rect 108099 131085 108127 131113
rect 108161 131085 108189 131113
rect 108099 131023 108127 131051
rect 108161 131023 108189 131051
rect 108099 130961 108127 130989
rect 108161 130961 108189 130989
rect 100419 128147 100447 128175
rect 100481 128147 100509 128175
rect 100419 128085 100447 128113
rect 100481 128085 100509 128113
rect 100419 128023 100447 128051
rect 100481 128023 100509 128051
rect 100419 127961 100447 127989
rect 100481 127961 100509 127989
rect 110277 128147 110305 128175
rect 110339 128147 110367 128175
rect 110401 128147 110429 128175
rect 110463 128147 110491 128175
rect 110277 128085 110305 128113
rect 110339 128085 110367 128113
rect 110401 128085 110429 128113
rect 110463 128085 110491 128113
rect 110277 128023 110305 128051
rect 110339 128023 110367 128051
rect 110401 128023 110429 128051
rect 110463 128023 110491 128051
rect 110277 127961 110305 127989
rect 110339 127961 110367 127989
rect 110401 127961 110429 127989
rect 110463 127961 110491 127989
rect 96777 122147 96805 122175
rect 96839 122147 96867 122175
rect 96901 122147 96929 122175
rect 96963 122147 96991 122175
rect 96777 122085 96805 122113
rect 96839 122085 96867 122113
rect 96901 122085 96929 122113
rect 96963 122085 96991 122113
rect 96777 122023 96805 122051
rect 96839 122023 96867 122051
rect 96901 122023 96929 122051
rect 96963 122023 96991 122051
rect 96777 121961 96805 121989
rect 96839 121961 96867 121989
rect 96901 121961 96929 121989
rect 96963 121961 96991 121989
rect 108099 122147 108127 122175
rect 108161 122147 108189 122175
rect 108099 122085 108127 122113
rect 108161 122085 108189 122113
rect 108099 122023 108127 122051
rect 108161 122023 108189 122051
rect 108099 121961 108127 121989
rect 108161 121961 108189 121989
rect 100419 119147 100447 119175
rect 100481 119147 100509 119175
rect 100419 119085 100447 119113
rect 100481 119085 100509 119113
rect 100419 119023 100447 119051
rect 100481 119023 100509 119051
rect 100419 118961 100447 118989
rect 100481 118961 100509 118989
rect 110277 119147 110305 119175
rect 110339 119147 110367 119175
rect 110401 119147 110429 119175
rect 110463 119147 110491 119175
rect 110277 119085 110305 119113
rect 110339 119085 110367 119113
rect 110401 119085 110429 119113
rect 110463 119085 110491 119113
rect 110277 119023 110305 119051
rect 110339 119023 110367 119051
rect 110401 119023 110429 119051
rect 110463 119023 110491 119051
rect 110277 118961 110305 118989
rect 110339 118961 110367 118989
rect 110401 118961 110429 118989
rect 110463 118961 110491 118989
rect 96777 113147 96805 113175
rect 96839 113147 96867 113175
rect 96901 113147 96929 113175
rect 96963 113147 96991 113175
rect 96777 113085 96805 113113
rect 96839 113085 96867 113113
rect 96901 113085 96929 113113
rect 96963 113085 96991 113113
rect 96777 113023 96805 113051
rect 96839 113023 96867 113051
rect 96901 113023 96929 113051
rect 96963 113023 96991 113051
rect 96777 112961 96805 112989
rect 96839 112961 96867 112989
rect 96901 112961 96929 112989
rect 96963 112961 96991 112989
rect 108099 113147 108127 113175
rect 108161 113147 108189 113175
rect 108099 113085 108127 113113
rect 108161 113085 108189 113113
rect 108099 113023 108127 113051
rect 108161 113023 108189 113051
rect 108099 112961 108127 112989
rect 108161 112961 108189 112989
rect 100419 110147 100447 110175
rect 100481 110147 100509 110175
rect 100419 110085 100447 110113
rect 100481 110085 100509 110113
rect 100419 110023 100447 110051
rect 100481 110023 100509 110051
rect 100419 109961 100447 109989
rect 100481 109961 100509 109989
rect 110277 110147 110305 110175
rect 110339 110147 110367 110175
rect 110401 110147 110429 110175
rect 110463 110147 110491 110175
rect 110277 110085 110305 110113
rect 110339 110085 110367 110113
rect 110401 110085 110429 110113
rect 110463 110085 110491 110113
rect 110277 110023 110305 110051
rect 110339 110023 110367 110051
rect 110401 110023 110429 110051
rect 110463 110023 110491 110051
rect 110277 109961 110305 109989
rect 110339 109961 110367 109989
rect 110401 109961 110429 109989
rect 110463 109961 110491 109989
rect 96777 104147 96805 104175
rect 96839 104147 96867 104175
rect 96901 104147 96929 104175
rect 96963 104147 96991 104175
rect 96777 104085 96805 104113
rect 96839 104085 96867 104113
rect 96901 104085 96929 104113
rect 96963 104085 96991 104113
rect 96777 104023 96805 104051
rect 96839 104023 96867 104051
rect 96901 104023 96929 104051
rect 96963 104023 96991 104051
rect 96777 103961 96805 103989
rect 96839 103961 96867 103989
rect 96901 103961 96929 103989
rect 96963 103961 96991 103989
rect 108099 104147 108127 104175
rect 108161 104147 108189 104175
rect 108099 104085 108127 104113
rect 108161 104085 108189 104113
rect 108099 104023 108127 104051
rect 108161 104023 108189 104051
rect 108099 103961 108127 103989
rect 108161 103961 108189 103989
rect 100419 101147 100447 101175
rect 100481 101147 100509 101175
rect 100419 101085 100447 101113
rect 100481 101085 100509 101113
rect 100419 101023 100447 101051
rect 100481 101023 100509 101051
rect 100419 100961 100447 100989
rect 100481 100961 100509 100989
rect 110277 101147 110305 101175
rect 110339 101147 110367 101175
rect 110401 101147 110429 101175
rect 110463 101147 110491 101175
rect 110277 101085 110305 101113
rect 110339 101085 110367 101113
rect 110401 101085 110429 101113
rect 110463 101085 110491 101113
rect 110277 101023 110305 101051
rect 110339 101023 110367 101051
rect 110401 101023 110429 101051
rect 110463 101023 110491 101051
rect 110277 100961 110305 100989
rect 110339 100961 110367 100989
rect 110401 100961 110429 100989
rect 110463 100961 110491 100989
rect 96777 95147 96805 95175
rect 96839 95147 96867 95175
rect 96901 95147 96929 95175
rect 96963 95147 96991 95175
rect 96777 95085 96805 95113
rect 96839 95085 96867 95113
rect 96901 95085 96929 95113
rect 96963 95085 96991 95113
rect 96777 95023 96805 95051
rect 96839 95023 96867 95051
rect 96901 95023 96929 95051
rect 96963 95023 96991 95051
rect 96777 94961 96805 94989
rect 96839 94961 96867 94989
rect 96901 94961 96929 94989
rect 96963 94961 96991 94989
rect 108099 95147 108127 95175
rect 108161 95147 108189 95175
rect 108099 95085 108127 95113
rect 108161 95085 108189 95113
rect 108099 95023 108127 95051
rect 108161 95023 108189 95051
rect 108099 94961 108127 94989
rect 108161 94961 108189 94989
rect 100419 92147 100447 92175
rect 100481 92147 100509 92175
rect 100419 92085 100447 92113
rect 100481 92085 100509 92113
rect 100419 92023 100447 92051
rect 100481 92023 100509 92051
rect 100419 91961 100447 91989
rect 100481 91961 100509 91989
rect 110277 92147 110305 92175
rect 110339 92147 110367 92175
rect 110401 92147 110429 92175
rect 110463 92147 110491 92175
rect 110277 92085 110305 92113
rect 110339 92085 110367 92113
rect 110401 92085 110429 92113
rect 110463 92085 110491 92113
rect 110277 92023 110305 92051
rect 110339 92023 110367 92051
rect 110401 92023 110429 92051
rect 110463 92023 110491 92051
rect 110277 91961 110305 91989
rect 110339 91961 110367 91989
rect 110401 91961 110429 91989
rect 110463 91961 110491 91989
rect 96777 86147 96805 86175
rect 96839 86147 96867 86175
rect 96901 86147 96929 86175
rect 96963 86147 96991 86175
rect 96777 86085 96805 86113
rect 96839 86085 96867 86113
rect 96901 86085 96929 86113
rect 96963 86085 96991 86113
rect 96777 86023 96805 86051
rect 96839 86023 96867 86051
rect 96901 86023 96929 86051
rect 96963 86023 96991 86051
rect 96777 85961 96805 85989
rect 96839 85961 96867 85989
rect 96901 85961 96929 85989
rect 96963 85961 96991 85989
rect 108099 86147 108127 86175
rect 108161 86147 108189 86175
rect 108099 86085 108127 86113
rect 108161 86085 108189 86113
rect 108099 86023 108127 86051
rect 108161 86023 108189 86051
rect 108099 85961 108127 85989
rect 108161 85961 108189 85989
rect 100419 83147 100447 83175
rect 100481 83147 100509 83175
rect 100419 83085 100447 83113
rect 100481 83085 100509 83113
rect 100419 83023 100447 83051
rect 100481 83023 100509 83051
rect 100419 82961 100447 82989
rect 100481 82961 100509 82989
rect 110277 83147 110305 83175
rect 110339 83147 110367 83175
rect 110401 83147 110429 83175
rect 110463 83147 110491 83175
rect 110277 83085 110305 83113
rect 110339 83085 110367 83113
rect 110401 83085 110429 83113
rect 110463 83085 110491 83113
rect 110277 83023 110305 83051
rect 110339 83023 110367 83051
rect 110401 83023 110429 83051
rect 110463 83023 110491 83051
rect 110277 82961 110305 82989
rect 110339 82961 110367 82989
rect 110401 82961 110429 82989
rect 110463 82961 110491 82989
rect 96777 77147 96805 77175
rect 96839 77147 96867 77175
rect 96901 77147 96929 77175
rect 96963 77147 96991 77175
rect 96777 77085 96805 77113
rect 96839 77085 96867 77113
rect 96901 77085 96929 77113
rect 96963 77085 96991 77113
rect 96777 77023 96805 77051
rect 96839 77023 96867 77051
rect 96901 77023 96929 77051
rect 96963 77023 96991 77051
rect 96777 76961 96805 76989
rect 96839 76961 96867 76989
rect 96901 76961 96929 76989
rect 96963 76961 96991 76989
rect 108099 77147 108127 77175
rect 108161 77147 108189 77175
rect 108099 77085 108127 77113
rect 108161 77085 108189 77113
rect 108099 77023 108127 77051
rect 108161 77023 108189 77051
rect 108099 76961 108127 76989
rect 108161 76961 108189 76989
rect 100419 74147 100447 74175
rect 100481 74147 100509 74175
rect 100419 74085 100447 74113
rect 100481 74085 100509 74113
rect 100419 74023 100447 74051
rect 100481 74023 100509 74051
rect 100419 73961 100447 73989
rect 100481 73961 100509 73989
rect 110277 74147 110305 74175
rect 110339 74147 110367 74175
rect 110401 74147 110429 74175
rect 110463 74147 110491 74175
rect 110277 74085 110305 74113
rect 110339 74085 110367 74113
rect 110401 74085 110429 74113
rect 110463 74085 110491 74113
rect 110277 74023 110305 74051
rect 110339 74023 110367 74051
rect 110401 74023 110429 74051
rect 110463 74023 110491 74051
rect 110277 73961 110305 73989
rect 110339 73961 110367 73989
rect 110401 73961 110429 73989
rect 110463 73961 110491 73989
rect 96777 68147 96805 68175
rect 96839 68147 96867 68175
rect 96901 68147 96929 68175
rect 96963 68147 96991 68175
rect 96777 68085 96805 68113
rect 96839 68085 96867 68113
rect 96901 68085 96929 68113
rect 96963 68085 96991 68113
rect 96777 68023 96805 68051
rect 96839 68023 96867 68051
rect 96901 68023 96929 68051
rect 96963 68023 96991 68051
rect 96777 67961 96805 67989
rect 96839 67961 96867 67989
rect 96901 67961 96929 67989
rect 96963 67961 96991 67989
rect 108099 68147 108127 68175
rect 108161 68147 108189 68175
rect 108099 68085 108127 68113
rect 108161 68085 108189 68113
rect 108099 68023 108127 68051
rect 108161 68023 108189 68051
rect 108099 67961 108127 67989
rect 108161 67961 108189 67989
rect 100419 65147 100447 65175
rect 100481 65147 100509 65175
rect 100419 65085 100447 65113
rect 100481 65085 100509 65113
rect 100419 65023 100447 65051
rect 100481 65023 100509 65051
rect 100419 64961 100447 64989
rect 100481 64961 100509 64989
rect 110277 65147 110305 65175
rect 110339 65147 110367 65175
rect 110401 65147 110429 65175
rect 110463 65147 110491 65175
rect 110277 65085 110305 65113
rect 110339 65085 110367 65113
rect 110401 65085 110429 65113
rect 110463 65085 110491 65113
rect 110277 65023 110305 65051
rect 110339 65023 110367 65051
rect 110401 65023 110429 65051
rect 110463 65023 110491 65051
rect 110277 64961 110305 64989
rect 110339 64961 110367 64989
rect 110401 64961 110429 64989
rect 110463 64961 110491 64989
rect 96777 59147 96805 59175
rect 96839 59147 96867 59175
rect 96901 59147 96929 59175
rect 96963 59147 96991 59175
rect 96777 59085 96805 59113
rect 96839 59085 96867 59113
rect 96901 59085 96929 59113
rect 96963 59085 96991 59113
rect 96777 59023 96805 59051
rect 96839 59023 96867 59051
rect 96901 59023 96929 59051
rect 96963 59023 96991 59051
rect 96777 58961 96805 58989
rect 96839 58961 96867 58989
rect 96901 58961 96929 58989
rect 96963 58961 96991 58989
rect 108099 59147 108127 59175
rect 108161 59147 108189 59175
rect 108099 59085 108127 59113
rect 108161 59085 108189 59113
rect 108099 59023 108127 59051
rect 108161 59023 108189 59051
rect 108099 58961 108127 58989
rect 108161 58961 108189 58989
rect 100419 56147 100447 56175
rect 100481 56147 100509 56175
rect 100419 56085 100447 56113
rect 100481 56085 100509 56113
rect 100419 56023 100447 56051
rect 100481 56023 100509 56051
rect 100419 55961 100447 55989
rect 100481 55961 100509 55989
rect 110277 56147 110305 56175
rect 110339 56147 110367 56175
rect 110401 56147 110429 56175
rect 110463 56147 110491 56175
rect 110277 56085 110305 56113
rect 110339 56085 110367 56113
rect 110401 56085 110429 56113
rect 110463 56085 110491 56113
rect 110277 56023 110305 56051
rect 110339 56023 110367 56051
rect 110401 56023 110429 56051
rect 110463 56023 110491 56051
rect 110277 55961 110305 55989
rect 110339 55961 110367 55989
rect 110401 55961 110429 55989
rect 110463 55961 110491 55989
rect 96777 50147 96805 50175
rect 96839 50147 96867 50175
rect 96901 50147 96929 50175
rect 96963 50147 96991 50175
rect 96777 50085 96805 50113
rect 96839 50085 96867 50113
rect 96901 50085 96929 50113
rect 96963 50085 96991 50113
rect 96777 50023 96805 50051
rect 96839 50023 96867 50051
rect 96901 50023 96929 50051
rect 96963 50023 96991 50051
rect 96777 49961 96805 49989
rect 96839 49961 96867 49989
rect 96901 49961 96929 49989
rect 96963 49961 96991 49989
rect 108099 50147 108127 50175
rect 108161 50147 108189 50175
rect 108099 50085 108127 50113
rect 108161 50085 108189 50113
rect 108099 50023 108127 50051
rect 108161 50023 108189 50051
rect 108099 49961 108127 49989
rect 108161 49961 108189 49989
rect 100419 47147 100447 47175
rect 100481 47147 100509 47175
rect 100419 47085 100447 47113
rect 100481 47085 100509 47113
rect 100419 47023 100447 47051
rect 100481 47023 100509 47051
rect 100419 46961 100447 46989
rect 100481 46961 100509 46989
rect 110277 47147 110305 47175
rect 110339 47147 110367 47175
rect 110401 47147 110429 47175
rect 110463 47147 110491 47175
rect 110277 47085 110305 47113
rect 110339 47085 110367 47113
rect 110401 47085 110429 47113
rect 110463 47085 110491 47113
rect 110277 47023 110305 47051
rect 110339 47023 110367 47051
rect 110401 47023 110429 47051
rect 110463 47023 110491 47051
rect 110277 46961 110305 46989
rect 110339 46961 110367 46989
rect 110401 46961 110429 46989
rect 110463 46961 110491 46989
rect 96777 41147 96805 41175
rect 96839 41147 96867 41175
rect 96901 41147 96929 41175
rect 96963 41147 96991 41175
rect 96777 41085 96805 41113
rect 96839 41085 96867 41113
rect 96901 41085 96929 41113
rect 96963 41085 96991 41113
rect 96777 41023 96805 41051
rect 96839 41023 96867 41051
rect 96901 41023 96929 41051
rect 96963 41023 96991 41051
rect 96777 40961 96805 40989
rect 96839 40961 96867 40989
rect 96901 40961 96929 40989
rect 96963 40961 96991 40989
rect 108099 41147 108127 41175
rect 108161 41147 108189 41175
rect 108099 41085 108127 41113
rect 108161 41085 108189 41113
rect 108099 41023 108127 41051
rect 108161 41023 108189 41051
rect 108099 40961 108127 40989
rect 108161 40961 108189 40989
rect 100419 38147 100447 38175
rect 100481 38147 100509 38175
rect 100419 38085 100447 38113
rect 100481 38085 100509 38113
rect 100419 38023 100447 38051
rect 100481 38023 100509 38051
rect 100419 37961 100447 37989
rect 100481 37961 100509 37989
rect 110277 38147 110305 38175
rect 110339 38147 110367 38175
rect 110401 38147 110429 38175
rect 110463 38147 110491 38175
rect 110277 38085 110305 38113
rect 110339 38085 110367 38113
rect 110401 38085 110429 38113
rect 110463 38085 110491 38113
rect 110277 38023 110305 38051
rect 110339 38023 110367 38051
rect 110401 38023 110429 38051
rect 110463 38023 110491 38051
rect 110277 37961 110305 37989
rect 110339 37961 110367 37989
rect 110401 37961 110429 37989
rect 110463 37961 110491 37989
rect 96777 32147 96805 32175
rect 96839 32147 96867 32175
rect 96901 32147 96929 32175
rect 96963 32147 96991 32175
rect 96777 32085 96805 32113
rect 96839 32085 96867 32113
rect 96901 32085 96929 32113
rect 96963 32085 96991 32113
rect 96777 32023 96805 32051
rect 96839 32023 96867 32051
rect 96901 32023 96929 32051
rect 96963 32023 96991 32051
rect 96777 31961 96805 31989
rect 96839 31961 96867 31989
rect 96901 31961 96929 31989
rect 96963 31961 96991 31989
rect 108099 32147 108127 32175
rect 108161 32147 108189 32175
rect 108099 32085 108127 32113
rect 108161 32085 108189 32113
rect 108099 32023 108127 32051
rect 108161 32023 108189 32051
rect 108099 31961 108127 31989
rect 108161 31961 108189 31989
rect 100419 29147 100447 29175
rect 100481 29147 100509 29175
rect 100419 29085 100447 29113
rect 100481 29085 100509 29113
rect 100419 29023 100447 29051
rect 100481 29023 100509 29051
rect 100419 28961 100447 28989
rect 100481 28961 100509 28989
rect 110277 29147 110305 29175
rect 110339 29147 110367 29175
rect 110401 29147 110429 29175
rect 110463 29147 110491 29175
rect 110277 29085 110305 29113
rect 110339 29085 110367 29113
rect 110401 29085 110429 29113
rect 110463 29085 110491 29113
rect 110277 29023 110305 29051
rect 110339 29023 110367 29051
rect 110401 29023 110429 29051
rect 110463 29023 110491 29051
rect 110277 28961 110305 28989
rect 110339 28961 110367 28989
rect 110401 28961 110429 28989
rect 110463 28961 110491 28989
rect 96777 23147 96805 23175
rect 96839 23147 96867 23175
rect 96901 23147 96929 23175
rect 96963 23147 96991 23175
rect 96777 23085 96805 23113
rect 96839 23085 96867 23113
rect 96901 23085 96929 23113
rect 96963 23085 96991 23113
rect 96777 23023 96805 23051
rect 96839 23023 96867 23051
rect 96901 23023 96929 23051
rect 96963 23023 96991 23051
rect 96777 22961 96805 22989
rect 96839 22961 96867 22989
rect 96901 22961 96929 22989
rect 96963 22961 96991 22989
rect 108099 23147 108127 23175
rect 108161 23147 108189 23175
rect 108099 23085 108127 23113
rect 108161 23085 108189 23113
rect 108099 23023 108127 23051
rect 108161 23023 108189 23051
rect 108099 22961 108127 22989
rect 108161 22961 108189 22989
rect 100419 20147 100447 20175
rect 100481 20147 100509 20175
rect 100419 20085 100447 20113
rect 100481 20085 100509 20113
rect 100419 20023 100447 20051
rect 100481 20023 100509 20051
rect 100419 19961 100447 19989
rect 100481 19961 100509 19989
rect 110277 20147 110305 20175
rect 110339 20147 110367 20175
rect 110401 20147 110429 20175
rect 110463 20147 110491 20175
rect 110277 20085 110305 20113
rect 110339 20085 110367 20113
rect 110401 20085 110429 20113
rect 110463 20085 110491 20113
rect 110277 20023 110305 20051
rect 110339 20023 110367 20051
rect 110401 20023 110429 20051
rect 110463 20023 110491 20051
rect 110277 19961 110305 19989
rect 110339 19961 110367 19989
rect 110401 19961 110429 19989
rect 110463 19961 110491 19989
rect 96777 14147 96805 14175
rect 96839 14147 96867 14175
rect 96901 14147 96929 14175
rect 96963 14147 96991 14175
rect 96777 14085 96805 14113
rect 96839 14085 96867 14113
rect 96901 14085 96929 14113
rect 96963 14085 96991 14113
rect 96777 14023 96805 14051
rect 96839 14023 96867 14051
rect 96901 14023 96929 14051
rect 96963 14023 96991 14051
rect 96777 13961 96805 13989
rect 96839 13961 96867 13989
rect 96901 13961 96929 13989
rect 96963 13961 96991 13989
rect 108099 14147 108127 14175
rect 108161 14147 108189 14175
rect 108099 14085 108127 14113
rect 108161 14085 108189 14113
rect 108099 14023 108127 14051
rect 108161 14023 108189 14051
rect 108099 13961 108127 13989
rect 108161 13961 108189 13989
rect 100419 11147 100447 11175
rect 100481 11147 100509 11175
rect 100419 11085 100447 11113
rect 100481 11085 100509 11113
rect 100419 11023 100447 11051
rect 100481 11023 100509 11051
rect 100419 10961 100447 10989
rect 100481 10961 100509 10989
rect 110277 11147 110305 11175
rect 110339 11147 110367 11175
rect 110401 11147 110429 11175
rect 110463 11147 110491 11175
rect 110277 11085 110305 11113
rect 110339 11085 110367 11113
rect 110401 11085 110429 11113
rect 110463 11085 110491 11113
rect 110277 11023 110305 11051
rect 110339 11023 110367 11051
rect 110401 11023 110429 11051
rect 110463 11023 110491 11051
rect 110277 10961 110305 10989
rect 110339 10961 110367 10989
rect 110401 10961 110429 10989
rect 110463 10961 110491 10989
rect 96777 5147 96805 5175
rect 96839 5147 96867 5175
rect 96901 5147 96929 5175
rect 96963 5147 96991 5175
rect 96777 5085 96805 5113
rect 96839 5085 96867 5113
rect 96901 5085 96929 5113
rect 96963 5085 96991 5113
rect 96777 5023 96805 5051
rect 96839 5023 96867 5051
rect 96901 5023 96929 5051
rect 96963 5023 96991 5051
rect 96777 4961 96805 4989
rect 96839 4961 96867 4989
rect 96901 4961 96929 4989
rect 96963 4961 96991 4989
rect 108099 5147 108127 5175
rect 108161 5147 108189 5175
rect 108099 5085 108127 5113
rect 108161 5085 108189 5113
rect 108099 5023 108127 5051
rect 108161 5023 108189 5051
rect 108099 4961 108127 4989
rect 108161 4961 108189 4989
rect 96777 -588 96805 -560
rect 96839 -588 96867 -560
rect 96901 -588 96929 -560
rect 96963 -588 96991 -560
rect 96777 -650 96805 -622
rect 96839 -650 96867 -622
rect 96901 -650 96929 -622
rect 96963 -650 96991 -622
rect 96777 -712 96805 -684
rect 96839 -712 96867 -684
rect 96901 -712 96929 -684
rect 96963 -712 96991 -684
rect 96777 -774 96805 -746
rect 96839 -774 96867 -746
rect 96901 -774 96929 -746
rect 96963 -774 96991 -746
rect 110277 2147 110305 2175
rect 110339 2147 110367 2175
rect 110401 2147 110429 2175
rect 110463 2147 110491 2175
rect 110277 2085 110305 2113
rect 110339 2085 110367 2113
rect 110401 2085 110429 2113
rect 110463 2085 110491 2113
rect 110277 2023 110305 2051
rect 110339 2023 110367 2051
rect 110401 2023 110429 2051
rect 110463 2023 110491 2051
rect 110277 1961 110305 1989
rect 110339 1961 110367 1989
rect 110401 1961 110429 1989
rect 110463 1961 110491 1989
rect 110277 -108 110305 -80
rect 110339 -108 110367 -80
rect 110401 -108 110429 -80
rect 110463 -108 110491 -80
rect 110277 -170 110305 -142
rect 110339 -170 110367 -142
rect 110401 -170 110429 -142
rect 110463 -170 110491 -142
rect 110277 -232 110305 -204
rect 110339 -232 110367 -204
rect 110401 -232 110429 -204
rect 110463 -232 110491 -204
rect 110277 -294 110305 -266
rect 110339 -294 110367 -266
rect 110401 -294 110429 -266
rect 110463 -294 110491 -266
rect 112137 299058 112165 299086
rect 112199 299058 112227 299086
rect 112261 299058 112289 299086
rect 112323 299058 112351 299086
rect 112137 298996 112165 299024
rect 112199 298996 112227 299024
rect 112261 298996 112289 299024
rect 112323 298996 112351 299024
rect 112137 298934 112165 298962
rect 112199 298934 112227 298962
rect 112261 298934 112289 298962
rect 112323 298934 112351 298962
rect 112137 298872 112165 298900
rect 112199 298872 112227 298900
rect 112261 298872 112289 298900
rect 112323 298872 112351 298900
rect 112137 293147 112165 293175
rect 112199 293147 112227 293175
rect 112261 293147 112289 293175
rect 112323 293147 112351 293175
rect 112137 293085 112165 293113
rect 112199 293085 112227 293113
rect 112261 293085 112289 293113
rect 112323 293085 112351 293113
rect 112137 293023 112165 293051
rect 112199 293023 112227 293051
rect 112261 293023 112289 293051
rect 112323 293023 112351 293051
rect 112137 292961 112165 292989
rect 112199 292961 112227 292989
rect 112261 292961 112289 292989
rect 112323 292961 112351 292989
rect 112137 284147 112165 284175
rect 112199 284147 112227 284175
rect 112261 284147 112289 284175
rect 112323 284147 112351 284175
rect 112137 284085 112165 284113
rect 112199 284085 112227 284113
rect 112261 284085 112289 284113
rect 112323 284085 112351 284113
rect 112137 284023 112165 284051
rect 112199 284023 112227 284051
rect 112261 284023 112289 284051
rect 112323 284023 112351 284051
rect 112137 283961 112165 283989
rect 112199 283961 112227 283989
rect 112261 283961 112289 283989
rect 112323 283961 112351 283989
rect 112137 275147 112165 275175
rect 112199 275147 112227 275175
rect 112261 275147 112289 275175
rect 112323 275147 112351 275175
rect 112137 275085 112165 275113
rect 112199 275085 112227 275113
rect 112261 275085 112289 275113
rect 112323 275085 112351 275113
rect 112137 275023 112165 275051
rect 112199 275023 112227 275051
rect 112261 275023 112289 275051
rect 112323 275023 112351 275051
rect 112137 274961 112165 274989
rect 112199 274961 112227 274989
rect 112261 274961 112289 274989
rect 112323 274961 112351 274989
rect 112137 266147 112165 266175
rect 112199 266147 112227 266175
rect 112261 266147 112289 266175
rect 112323 266147 112351 266175
rect 112137 266085 112165 266113
rect 112199 266085 112227 266113
rect 112261 266085 112289 266113
rect 112323 266085 112351 266113
rect 112137 266023 112165 266051
rect 112199 266023 112227 266051
rect 112261 266023 112289 266051
rect 112323 266023 112351 266051
rect 112137 265961 112165 265989
rect 112199 265961 112227 265989
rect 112261 265961 112289 265989
rect 112323 265961 112351 265989
rect 112137 257147 112165 257175
rect 112199 257147 112227 257175
rect 112261 257147 112289 257175
rect 112323 257147 112351 257175
rect 112137 257085 112165 257113
rect 112199 257085 112227 257113
rect 112261 257085 112289 257113
rect 112323 257085 112351 257113
rect 112137 257023 112165 257051
rect 112199 257023 112227 257051
rect 112261 257023 112289 257051
rect 112323 257023 112351 257051
rect 112137 256961 112165 256989
rect 112199 256961 112227 256989
rect 112261 256961 112289 256989
rect 112323 256961 112351 256989
rect 112137 248147 112165 248175
rect 112199 248147 112227 248175
rect 112261 248147 112289 248175
rect 112323 248147 112351 248175
rect 112137 248085 112165 248113
rect 112199 248085 112227 248113
rect 112261 248085 112289 248113
rect 112323 248085 112351 248113
rect 112137 248023 112165 248051
rect 112199 248023 112227 248051
rect 112261 248023 112289 248051
rect 112323 248023 112351 248051
rect 112137 247961 112165 247989
rect 112199 247961 112227 247989
rect 112261 247961 112289 247989
rect 112323 247961 112351 247989
rect 112137 239147 112165 239175
rect 112199 239147 112227 239175
rect 112261 239147 112289 239175
rect 112323 239147 112351 239175
rect 112137 239085 112165 239113
rect 112199 239085 112227 239113
rect 112261 239085 112289 239113
rect 112323 239085 112351 239113
rect 112137 239023 112165 239051
rect 112199 239023 112227 239051
rect 112261 239023 112289 239051
rect 112323 239023 112351 239051
rect 112137 238961 112165 238989
rect 112199 238961 112227 238989
rect 112261 238961 112289 238989
rect 112323 238961 112351 238989
rect 112137 230147 112165 230175
rect 112199 230147 112227 230175
rect 112261 230147 112289 230175
rect 112323 230147 112351 230175
rect 112137 230085 112165 230113
rect 112199 230085 112227 230113
rect 112261 230085 112289 230113
rect 112323 230085 112351 230113
rect 112137 230023 112165 230051
rect 112199 230023 112227 230051
rect 112261 230023 112289 230051
rect 112323 230023 112351 230051
rect 112137 229961 112165 229989
rect 112199 229961 112227 229989
rect 112261 229961 112289 229989
rect 112323 229961 112351 229989
rect 112137 221147 112165 221175
rect 112199 221147 112227 221175
rect 112261 221147 112289 221175
rect 112323 221147 112351 221175
rect 112137 221085 112165 221113
rect 112199 221085 112227 221113
rect 112261 221085 112289 221113
rect 112323 221085 112351 221113
rect 112137 221023 112165 221051
rect 112199 221023 112227 221051
rect 112261 221023 112289 221051
rect 112323 221023 112351 221051
rect 112137 220961 112165 220989
rect 112199 220961 112227 220989
rect 112261 220961 112289 220989
rect 112323 220961 112351 220989
rect 112137 212147 112165 212175
rect 112199 212147 112227 212175
rect 112261 212147 112289 212175
rect 112323 212147 112351 212175
rect 112137 212085 112165 212113
rect 112199 212085 112227 212113
rect 112261 212085 112289 212113
rect 112323 212085 112351 212113
rect 112137 212023 112165 212051
rect 112199 212023 112227 212051
rect 112261 212023 112289 212051
rect 112323 212023 112351 212051
rect 112137 211961 112165 211989
rect 112199 211961 112227 211989
rect 112261 211961 112289 211989
rect 112323 211961 112351 211989
rect 112137 203147 112165 203175
rect 112199 203147 112227 203175
rect 112261 203147 112289 203175
rect 112323 203147 112351 203175
rect 112137 203085 112165 203113
rect 112199 203085 112227 203113
rect 112261 203085 112289 203113
rect 112323 203085 112351 203113
rect 112137 203023 112165 203051
rect 112199 203023 112227 203051
rect 112261 203023 112289 203051
rect 112323 203023 112351 203051
rect 112137 202961 112165 202989
rect 112199 202961 112227 202989
rect 112261 202961 112289 202989
rect 112323 202961 112351 202989
rect 112137 194147 112165 194175
rect 112199 194147 112227 194175
rect 112261 194147 112289 194175
rect 112323 194147 112351 194175
rect 112137 194085 112165 194113
rect 112199 194085 112227 194113
rect 112261 194085 112289 194113
rect 112323 194085 112351 194113
rect 112137 194023 112165 194051
rect 112199 194023 112227 194051
rect 112261 194023 112289 194051
rect 112323 194023 112351 194051
rect 112137 193961 112165 193989
rect 112199 193961 112227 193989
rect 112261 193961 112289 193989
rect 112323 193961 112351 193989
rect 112137 185147 112165 185175
rect 112199 185147 112227 185175
rect 112261 185147 112289 185175
rect 112323 185147 112351 185175
rect 112137 185085 112165 185113
rect 112199 185085 112227 185113
rect 112261 185085 112289 185113
rect 112323 185085 112351 185113
rect 112137 185023 112165 185051
rect 112199 185023 112227 185051
rect 112261 185023 112289 185051
rect 112323 185023 112351 185051
rect 112137 184961 112165 184989
rect 112199 184961 112227 184989
rect 112261 184961 112289 184989
rect 112323 184961 112351 184989
rect 112137 176147 112165 176175
rect 112199 176147 112227 176175
rect 112261 176147 112289 176175
rect 112323 176147 112351 176175
rect 112137 176085 112165 176113
rect 112199 176085 112227 176113
rect 112261 176085 112289 176113
rect 112323 176085 112351 176113
rect 112137 176023 112165 176051
rect 112199 176023 112227 176051
rect 112261 176023 112289 176051
rect 112323 176023 112351 176051
rect 112137 175961 112165 175989
rect 112199 175961 112227 175989
rect 112261 175961 112289 175989
rect 112323 175961 112351 175989
rect 125637 298578 125665 298606
rect 125699 298578 125727 298606
rect 125761 298578 125789 298606
rect 125823 298578 125851 298606
rect 125637 298516 125665 298544
rect 125699 298516 125727 298544
rect 125761 298516 125789 298544
rect 125823 298516 125851 298544
rect 125637 298454 125665 298482
rect 125699 298454 125727 298482
rect 125761 298454 125789 298482
rect 125823 298454 125851 298482
rect 125637 298392 125665 298420
rect 125699 298392 125727 298420
rect 125761 298392 125789 298420
rect 125823 298392 125851 298420
rect 125637 290147 125665 290175
rect 125699 290147 125727 290175
rect 125761 290147 125789 290175
rect 125823 290147 125851 290175
rect 125637 290085 125665 290113
rect 125699 290085 125727 290113
rect 125761 290085 125789 290113
rect 125823 290085 125851 290113
rect 125637 290023 125665 290051
rect 125699 290023 125727 290051
rect 125761 290023 125789 290051
rect 125823 290023 125851 290051
rect 125637 289961 125665 289989
rect 125699 289961 125727 289989
rect 125761 289961 125789 289989
rect 125823 289961 125851 289989
rect 125637 281147 125665 281175
rect 125699 281147 125727 281175
rect 125761 281147 125789 281175
rect 125823 281147 125851 281175
rect 125637 281085 125665 281113
rect 125699 281085 125727 281113
rect 125761 281085 125789 281113
rect 125823 281085 125851 281113
rect 125637 281023 125665 281051
rect 125699 281023 125727 281051
rect 125761 281023 125789 281051
rect 125823 281023 125851 281051
rect 125637 280961 125665 280989
rect 125699 280961 125727 280989
rect 125761 280961 125789 280989
rect 125823 280961 125851 280989
rect 125637 272147 125665 272175
rect 125699 272147 125727 272175
rect 125761 272147 125789 272175
rect 125823 272147 125851 272175
rect 125637 272085 125665 272113
rect 125699 272085 125727 272113
rect 125761 272085 125789 272113
rect 125823 272085 125851 272113
rect 125637 272023 125665 272051
rect 125699 272023 125727 272051
rect 125761 272023 125789 272051
rect 125823 272023 125851 272051
rect 125637 271961 125665 271989
rect 125699 271961 125727 271989
rect 125761 271961 125789 271989
rect 125823 271961 125851 271989
rect 125637 263147 125665 263175
rect 125699 263147 125727 263175
rect 125761 263147 125789 263175
rect 125823 263147 125851 263175
rect 125637 263085 125665 263113
rect 125699 263085 125727 263113
rect 125761 263085 125789 263113
rect 125823 263085 125851 263113
rect 125637 263023 125665 263051
rect 125699 263023 125727 263051
rect 125761 263023 125789 263051
rect 125823 263023 125851 263051
rect 125637 262961 125665 262989
rect 125699 262961 125727 262989
rect 125761 262961 125789 262989
rect 125823 262961 125851 262989
rect 125637 254147 125665 254175
rect 125699 254147 125727 254175
rect 125761 254147 125789 254175
rect 125823 254147 125851 254175
rect 125637 254085 125665 254113
rect 125699 254085 125727 254113
rect 125761 254085 125789 254113
rect 125823 254085 125851 254113
rect 125637 254023 125665 254051
rect 125699 254023 125727 254051
rect 125761 254023 125789 254051
rect 125823 254023 125851 254051
rect 125637 253961 125665 253989
rect 125699 253961 125727 253989
rect 125761 253961 125789 253989
rect 125823 253961 125851 253989
rect 125637 245147 125665 245175
rect 125699 245147 125727 245175
rect 125761 245147 125789 245175
rect 125823 245147 125851 245175
rect 125637 245085 125665 245113
rect 125699 245085 125727 245113
rect 125761 245085 125789 245113
rect 125823 245085 125851 245113
rect 125637 245023 125665 245051
rect 125699 245023 125727 245051
rect 125761 245023 125789 245051
rect 125823 245023 125851 245051
rect 125637 244961 125665 244989
rect 125699 244961 125727 244989
rect 125761 244961 125789 244989
rect 125823 244961 125851 244989
rect 125637 236147 125665 236175
rect 125699 236147 125727 236175
rect 125761 236147 125789 236175
rect 125823 236147 125851 236175
rect 125637 236085 125665 236113
rect 125699 236085 125727 236113
rect 125761 236085 125789 236113
rect 125823 236085 125851 236113
rect 125637 236023 125665 236051
rect 125699 236023 125727 236051
rect 125761 236023 125789 236051
rect 125823 236023 125851 236051
rect 125637 235961 125665 235989
rect 125699 235961 125727 235989
rect 125761 235961 125789 235989
rect 125823 235961 125851 235989
rect 125637 227147 125665 227175
rect 125699 227147 125727 227175
rect 125761 227147 125789 227175
rect 125823 227147 125851 227175
rect 125637 227085 125665 227113
rect 125699 227085 125727 227113
rect 125761 227085 125789 227113
rect 125823 227085 125851 227113
rect 125637 227023 125665 227051
rect 125699 227023 125727 227051
rect 125761 227023 125789 227051
rect 125823 227023 125851 227051
rect 125637 226961 125665 226989
rect 125699 226961 125727 226989
rect 125761 226961 125789 226989
rect 125823 226961 125851 226989
rect 125637 218147 125665 218175
rect 125699 218147 125727 218175
rect 125761 218147 125789 218175
rect 125823 218147 125851 218175
rect 125637 218085 125665 218113
rect 125699 218085 125727 218113
rect 125761 218085 125789 218113
rect 125823 218085 125851 218113
rect 125637 218023 125665 218051
rect 125699 218023 125727 218051
rect 125761 218023 125789 218051
rect 125823 218023 125851 218051
rect 125637 217961 125665 217989
rect 125699 217961 125727 217989
rect 125761 217961 125789 217989
rect 125823 217961 125851 217989
rect 125637 209147 125665 209175
rect 125699 209147 125727 209175
rect 125761 209147 125789 209175
rect 125823 209147 125851 209175
rect 125637 209085 125665 209113
rect 125699 209085 125727 209113
rect 125761 209085 125789 209113
rect 125823 209085 125851 209113
rect 125637 209023 125665 209051
rect 125699 209023 125727 209051
rect 125761 209023 125789 209051
rect 125823 209023 125851 209051
rect 125637 208961 125665 208989
rect 125699 208961 125727 208989
rect 125761 208961 125789 208989
rect 125823 208961 125851 208989
rect 125637 200147 125665 200175
rect 125699 200147 125727 200175
rect 125761 200147 125789 200175
rect 125823 200147 125851 200175
rect 125637 200085 125665 200113
rect 125699 200085 125727 200113
rect 125761 200085 125789 200113
rect 125823 200085 125851 200113
rect 125637 200023 125665 200051
rect 125699 200023 125727 200051
rect 125761 200023 125789 200051
rect 125823 200023 125851 200051
rect 125637 199961 125665 199989
rect 125699 199961 125727 199989
rect 125761 199961 125789 199989
rect 125823 199961 125851 199989
rect 125637 191147 125665 191175
rect 125699 191147 125727 191175
rect 125761 191147 125789 191175
rect 125823 191147 125851 191175
rect 125637 191085 125665 191113
rect 125699 191085 125727 191113
rect 125761 191085 125789 191113
rect 125823 191085 125851 191113
rect 125637 191023 125665 191051
rect 125699 191023 125727 191051
rect 125761 191023 125789 191051
rect 125823 191023 125851 191051
rect 125637 190961 125665 190989
rect 125699 190961 125727 190989
rect 125761 190961 125789 190989
rect 125823 190961 125851 190989
rect 125637 182147 125665 182175
rect 125699 182147 125727 182175
rect 125761 182147 125789 182175
rect 125823 182147 125851 182175
rect 125637 182085 125665 182113
rect 125699 182085 125727 182113
rect 125761 182085 125789 182113
rect 125823 182085 125851 182113
rect 125637 182023 125665 182051
rect 125699 182023 125727 182051
rect 125761 182023 125789 182051
rect 125823 182023 125851 182051
rect 125637 181961 125665 181989
rect 125699 181961 125727 181989
rect 125761 181961 125789 181989
rect 125823 181961 125851 181989
rect 115779 173147 115807 173175
rect 115841 173147 115869 173175
rect 115779 173085 115807 173113
rect 115841 173085 115869 173113
rect 115779 173023 115807 173051
rect 115841 173023 115869 173051
rect 115779 172961 115807 172989
rect 115841 172961 115869 172989
rect 125637 173147 125665 173175
rect 125699 173147 125727 173175
rect 125761 173147 125789 173175
rect 125823 173147 125851 173175
rect 125637 173085 125665 173113
rect 125699 173085 125727 173113
rect 125761 173085 125789 173113
rect 125823 173085 125851 173113
rect 125637 173023 125665 173051
rect 125699 173023 125727 173051
rect 125761 173023 125789 173051
rect 125823 173023 125851 173051
rect 125637 172961 125665 172989
rect 125699 172961 125727 172989
rect 125761 172961 125789 172989
rect 125823 172961 125851 172989
rect 112137 167147 112165 167175
rect 112199 167147 112227 167175
rect 112261 167147 112289 167175
rect 112323 167147 112351 167175
rect 112137 167085 112165 167113
rect 112199 167085 112227 167113
rect 112261 167085 112289 167113
rect 112323 167085 112351 167113
rect 112137 167023 112165 167051
rect 112199 167023 112227 167051
rect 112261 167023 112289 167051
rect 112323 167023 112351 167051
rect 112137 166961 112165 166989
rect 112199 166961 112227 166989
rect 112261 166961 112289 166989
rect 112323 166961 112351 166989
rect 123459 167147 123487 167175
rect 123521 167147 123549 167175
rect 123459 167085 123487 167113
rect 123521 167085 123549 167113
rect 123459 167023 123487 167051
rect 123521 167023 123549 167051
rect 123459 166961 123487 166989
rect 123521 166961 123549 166989
rect 115779 164147 115807 164175
rect 115841 164147 115869 164175
rect 115779 164085 115807 164113
rect 115841 164085 115869 164113
rect 115779 164023 115807 164051
rect 115841 164023 115869 164051
rect 115779 163961 115807 163989
rect 115841 163961 115869 163989
rect 125637 164147 125665 164175
rect 125699 164147 125727 164175
rect 125761 164147 125789 164175
rect 125823 164147 125851 164175
rect 125637 164085 125665 164113
rect 125699 164085 125727 164113
rect 125761 164085 125789 164113
rect 125823 164085 125851 164113
rect 125637 164023 125665 164051
rect 125699 164023 125727 164051
rect 125761 164023 125789 164051
rect 125823 164023 125851 164051
rect 125637 163961 125665 163989
rect 125699 163961 125727 163989
rect 125761 163961 125789 163989
rect 125823 163961 125851 163989
rect 112137 158147 112165 158175
rect 112199 158147 112227 158175
rect 112261 158147 112289 158175
rect 112323 158147 112351 158175
rect 112137 158085 112165 158113
rect 112199 158085 112227 158113
rect 112261 158085 112289 158113
rect 112323 158085 112351 158113
rect 112137 158023 112165 158051
rect 112199 158023 112227 158051
rect 112261 158023 112289 158051
rect 112323 158023 112351 158051
rect 112137 157961 112165 157989
rect 112199 157961 112227 157989
rect 112261 157961 112289 157989
rect 112323 157961 112351 157989
rect 123459 158147 123487 158175
rect 123521 158147 123549 158175
rect 123459 158085 123487 158113
rect 123521 158085 123549 158113
rect 123459 158023 123487 158051
rect 123521 158023 123549 158051
rect 123459 157961 123487 157989
rect 123521 157961 123549 157989
rect 115779 155147 115807 155175
rect 115841 155147 115869 155175
rect 115779 155085 115807 155113
rect 115841 155085 115869 155113
rect 115779 155023 115807 155051
rect 115841 155023 115869 155051
rect 115779 154961 115807 154989
rect 115841 154961 115869 154989
rect 125637 155147 125665 155175
rect 125699 155147 125727 155175
rect 125761 155147 125789 155175
rect 125823 155147 125851 155175
rect 125637 155085 125665 155113
rect 125699 155085 125727 155113
rect 125761 155085 125789 155113
rect 125823 155085 125851 155113
rect 125637 155023 125665 155051
rect 125699 155023 125727 155051
rect 125761 155023 125789 155051
rect 125823 155023 125851 155051
rect 125637 154961 125665 154989
rect 125699 154961 125727 154989
rect 125761 154961 125789 154989
rect 125823 154961 125851 154989
rect 112137 149147 112165 149175
rect 112199 149147 112227 149175
rect 112261 149147 112289 149175
rect 112323 149147 112351 149175
rect 112137 149085 112165 149113
rect 112199 149085 112227 149113
rect 112261 149085 112289 149113
rect 112323 149085 112351 149113
rect 112137 149023 112165 149051
rect 112199 149023 112227 149051
rect 112261 149023 112289 149051
rect 112323 149023 112351 149051
rect 112137 148961 112165 148989
rect 112199 148961 112227 148989
rect 112261 148961 112289 148989
rect 112323 148961 112351 148989
rect 123459 149147 123487 149175
rect 123521 149147 123549 149175
rect 123459 149085 123487 149113
rect 123521 149085 123549 149113
rect 123459 149023 123487 149051
rect 123521 149023 123549 149051
rect 123459 148961 123487 148989
rect 123521 148961 123549 148989
rect 115779 146147 115807 146175
rect 115841 146147 115869 146175
rect 115779 146085 115807 146113
rect 115841 146085 115869 146113
rect 115779 146023 115807 146051
rect 115841 146023 115869 146051
rect 115779 145961 115807 145989
rect 115841 145961 115869 145989
rect 125637 146147 125665 146175
rect 125699 146147 125727 146175
rect 125761 146147 125789 146175
rect 125823 146147 125851 146175
rect 125637 146085 125665 146113
rect 125699 146085 125727 146113
rect 125761 146085 125789 146113
rect 125823 146085 125851 146113
rect 125637 146023 125665 146051
rect 125699 146023 125727 146051
rect 125761 146023 125789 146051
rect 125823 146023 125851 146051
rect 125637 145961 125665 145989
rect 125699 145961 125727 145989
rect 125761 145961 125789 145989
rect 125823 145961 125851 145989
rect 112137 140147 112165 140175
rect 112199 140147 112227 140175
rect 112261 140147 112289 140175
rect 112323 140147 112351 140175
rect 112137 140085 112165 140113
rect 112199 140085 112227 140113
rect 112261 140085 112289 140113
rect 112323 140085 112351 140113
rect 112137 140023 112165 140051
rect 112199 140023 112227 140051
rect 112261 140023 112289 140051
rect 112323 140023 112351 140051
rect 112137 139961 112165 139989
rect 112199 139961 112227 139989
rect 112261 139961 112289 139989
rect 112323 139961 112351 139989
rect 123459 140147 123487 140175
rect 123521 140147 123549 140175
rect 123459 140085 123487 140113
rect 123521 140085 123549 140113
rect 123459 140023 123487 140051
rect 123521 140023 123549 140051
rect 123459 139961 123487 139989
rect 123521 139961 123549 139989
rect 115779 137147 115807 137175
rect 115841 137147 115869 137175
rect 115779 137085 115807 137113
rect 115841 137085 115869 137113
rect 115779 137023 115807 137051
rect 115841 137023 115869 137051
rect 115779 136961 115807 136989
rect 115841 136961 115869 136989
rect 125637 137147 125665 137175
rect 125699 137147 125727 137175
rect 125761 137147 125789 137175
rect 125823 137147 125851 137175
rect 125637 137085 125665 137113
rect 125699 137085 125727 137113
rect 125761 137085 125789 137113
rect 125823 137085 125851 137113
rect 125637 137023 125665 137051
rect 125699 137023 125727 137051
rect 125761 137023 125789 137051
rect 125823 137023 125851 137051
rect 125637 136961 125665 136989
rect 125699 136961 125727 136989
rect 125761 136961 125789 136989
rect 125823 136961 125851 136989
rect 112137 131147 112165 131175
rect 112199 131147 112227 131175
rect 112261 131147 112289 131175
rect 112323 131147 112351 131175
rect 112137 131085 112165 131113
rect 112199 131085 112227 131113
rect 112261 131085 112289 131113
rect 112323 131085 112351 131113
rect 112137 131023 112165 131051
rect 112199 131023 112227 131051
rect 112261 131023 112289 131051
rect 112323 131023 112351 131051
rect 112137 130961 112165 130989
rect 112199 130961 112227 130989
rect 112261 130961 112289 130989
rect 112323 130961 112351 130989
rect 123459 131147 123487 131175
rect 123521 131147 123549 131175
rect 123459 131085 123487 131113
rect 123521 131085 123549 131113
rect 123459 131023 123487 131051
rect 123521 131023 123549 131051
rect 123459 130961 123487 130989
rect 123521 130961 123549 130989
rect 115779 128147 115807 128175
rect 115841 128147 115869 128175
rect 115779 128085 115807 128113
rect 115841 128085 115869 128113
rect 115779 128023 115807 128051
rect 115841 128023 115869 128051
rect 115779 127961 115807 127989
rect 115841 127961 115869 127989
rect 125637 128147 125665 128175
rect 125699 128147 125727 128175
rect 125761 128147 125789 128175
rect 125823 128147 125851 128175
rect 125637 128085 125665 128113
rect 125699 128085 125727 128113
rect 125761 128085 125789 128113
rect 125823 128085 125851 128113
rect 125637 128023 125665 128051
rect 125699 128023 125727 128051
rect 125761 128023 125789 128051
rect 125823 128023 125851 128051
rect 125637 127961 125665 127989
rect 125699 127961 125727 127989
rect 125761 127961 125789 127989
rect 125823 127961 125851 127989
rect 112137 122147 112165 122175
rect 112199 122147 112227 122175
rect 112261 122147 112289 122175
rect 112323 122147 112351 122175
rect 112137 122085 112165 122113
rect 112199 122085 112227 122113
rect 112261 122085 112289 122113
rect 112323 122085 112351 122113
rect 112137 122023 112165 122051
rect 112199 122023 112227 122051
rect 112261 122023 112289 122051
rect 112323 122023 112351 122051
rect 112137 121961 112165 121989
rect 112199 121961 112227 121989
rect 112261 121961 112289 121989
rect 112323 121961 112351 121989
rect 123459 122147 123487 122175
rect 123521 122147 123549 122175
rect 123459 122085 123487 122113
rect 123521 122085 123549 122113
rect 123459 122023 123487 122051
rect 123521 122023 123549 122051
rect 123459 121961 123487 121989
rect 123521 121961 123549 121989
rect 115779 119147 115807 119175
rect 115841 119147 115869 119175
rect 115779 119085 115807 119113
rect 115841 119085 115869 119113
rect 115779 119023 115807 119051
rect 115841 119023 115869 119051
rect 115779 118961 115807 118989
rect 115841 118961 115869 118989
rect 125637 119147 125665 119175
rect 125699 119147 125727 119175
rect 125761 119147 125789 119175
rect 125823 119147 125851 119175
rect 125637 119085 125665 119113
rect 125699 119085 125727 119113
rect 125761 119085 125789 119113
rect 125823 119085 125851 119113
rect 125637 119023 125665 119051
rect 125699 119023 125727 119051
rect 125761 119023 125789 119051
rect 125823 119023 125851 119051
rect 125637 118961 125665 118989
rect 125699 118961 125727 118989
rect 125761 118961 125789 118989
rect 125823 118961 125851 118989
rect 112137 113147 112165 113175
rect 112199 113147 112227 113175
rect 112261 113147 112289 113175
rect 112323 113147 112351 113175
rect 112137 113085 112165 113113
rect 112199 113085 112227 113113
rect 112261 113085 112289 113113
rect 112323 113085 112351 113113
rect 112137 113023 112165 113051
rect 112199 113023 112227 113051
rect 112261 113023 112289 113051
rect 112323 113023 112351 113051
rect 112137 112961 112165 112989
rect 112199 112961 112227 112989
rect 112261 112961 112289 112989
rect 112323 112961 112351 112989
rect 123459 113147 123487 113175
rect 123521 113147 123549 113175
rect 123459 113085 123487 113113
rect 123521 113085 123549 113113
rect 123459 113023 123487 113051
rect 123521 113023 123549 113051
rect 123459 112961 123487 112989
rect 123521 112961 123549 112989
rect 115779 110147 115807 110175
rect 115841 110147 115869 110175
rect 115779 110085 115807 110113
rect 115841 110085 115869 110113
rect 115779 110023 115807 110051
rect 115841 110023 115869 110051
rect 115779 109961 115807 109989
rect 115841 109961 115869 109989
rect 125637 110147 125665 110175
rect 125699 110147 125727 110175
rect 125761 110147 125789 110175
rect 125823 110147 125851 110175
rect 125637 110085 125665 110113
rect 125699 110085 125727 110113
rect 125761 110085 125789 110113
rect 125823 110085 125851 110113
rect 125637 110023 125665 110051
rect 125699 110023 125727 110051
rect 125761 110023 125789 110051
rect 125823 110023 125851 110051
rect 125637 109961 125665 109989
rect 125699 109961 125727 109989
rect 125761 109961 125789 109989
rect 125823 109961 125851 109989
rect 112137 104147 112165 104175
rect 112199 104147 112227 104175
rect 112261 104147 112289 104175
rect 112323 104147 112351 104175
rect 112137 104085 112165 104113
rect 112199 104085 112227 104113
rect 112261 104085 112289 104113
rect 112323 104085 112351 104113
rect 112137 104023 112165 104051
rect 112199 104023 112227 104051
rect 112261 104023 112289 104051
rect 112323 104023 112351 104051
rect 112137 103961 112165 103989
rect 112199 103961 112227 103989
rect 112261 103961 112289 103989
rect 112323 103961 112351 103989
rect 123459 104147 123487 104175
rect 123521 104147 123549 104175
rect 123459 104085 123487 104113
rect 123521 104085 123549 104113
rect 123459 104023 123487 104051
rect 123521 104023 123549 104051
rect 123459 103961 123487 103989
rect 123521 103961 123549 103989
rect 115779 101147 115807 101175
rect 115841 101147 115869 101175
rect 115779 101085 115807 101113
rect 115841 101085 115869 101113
rect 115779 101023 115807 101051
rect 115841 101023 115869 101051
rect 115779 100961 115807 100989
rect 115841 100961 115869 100989
rect 125637 101147 125665 101175
rect 125699 101147 125727 101175
rect 125761 101147 125789 101175
rect 125823 101147 125851 101175
rect 125637 101085 125665 101113
rect 125699 101085 125727 101113
rect 125761 101085 125789 101113
rect 125823 101085 125851 101113
rect 125637 101023 125665 101051
rect 125699 101023 125727 101051
rect 125761 101023 125789 101051
rect 125823 101023 125851 101051
rect 125637 100961 125665 100989
rect 125699 100961 125727 100989
rect 125761 100961 125789 100989
rect 125823 100961 125851 100989
rect 112137 95147 112165 95175
rect 112199 95147 112227 95175
rect 112261 95147 112289 95175
rect 112323 95147 112351 95175
rect 112137 95085 112165 95113
rect 112199 95085 112227 95113
rect 112261 95085 112289 95113
rect 112323 95085 112351 95113
rect 112137 95023 112165 95051
rect 112199 95023 112227 95051
rect 112261 95023 112289 95051
rect 112323 95023 112351 95051
rect 112137 94961 112165 94989
rect 112199 94961 112227 94989
rect 112261 94961 112289 94989
rect 112323 94961 112351 94989
rect 123459 95147 123487 95175
rect 123521 95147 123549 95175
rect 123459 95085 123487 95113
rect 123521 95085 123549 95113
rect 123459 95023 123487 95051
rect 123521 95023 123549 95051
rect 123459 94961 123487 94989
rect 123521 94961 123549 94989
rect 115779 92147 115807 92175
rect 115841 92147 115869 92175
rect 115779 92085 115807 92113
rect 115841 92085 115869 92113
rect 115779 92023 115807 92051
rect 115841 92023 115869 92051
rect 115779 91961 115807 91989
rect 115841 91961 115869 91989
rect 125637 92147 125665 92175
rect 125699 92147 125727 92175
rect 125761 92147 125789 92175
rect 125823 92147 125851 92175
rect 125637 92085 125665 92113
rect 125699 92085 125727 92113
rect 125761 92085 125789 92113
rect 125823 92085 125851 92113
rect 125637 92023 125665 92051
rect 125699 92023 125727 92051
rect 125761 92023 125789 92051
rect 125823 92023 125851 92051
rect 125637 91961 125665 91989
rect 125699 91961 125727 91989
rect 125761 91961 125789 91989
rect 125823 91961 125851 91989
rect 112137 86147 112165 86175
rect 112199 86147 112227 86175
rect 112261 86147 112289 86175
rect 112323 86147 112351 86175
rect 112137 86085 112165 86113
rect 112199 86085 112227 86113
rect 112261 86085 112289 86113
rect 112323 86085 112351 86113
rect 112137 86023 112165 86051
rect 112199 86023 112227 86051
rect 112261 86023 112289 86051
rect 112323 86023 112351 86051
rect 112137 85961 112165 85989
rect 112199 85961 112227 85989
rect 112261 85961 112289 85989
rect 112323 85961 112351 85989
rect 123459 86147 123487 86175
rect 123521 86147 123549 86175
rect 123459 86085 123487 86113
rect 123521 86085 123549 86113
rect 123459 86023 123487 86051
rect 123521 86023 123549 86051
rect 123459 85961 123487 85989
rect 123521 85961 123549 85989
rect 115779 83147 115807 83175
rect 115841 83147 115869 83175
rect 115779 83085 115807 83113
rect 115841 83085 115869 83113
rect 115779 83023 115807 83051
rect 115841 83023 115869 83051
rect 115779 82961 115807 82989
rect 115841 82961 115869 82989
rect 125637 83147 125665 83175
rect 125699 83147 125727 83175
rect 125761 83147 125789 83175
rect 125823 83147 125851 83175
rect 125637 83085 125665 83113
rect 125699 83085 125727 83113
rect 125761 83085 125789 83113
rect 125823 83085 125851 83113
rect 125637 83023 125665 83051
rect 125699 83023 125727 83051
rect 125761 83023 125789 83051
rect 125823 83023 125851 83051
rect 125637 82961 125665 82989
rect 125699 82961 125727 82989
rect 125761 82961 125789 82989
rect 125823 82961 125851 82989
rect 112137 77147 112165 77175
rect 112199 77147 112227 77175
rect 112261 77147 112289 77175
rect 112323 77147 112351 77175
rect 112137 77085 112165 77113
rect 112199 77085 112227 77113
rect 112261 77085 112289 77113
rect 112323 77085 112351 77113
rect 112137 77023 112165 77051
rect 112199 77023 112227 77051
rect 112261 77023 112289 77051
rect 112323 77023 112351 77051
rect 112137 76961 112165 76989
rect 112199 76961 112227 76989
rect 112261 76961 112289 76989
rect 112323 76961 112351 76989
rect 123459 77147 123487 77175
rect 123521 77147 123549 77175
rect 123459 77085 123487 77113
rect 123521 77085 123549 77113
rect 123459 77023 123487 77051
rect 123521 77023 123549 77051
rect 123459 76961 123487 76989
rect 123521 76961 123549 76989
rect 115779 74147 115807 74175
rect 115841 74147 115869 74175
rect 115779 74085 115807 74113
rect 115841 74085 115869 74113
rect 115779 74023 115807 74051
rect 115841 74023 115869 74051
rect 115779 73961 115807 73989
rect 115841 73961 115869 73989
rect 125637 74147 125665 74175
rect 125699 74147 125727 74175
rect 125761 74147 125789 74175
rect 125823 74147 125851 74175
rect 125637 74085 125665 74113
rect 125699 74085 125727 74113
rect 125761 74085 125789 74113
rect 125823 74085 125851 74113
rect 125637 74023 125665 74051
rect 125699 74023 125727 74051
rect 125761 74023 125789 74051
rect 125823 74023 125851 74051
rect 125637 73961 125665 73989
rect 125699 73961 125727 73989
rect 125761 73961 125789 73989
rect 125823 73961 125851 73989
rect 112137 68147 112165 68175
rect 112199 68147 112227 68175
rect 112261 68147 112289 68175
rect 112323 68147 112351 68175
rect 112137 68085 112165 68113
rect 112199 68085 112227 68113
rect 112261 68085 112289 68113
rect 112323 68085 112351 68113
rect 112137 68023 112165 68051
rect 112199 68023 112227 68051
rect 112261 68023 112289 68051
rect 112323 68023 112351 68051
rect 112137 67961 112165 67989
rect 112199 67961 112227 67989
rect 112261 67961 112289 67989
rect 112323 67961 112351 67989
rect 123459 68147 123487 68175
rect 123521 68147 123549 68175
rect 123459 68085 123487 68113
rect 123521 68085 123549 68113
rect 123459 68023 123487 68051
rect 123521 68023 123549 68051
rect 123459 67961 123487 67989
rect 123521 67961 123549 67989
rect 115779 65147 115807 65175
rect 115841 65147 115869 65175
rect 115779 65085 115807 65113
rect 115841 65085 115869 65113
rect 115779 65023 115807 65051
rect 115841 65023 115869 65051
rect 115779 64961 115807 64989
rect 115841 64961 115869 64989
rect 125637 65147 125665 65175
rect 125699 65147 125727 65175
rect 125761 65147 125789 65175
rect 125823 65147 125851 65175
rect 125637 65085 125665 65113
rect 125699 65085 125727 65113
rect 125761 65085 125789 65113
rect 125823 65085 125851 65113
rect 125637 65023 125665 65051
rect 125699 65023 125727 65051
rect 125761 65023 125789 65051
rect 125823 65023 125851 65051
rect 125637 64961 125665 64989
rect 125699 64961 125727 64989
rect 125761 64961 125789 64989
rect 125823 64961 125851 64989
rect 112137 59147 112165 59175
rect 112199 59147 112227 59175
rect 112261 59147 112289 59175
rect 112323 59147 112351 59175
rect 112137 59085 112165 59113
rect 112199 59085 112227 59113
rect 112261 59085 112289 59113
rect 112323 59085 112351 59113
rect 112137 59023 112165 59051
rect 112199 59023 112227 59051
rect 112261 59023 112289 59051
rect 112323 59023 112351 59051
rect 112137 58961 112165 58989
rect 112199 58961 112227 58989
rect 112261 58961 112289 58989
rect 112323 58961 112351 58989
rect 123459 59147 123487 59175
rect 123521 59147 123549 59175
rect 123459 59085 123487 59113
rect 123521 59085 123549 59113
rect 123459 59023 123487 59051
rect 123521 59023 123549 59051
rect 123459 58961 123487 58989
rect 123521 58961 123549 58989
rect 115779 56147 115807 56175
rect 115841 56147 115869 56175
rect 115779 56085 115807 56113
rect 115841 56085 115869 56113
rect 115779 56023 115807 56051
rect 115841 56023 115869 56051
rect 115779 55961 115807 55989
rect 115841 55961 115869 55989
rect 125637 56147 125665 56175
rect 125699 56147 125727 56175
rect 125761 56147 125789 56175
rect 125823 56147 125851 56175
rect 125637 56085 125665 56113
rect 125699 56085 125727 56113
rect 125761 56085 125789 56113
rect 125823 56085 125851 56113
rect 125637 56023 125665 56051
rect 125699 56023 125727 56051
rect 125761 56023 125789 56051
rect 125823 56023 125851 56051
rect 125637 55961 125665 55989
rect 125699 55961 125727 55989
rect 125761 55961 125789 55989
rect 125823 55961 125851 55989
rect 112137 50147 112165 50175
rect 112199 50147 112227 50175
rect 112261 50147 112289 50175
rect 112323 50147 112351 50175
rect 112137 50085 112165 50113
rect 112199 50085 112227 50113
rect 112261 50085 112289 50113
rect 112323 50085 112351 50113
rect 112137 50023 112165 50051
rect 112199 50023 112227 50051
rect 112261 50023 112289 50051
rect 112323 50023 112351 50051
rect 112137 49961 112165 49989
rect 112199 49961 112227 49989
rect 112261 49961 112289 49989
rect 112323 49961 112351 49989
rect 123459 50147 123487 50175
rect 123521 50147 123549 50175
rect 123459 50085 123487 50113
rect 123521 50085 123549 50113
rect 123459 50023 123487 50051
rect 123521 50023 123549 50051
rect 123459 49961 123487 49989
rect 123521 49961 123549 49989
rect 115779 47147 115807 47175
rect 115841 47147 115869 47175
rect 115779 47085 115807 47113
rect 115841 47085 115869 47113
rect 115779 47023 115807 47051
rect 115841 47023 115869 47051
rect 115779 46961 115807 46989
rect 115841 46961 115869 46989
rect 125637 47147 125665 47175
rect 125699 47147 125727 47175
rect 125761 47147 125789 47175
rect 125823 47147 125851 47175
rect 125637 47085 125665 47113
rect 125699 47085 125727 47113
rect 125761 47085 125789 47113
rect 125823 47085 125851 47113
rect 125637 47023 125665 47051
rect 125699 47023 125727 47051
rect 125761 47023 125789 47051
rect 125823 47023 125851 47051
rect 125637 46961 125665 46989
rect 125699 46961 125727 46989
rect 125761 46961 125789 46989
rect 125823 46961 125851 46989
rect 112137 41147 112165 41175
rect 112199 41147 112227 41175
rect 112261 41147 112289 41175
rect 112323 41147 112351 41175
rect 112137 41085 112165 41113
rect 112199 41085 112227 41113
rect 112261 41085 112289 41113
rect 112323 41085 112351 41113
rect 112137 41023 112165 41051
rect 112199 41023 112227 41051
rect 112261 41023 112289 41051
rect 112323 41023 112351 41051
rect 112137 40961 112165 40989
rect 112199 40961 112227 40989
rect 112261 40961 112289 40989
rect 112323 40961 112351 40989
rect 123459 41147 123487 41175
rect 123521 41147 123549 41175
rect 123459 41085 123487 41113
rect 123521 41085 123549 41113
rect 123459 41023 123487 41051
rect 123521 41023 123549 41051
rect 123459 40961 123487 40989
rect 123521 40961 123549 40989
rect 115779 38147 115807 38175
rect 115841 38147 115869 38175
rect 115779 38085 115807 38113
rect 115841 38085 115869 38113
rect 115779 38023 115807 38051
rect 115841 38023 115869 38051
rect 115779 37961 115807 37989
rect 115841 37961 115869 37989
rect 125637 38147 125665 38175
rect 125699 38147 125727 38175
rect 125761 38147 125789 38175
rect 125823 38147 125851 38175
rect 125637 38085 125665 38113
rect 125699 38085 125727 38113
rect 125761 38085 125789 38113
rect 125823 38085 125851 38113
rect 125637 38023 125665 38051
rect 125699 38023 125727 38051
rect 125761 38023 125789 38051
rect 125823 38023 125851 38051
rect 125637 37961 125665 37989
rect 125699 37961 125727 37989
rect 125761 37961 125789 37989
rect 125823 37961 125851 37989
rect 112137 32147 112165 32175
rect 112199 32147 112227 32175
rect 112261 32147 112289 32175
rect 112323 32147 112351 32175
rect 112137 32085 112165 32113
rect 112199 32085 112227 32113
rect 112261 32085 112289 32113
rect 112323 32085 112351 32113
rect 112137 32023 112165 32051
rect 112199 32023 112227 32051
rect 112261 32023 112289 32051
rect 112323 32023 112351 32051
rect 112137 31961 112165 31989
rect 112199 31961 112227 31989
rect 112261 31961 112289 31989
rect 112323 31961 112351 31989
rect 123459 32147 123487 32175
rect 123521 32147 123549 32175
rect 123459 32085 123487 32113
rect 123521 32085 123549 32113
rect 123459 32023 123487 32051
rect 123521 32023 123549 32051
rect 123459 31961 123487 31989
rect 123521 31961 123549 31989
rect 115779 29147 115807 29175
rect 115841 29147 115869 29175
rect 115779 29085 115807 29113
rect 115841 29085 115869 29113
rect 115779 29023 115807 29051
rect 115841 29023 115869 29051
rect 115779 28961 115807 28989
rect 115841 28961 115869 28989
rect 125637 29147 125665 29175
rect 125699 29147 125727 29175
rect 125761 29147 125789 29175
rect 125823 29147 125851 29175
rect 125637 29085 125665 29113
rect 125699 29085 125727 29113
rect 125761 29085 125789 29113
rect 125823 29085 125851 29113
rect 125637 29023 125665 29051
rect 125699 29023 125727 29051
rect 125761 29023 125789 29051
rect 125823 29023 125851 29051
rect 125637 28961 125665 28989
rect 125699 28961 125727 28989
rect 125761 28961 125789 28989
rect 125823 28961 125851 28989
rect 112137 23147 112165 23175
rect 112199 23147 112227 23175
rect 112261 23147 112289 23175
rect 112323 23147 112351 23175
rect 112137 23085 112165 23113
rect 112199 23085 112227 23113
rect 112261 23085 112289 23113
rect 112323 23085 112351 23113
rect 112137 23023 112165 23051
rect 112199 23023 112227 23051
rect 112261 23023 112289 23051
rect 112323 23023 112351 23051
rect 112137 22961 112165 22989
rect 112199 22961 112227 22989
rect 112261 22961 112289 22989
rect 112323 22961 112351 22989
rect 123459 23147 123487 23175
rect 123521 23147 123549 23175
rect 123459 23085 123487 23113
rect 123521 23085 123549 23113
rect 123459 23023 123487 23051
rect 123521 23023 123549 23051
rect 123459 22961 123487 22989
rect 123521 22961 123549 22989
rect 115779 20147 115807 20175
rect 115841 20147 115869 20175
rect 115779 20085 115807 20113
rect 115841 20085 115869 20113
rect 115779 20023 115807 20051
rect 115841 20023 115869 20051
rect 115779 19961 115807 19989
rect 115841 19961 115869 19989
rect 125637 20147 125665 20175
rect 125699 20147 125727 20175
rect 125761 20147 125789 20175
rect 125823 20147 125851 20175
rect 125637 20085 125665 20113
rect 125699 20085 125727 20113
rect 125761 20085 125789 20113
rect 125823 20085 125851 20113
rect 125637 20023 125665 20051
rect 125699 20023 125727 20051
rect 125761 20023 125789 20051
rect 125823 20023 125851 20051
rect 125637 19961 125665 19989
rect 125699 19961 125727 19989
rect 125761 19961 125789 19989
rect 125823 19961 125851 19989
rect 112137 14147 112165 14175
rect 112199 14147 112227 14175
rect 112261 14147 112289 14175
rect 112323 14147 112351 14175
rect 112137 14085 112165 14113
rect 112199 14085 112227 14113
rect 112261 14085 112289 14113
rect 112323 14085 112351 14113
rect 112137 14023 112165 14051
rect 112199 14023 112227 14051
rect 112261 14023 112289 14051
rect 112323 14023 112351 14051
rect 112137 13961 112165 13989
rect 112199 13961 112227 13989
rect 112261 13961 112289 13989
rect 112323 13961 112351 13989
rect 123459 14147 123487 14175
rect 123521 14147 123549 14175
rect 123459 14085 123487 14113
rect 123521 14085 123549 14113
rect 123459 14023 123487 14051
rect 123521 14023 123549 14051
rect 123459 13961 123487 13989
rect 123521 13961 123549 13989
rect 115779 11147 115807 11175
rect 115841 11147 115869 11175
rect 115779 11085 115807 11113
rect 115841 11085 115869 11113
rect 115779 11023 115807 11051
rect 115841 11023 115869 11051
rect 115779 10961 115807 10989
rect 115841 10961 115869 10989
rect 125637 11147 125665 11175
rect 125699 11147 125727 11175
rect 125761 11147 125789 11175
rect 125823 11147 125851 11175
rect 125637 11085 125665 11113
rect 125699 11085 125727 11113
rect 125761 11085 125789 11113
rect 125823 11085 125851 11113
rect 125637 11023 125665 11051
rect 125699 11023 125727 11051
rect 125761 11023 125789 11051
rect 125823 11023 125851 11051
rect 125637 10961 125665 10989
rect 125699 10961 125727 10989
rect 125761 10961 125789 10989
rect 125823 10961 125851 10989
rect 112137 5147 112165 5175
rect 112199 5147 112227 5175
rect 112261 5147 112289 5175
rect 112323 5147 112351 5175
rect 112137 5085 112165 5113
rect 112199 5085 112227 5113
rect 112261 5085 112289 5113
rect 112323 5085 112351 5113
rect 112137 5023 112165 5051
rect 112199 5023 112227 5051
rect 112261 5023 112289 5051
rect 112323 5023 112351 5051
rect 112137 4961 112165 4989
rect 112199 4961 112227 4989
rect 112261 4961 112289 4989
rect 112323 4961 112351 4989
rect 123459 5147 123487 5175
rect 123521 5147 123549 5175
rect 123459 5085 123487 5113
rect 123521 5085 123549 5113
rect 123459 5023 123487 5051
rect 123521 5023 123549 5051
rect 123459 4961 123487 4989
rect 123521 4961 123549 4989
rect 112137 -588 112165 -560
rect 112199 -588 112227 -560
rect 112261 -588 112289 -560
rect 112323 -588 112351 -560
rect 112137 -650 112165 -622
rect 112199 -650 112227 -622
rect 112261 -650 112289 -622
rect 112323 -650 112351 -622
rect 112137 -712 112165 -684
rect 112199 -712 112227 -684
rect 112261 -712 112289 -684
rect 112323 -712 112351 -684
rect 112137 -774 112165 -746
rect 112199 -774 112227 -746
rect 112261 -774 112289 -746
rect 112323 -774 112351 -746
rect 125637 2147 125665 2175
rect 125699 2147 125727 2175
rect 125761 2147 125789 2175
rect 125823 2147 125851 2175
rect 125637 2085 125665 2113
rect 125699 2085 125727 2113
rect 125761 2085 125789 2113
rect 125823 2085 125851 2113
rect 125637 2023 125665 2051
rect 125699 2023 125727 2051
rect 125761 2023 125789 2051
rect 125823 2023 125851 2051
rect 125637 1961 125665 1989
rect 125699 1961 125727 1989
rect 125761 1961 125789 1989
rect 125823 1961 125851 1989
rect 125637 -108 125665 -80
rect 125699 -108 125727 -80
rect 125761 -108 125789 -80
rect 125823 -108 125851 -80
rect 125637 -170 125665 -142
rect 125699 -170 125727 -142
rect 125761 -170 125789 -142
rect 125823 -170 125851 -142
rect 125637 -232 125665 -204
rect 125699 -232 125727 -204
rect 125761 -232 125789 -204
rect 125823 -232 125851 -204
rect 125637 -294 125665 -266
rect 125699 -294 125727 -266
rect 125761 -294 125789 -266
rect 125823 -294 125851 -266
rect 127497 299058 127525 299086
rect 127559 299058 127587 299086
rect 127621 299058 127649 299086
rect 127683 299058 127711 299086
rect 127497 298996 127525 299024
rect 127559 298996 127587 299024
rect 127621 298996 127649 299024
rect 127683 298996 127711 299024
rect 127497 298934 127525 298962
rect 127559 298934 127587 298962
rect 127621 298934 127649 298962
rect 127683 298934 127711 298962
rect 127497 298872 127525 298900
rect 127559 298872 127587 298900
rect 127621 298872 127649 298900
rect 127683 298872 127711 298900
rect 127497 293147 127525 293175
rect 127559 293147 127587 293175
rect 127621 293147 127649 293175
rect 127683 293147 127711 293175
rect 127497 293085 127525 293113
rect 127559 293085 127587 293113
rect 127621 293085 127649 293113
rect 127683 293085 127711 293113
rect 127497 293023 127525 293051
rect 127559 293023 127587 293051
rect 127621 293023 127649 293051
rect 127683 293023 127711 293051
rect 127497 292961 127525 292989
rect 127559 292961 127587 292989
rect 127621 292961 127649 292989
rect 127683 292961 127711 292989
rect 127497 284147 127525 284175
rect 127559 284147 127587 284175
rect 127621 284147 127649 284175
rect 127683 284147 127711 284175
rect 127497 284085 127525 284113
rect 127559 284085 127587 284113
rect 127621 284085 127649 284113
rect 127683 284085 127711 284113
rect 127497 284023 127525 284051
rect 127559 284023 127587 284051
rect 127621 284023 127649 284051
rect 127683 284023 127711 284051
rect 127497 283961 127525 283989
rect 127559 283961 127587 283989
rect 127621 283961 127649 283989
rect 127683 283961 127711 283989
rect 127497 275147 127525 275175
rect 127559 275147 127587 275175
rect 127621 275147 127649 275175
rect 127683 275147 127711 275175
rect 127497 275085 127525 275113
rect 127559 275085 127587 275113
rect 127621 275085 127649 275113
rect 127683 275085 127711 275113
rect 127497 275023 127525 275051
rect 127559 275023 127587 275051
rect 127621 275023 127649 275051
rect 127683 275023 127711 275051
rect 127497 274961 127525 274989
rect 127559 274961 127587 274989
rect 127621 274961 127649 274989
rect 127683 274961 127711 274989
rect 127497 266147 127525 266175
rect 127559 266147 127587 266175
rect 127621 266147 127649 266175
rect 127683 266147 127711 266175
rect 127497 266085 127525 266113
rect 127559 266085 127587 266113
rect 127621 266085 127649 266113
rect 127683 266085 127711 266113
rect 127497 266023 127525 266051
rect 127559 266023 127587 266051
rect 127621 266023 127649 266051
rect 127683 266023 127711 266051
rect 127497 265961 127525 265989
rect 127559 265961 127587 265989
rect 127621 265961 127649 265989
rect 127683 265961 127711 265989
rect 127497 257147 127525 257175
rect 127559 257147 127587 257175
rect 127621 257147 127649 257175
rect 127683 257147 127711 257175
rect 127497 257085 127525 257113
rect 127559 257085 127587 257113
rect 127621 257085 127649 257113
rect 127683 257085 127711 257113
rect 127497 257023 127525 257051
rect 127559 257023 127587 257051
rect 127621 257023 127649 257051
rect 127683 257023 127711 257051
rect 127497 256961 127525 256989
rect 127559 256961 127587 256989
rect 127621 256961 127649 256989
rect 127683 256961 127711 256989
rect 127497 248147 127525 248175
rect 127559 248147 127587 248175
rect 127621 248147 127649 248175
rect 127683 248147 127711 248175
rect 127497 248085 127525 248113
rect 127559 248085 127587 248113
rect 127621 248085 127649 248113
rect 127683 248085 127711 248113
rect 127497 248023 127525 248051
rect 127559 248023 127587 248051
rect 127621 248023 127649 248051
rect 127683 248023 127711 248051
rect 127497 247961 127525 247989
rect 127559 247961 127587 247989
rect 127621 247961 127649 247989
rect 127683 247961 127711 247989
rect 127497 239147 127525 239175
rect 127559 239147 127587 239175
rect 127621 239147 127649 239175
rect 127683 239147 127711 239175
rect 127497 239085 127525 239113
rect 127559 239085 127587 239113
rect 127621 239085 127649 239113
rect 127683 239085 127711 239113
rect 127497 239023 127525 239051
rect 127559 239023 127587 239051
rect 127621 239023 127649 239051
rect 127683 239023 127711 239051
rect 127497 238961 127525 238989
rect 127559 238961 127587 238989
rect 127621 238961 127649 238989
rect 127683 238961 127711 238989
rect 127497 230147 127525 230175
rect 127559 230147 127587 230175
rect 127621 230147 127649 230175
rect 127683 230147 127711 230175
rect 127497 230085 127525 230113
rect 127559 230085 127587 230113
rect 127621 230085 127649 230113
rect 127683 230085 127711 230113
rect 127497 230023 127525 230051
rect 127559 230023 127587 230051
rect 127621 230023 127649 230051
rect 127683 230023 127711 230051
rect 127497 229961 127525 229989
rect 127559 229961 127587 229989
rect 127621 229961 127649 229989
rect 127683 229961 127711 229989
rect 127497 221147 127525 221175
rect 127559 221147 127587 221175
rect 127621 221147 127649 221175
rect 127683 221147 127711 221175
rect 127497 221085 127525 221113
rect 127559 221085 127587 221113
rect 127621 221085 127649 221113
rect 127683 221085 127711 221113
rect 127497 221023 127525 221051
rect 127559 221023 127587 221051
rect 127621 221023 127649 221051
rect 127683 221023 127711 221051
rect 127497 220961 127525 220989
rect 127559 220961 127587 220989
rect 127621 220961 127649 220989
rect 127683 220961 127711 220989
rect 127497 212147 127525 212175
rect 127559 212147 127587 212175
rect 127621 212147 127649 212175
rect 127683 212147 127711 212175
rect 127497 212085 127525 212113
rect 127559 212085 127587 212113
rect 127621 212085 127649 212113
rect 127683 212085 127711 212113
rect 127497 212023 127525 212051
rect 127559 212023 127587 212051
rect 127621 212023 127649 212051
rect 127683 212023 127711 212051
rect 127497 211961 127525 211989
rect 127559 211961 127587 211989
rect 127621 211961 127649 211989
rect 127683 211961 127711 211989
rect 127497 203147 127525 203175
rect 127559 203147 127587 203175
rect 127621 203147 127649 203175
rect 127683 203147 127711 203175
rect 127497 203085 127525 203113
rect 127559 203085 127587 203113
rect 127621 203085 127649 203113
rect 127683 203085 127711 203113
rect 127497 203023 127525 203051
rect 127559 203023 127587 203051
rect 127621 203023 127649 203051
rect 127683 203023 127711 203051
rect 127497 202961 127525 202989
rect 127559 202961 127587 202989
rect 127621 202961 127649 202989
rect 127683 202961 127711 202989
rect 127497 194147 127525 194175
rect 127559 194147 127587 194175
rect 127621 194147 127649 194175
rect 127683 194147 127711 194175
rect 127497 194085 127525 194113
rect 127559 194085 127587 194113
rect 127621 194085 127649 194113
rect 127683 194085 127711 194113
rect 127497 194023 127525 194051
rect 127559 194023 127587 194051
rect 127621 194023 127649 194051
rect 127683 194023 127711 194051
rect 127497 193961 127525 193989
rect 127559 193961 127587 193989
rect 127621 193961 127649 193989
rect 127683 193961 127711 193989
rect 127497 185147 127525 185175
rect 127559 185147 127587 185175
rect 127621 185147 127649 185175
rect 127683 185147 127711 185175
rect 127497 185085 127525 185113
rect 127559 185085 127587 185113
rect 127621 185085 127649 185113
rect 127683 185085 127711 185113
rect 127497 185023 127525 185051
rect 127559 185023 127587 185051
rect 127621 185023 127649 185051
rect 127683 185023 127711 185051
rect 127497 184961 127525 184989
rect 127559 184961 127587 184989
rect 127621 184961 127649 184989
rect 127683 184961 127711 184989
rect 127497 176147 127525 176175
rect 127559 176147 127587 176175
rect 127621 176147 127649 176175
rect 127683 176147 127711 176175
rect 127497 176085 127525 176113
rect 127559 176085 127587 176113
rect 127621 176085 127649 176113
rect 127683 176085 127711 176113
rect 127497 176023 127525 176051
rect 127559 176023 127587 176051
rect 127621 176023 127649 176051
rect 127683 176023 127711 176051
rect 127497 175961 127525 175989
rect 127559 175961 127587 175989
rect 127621 175961 127649 175989
rect 127683 175961 127711 175989
rect 140997 298578 141025 298606
rect 141059 298578 141087 298606
rect 141121 298578 141149 298606
rect 141183 298578 141211 298606
rect 140997 298516 141025 298544
rect 141059 298516 141087 298544
rect 141121 298516 141149 298544
rect 141183 298516 141211 298544
rect 140997 298454 141025 298482
rect 141059 298454 141087 298482
rect 141121 298454 141149 298482
rect 141183 298454 141211 298482
rect 140997 298392 141025 298420
rect 141059 298392 141087 298420
rect 141121 298392 141149 298420
rect 141183 298392 141211 298420
rect 140997 290147 141025 290175
rect 141059 290147 141087 290175
rect 141121 290147 141149 290175
rect 141183 290147 141211 290175
rect 140997 290085 141025 290113
rect 141059 290085 141087 290113
rect 141121 290085 141149 290113
rect 141183 290085 141211 290113
rect 140997 290023 141025 290051
rect 141059 290023 141087 290051
rect 141121 290023 141149 290051
rect 141183 290023 141211 290051
rect 140997 289961 141025 289989
rect 141059 289961 141087 289989
rect 141121 289961 141149 289989
rect 141183 289961 141211 289989
rect 140997 281147 141025 281175
rect 141059 281147 141087 281175
rect 141121 281147 141149 281175
rect 141183 281147 141211 281175
rect 140997 281085 141025 281113
rect 141059 281085 141087 281113
rect 141121 281085 141149 281113
rect 141183 281085 141211 281113
rect 140997 281023 141025 281051
rect 141059 281023 141087 281051
rect 141121 281023 141149 281051
rect 141183 281023 141211 281051
rect 140997 280961 141025 280989
rect 141059 280961 141087 280989
rect 141121 280961 141149 280989
rect 141183 280961 141211 280989
rect 140997 272147 141025 272175
rect 141059 272147 141087 272175
rect 141121 272147 141149 272175
rect 141183 272147 141211 272175
rect 140997 272085 141025 272113
rect 141059 272085 141087 272113
rect 141121 272085 141149 272113
rect 141183 272085 141211 272113
rect 140997 272023 141025 272051
rect 141059 272023 141087 272051
rect 141121 272023 141149 272051
rect 141183 272023 141211 272051
rect 140997 271961 141025 271989
rect 141059 271961 141087 271989
rect 141121 271961 141149 271989
rect 141183 271961 141211 271989
rect 140997 263147 141025 263175
rect 141059 263147 141087 263175
rect 141121 263147 141149 263175
rect 141183 263147 141211 263175
rect 140997 263085 141025 263113
rect 141059 263085 141087 263113
rect 141121 263085 141149 263113
rect 141183 263085 141211 263113
rect 140997 263023 141025 263051
rect 141059 263023 141087 263051
rect 141121 263023 141149 263051
rect 141183 263023 141211 263051
rect 140997 262961 141025 262989
rect 141059 262961 141087 262989
rect 141121 262961 141149 262989
rect 141183 262961 141211 262989
rect 140997 254147 141025 254175
rect 141059 254147 141087 254175
rect 141121 254147 141149 254175
rect 141183 254147 141211 254175
rect 140997 254085 141025 254113
rect 141059 254085 141087 254113
rect 141121 254085 141149 254113
rect 141183 254085 141211 254113
rect 140997 254023 141025 254051
rect 141059 254023 141087 254051
rect 141121 254023 141149 254051
rect 141183 254023 141211 254051
rect 140997 253961 141025 253989
rect 141059 253961 141087 253989
rect 141121 253961 141149 253989
rect 141183 253961 141211 253989
rect 140997 245147 141025 245175
rect 141059 245147 141087 245175
rect 141121 245147 141149 245175
rect 141183 245147 141211 245175
rect 140997 245085 141025 245113
rect 141059 245085 141087 245113
rect 141121 245085 141149 245113
rect 141183 245085 141211 245113
rect 140997 245023 141025 245051
rect 141059 245023 141087 245051
rect 141121 245023 141149 245051
rect 141183 245023 141211 245051
rect 140997 244961 141025 244989
rect 141059 244961 141087 244989
rect 141121 244961 141149 244989
rect 141183 244961 141211 244989
rect 140997 236147 141025 236175
rect 141059 236147 141087 236175
rect 141121 236147 141149 236175
rect 141183 236147 141211 236175
rect 140997 236085 141025 236113
rect 141059 236085 141087 236113
rect 141121 236085 141149 236113
rect 141183 236085 141211 236113
rect 140997 236023 141025 236051
rect 141059 236023 141087 236051
rect 141121 236023 141149 236051
rect 141183 236023 141211 236051
rect 140997 235961 141025 235989
rect 141059 235961 141087 235989
rect 141121 235961 141149 235989
rect 141183 235961 141211 235989
rect 140997 227147 141025 227175
rect 141059 227147 141087 227175
rect 141121 227147 141149 227175
rect 141183 227147 141211 227175
rect 140997 227085 141025 227113
rect 141059 227085 141087 227113
rect 141121 227085 141149 227113
rect 141183 227085 141211 227113
rect 140997 227023 141025 227051
rect 141059 227023 141087 227051
rect 141121 227023 141149 227051
rect 141183 227023 141211 227051
rect 140997 226961 141025 226989
rect 141059 226961 141087 226989
rect 141121 226961 141149 226989
rect 141183 226961 141211 226989
rect 140997 218147 141025 218175
rect 141059 218147 141087 218175
rect 141121 218147 141149 218175
rect 141183 218147 141211 218175
rect 140997 218085 141025 218113
rect 141059 218085 141087 218113
rect 141121 218085 141149 218113
rect 141183 218085 141211 218113
rect 140997 218023 141025 218051
rect 141059 218023 141087 218051
rect 141121 218023 141149 218051
rect 141183 218023 141211 218051
rect 140997 217961 141025 217989
rect 141059 217961 141087 217989
rect 141121 217961 141149 217989
rect 141183 217961 141211 217989
rect 140997 209147 141025 209175
rect 141059 209147 141087 209175
rect 141121 209147 141149 209175
rect 141183 209147 141211 209175
rect 140997 209085 141025 209113
rect 141059 209085 141087 209113
rect 141121 209085 141149 209113
rect 141183 209085 141211 209113
rect 140997 209023 141025 209051
rect 141059 209023 141087 209051
rect 141121 209023 141149 209051
rect 141183 209023 141211 209051
rect 140997 208961 141025 208989
rect 141059 208961 141087 208989
rect 141121 208961 141149 208989
rect 141183 208961 141211 208989
rect 140997 200147 141025 200175
rect 141059 200147 141087 200175
rect 141121 200147 141149 200175
rect 141183 200147 141211 200175
rect 140997 200085 141025 200113
rect 141059 200085 141087 200113
rect 141121 200085 141149 200113
rect 141183 200085 141211 200113
rect 140997 200023 141025 200051
rect 141059 200023 141087 200051
rect 141121 200023 141149 200051
rect 141183 200023 141211 200051
rect 140997 199961 141025 199989
rect 141059 199961 141087 199989
rect 141121 199961 141149 199989
rect 141183 199961 141211 199989
rect 140997 191147 141025 191175
rect 141059 191147 141087 191175
rect 141121 191147 141149 191175
rect 141183 191147 141211 191175
rect 140997 191085 141025 191113
rect 141059 191085 141087 191113
rect 141121 191085 141149 191113
rect 141183 191085 141211 191113
rect 140997 191023 141025 191051
rect 141059 191023 141087 191051
rect 141121 191023 141149 191051
rect 141183 191023 141211 191051
rect 140997 190961 141025 190989
rect 141059 190961 141087 190989
rect 141121 190961 141149 190989
rect 141183 190961 141211 190989
rect 140997 182147 141025 182175
rect 141059 182147 141087 182175
rect 141121 182147 141149 182175
rect 141183 182147 141211 182175
rect 140997 182085 141025 182113
rect 141059 182085 141087 182113
rect 141121 182085 141149 182113
rect 141183 182085 141211 182113
rect 140997 182023 141025 182051
rect 141059 182023 141087 182051
rect 141121 182023 141149 182051
rect 141183 182023 141211 182051
rect 140997 181961 141025 181989
rect 141059 181961 141087 181989
rect 141121 181961 141149 181989
rect 141183 181961 141211 181989
rect 131139 173147 131167 173175
rect 131201 173147 131229 173175
rect 131139 173085 131167 173113
rect 131201 173085 131229 173113
rect 131139 173023 131167 173051
rect 131201 173023 131229 173051
rect 131139 172961 131167 172989
rect 131201 172961 131229 172989
rect 140997 173147 141025 173175
rect 141059 173147 141087 173175
rect 141121 173147 141149 173175
rect 141183 173147 141211 173175
rect 140997 173085 141025 173113
rect 141059 173085 141087 173113
rect 141121 173085 141149 173113
rect 141183 173085 141211 173113
rect 140997 173023 141025 173051
rect 141059 173023 141087 173051
rect 141121 173023 141149 173051
rect 141183 173023 141211 173051
rect 140997 172961 141025 172989
rect 141059 172961 141087 172989
rect 141121 172961 141149 172989
rect 141183 172961 141211 172989
rect 127497 167147 127525 167175
rect 127559 167147 127587 167175
rect 127621 167147 127649 167175
rect 127683 167147 127711 167175
rect 127497 167085 127525 167113
rect 127559 167085 127587 167113
rect 127621 167085 127649 167113
rect 127683 167085 127711 167113
rect 127497 167023 127525 167051
rect 127559 167023 127587 167051
rect 127621 167023 127649 167051
rect 127683 167023 127711 167051
rect 127497 166961 127525 166989
rect 127559 166961 127587 166989
rect 127621 166961 127649 166989
rect 127683 166961 127711 166989
rect 138819 167147 138847 167175
rect 138881 167147 138909 167175
rect 138819 167085 138847 167113
rect 138881 167085 138909 167113
rect 138819 167023 138847 167051
rect 138881 167023 138909 167051
rect 138819 166961 138847 166989
rect 138881 166961 138909 166989
rect 131139 164147 131167 164175
rect 131201 164147 131229 164175
rect 131139 164085 131167 164113
rect 131201 164085 131229 164113
rect 131139 164023 131167 164051
rect 131201 164023 131229 164051
rect 131139 163961 131167 163989
rect 131201 163961 131229 163989
rect 140997 164147 141025 164175
rect 141059 164147 141087 164175
rect 141121 164147 141149 164175
rect 141183 164147 141211 164175
rect 140997 164085 141025 164113
rect 141059 164085 141087 164113
rect 141121 164085 141149 164113
rect 141183 164085 141211 164113
rect 140997 164023 141025 164051
rect 141059 164023 141087 164051
rect 141121 164023 141149 164051
rect 141183 164023 141211 164051
rect 140997 163961 141025 163989
rect 141059 163961 141087 163989
rect 141121 163961 141149 163989
rect 141183 163961 141211 163989
rect 127497 158147 127525 158175
rect 127559 158147 127587 158175
rect 127621 158147 127649 158175
rect 127683 158147 127711 158175
rect 127497 158085 127525 158113
rect 127559 158085 127587 158113
rect 127621 158085 127649 158113
rect 127683 158085 127711 158113
rect 127497 158023 127525 158051
rect 127559 158023 127587 158051
rect 127621 158023 127649 158051
rect 127683 158023 127711 158051
rect 127497 157961 127525 157989
rect 127559 157961 127587 157989
rect 127621 157961 127649 157989
rect 127683 157961 127711 157989
rect 138819 158147 138847 158175
rect 138881 158147 138909 158175
rect 138819 158085 138847 158113
rect 138881 158085 138909 158113
rect 138819 158023 138847 158051
rect 138881 158023 138909 158051
rect 138819 157961 138847 157989
rect 138881 157961 138909 157989
rect 131139 155147 131167 155175
rect 131201 155147 131229 155175
rect 131139 155085 131167 155113
rect 131201 155085 131229 155113
rect 131139 155023 131167 155051
rect 131201 155023 131229 155051
rect 131139 154961 131167 154989
rect 131201 154961 131229 154989
rect 140997 155147 141025 155175
rect 141059 155147 141087 155175
rect 141121 155147 141149 155175
rect 141183 155147 141211 155175
rect 140997 155085 141025 155113
rect 141059 155085 141087 155113
rect 141121 155085 141149 155113
rect 141183 155085 141211 155113
rect 140997 155023 141025 155051
rect 141059 155023 141087 155051
rect 141121 155023 141149 155051
rect 141183 155023 141211 155051
rect 140997 154961 141025 154989
rect 141059 154961 141087 154989
rect 141121 154961 141149 154989
rect 141183 154961 141211 154989
rect 127497 149147 127525 149175
rect 127559 149147 127587 149175
rect 127621 149147 127649 149175
rect 127683 149147 127711 149175
rect 127497 149085 127525 149113
rect 127559 149085 127587 149113
rect 127621 149085 127649 149113
rect 127683 149085 127711 149113
rect 127497 149023 127525 149051
rect 127559 149023 127587 149051
rect 127621 149023 127649 149051
rect 127683 149023 127711 149051
rect 127497 148961 127525 148989
rect 127559 148961 127587 148989
rect 127621 148961 127649 148989
rect 127683 148961 127711 148989
rect 138819 149147 138847 149175
rect 138881 149147 138909 149175
rect 138819 149085 138847 149113
rect 138881 149085 138909 149113
rect 138819 149023 138847 149051
rect 138881 149023 138909 149051
rect 138819 148961 138847 148989
rect 138881 148961 138909 148989
rect 131139 146147 131167 146175
rect 131201 146147 131229 146175
rect 131139 146085 131167 146113
rect 131201 146085 131229 146113
rect 131139 146023 131167 146051
rect 131201 146023 131229 146051
rect 131139 145961 131167 145989
rect 131201 145961 131229 145989
rect 140997 146147 141025 146175
rect 141059 146147 141087 146175
rect 141121 146147 141149 146175
rect 141183 146147 141211 146175
rect 140997 146085 141025 146113
rect 141059 146085 141087 146113
rect 141121 146085 141149 146113
rect 141183 146085 141211 146113
rect 140997 146023 141025 146051
rect 141059 146023 141087 146051
rect 141121 146023 141149 146051
rect 141183 146023 141211 146051
rect 140997 145961 141025 145989
rect 141059 145961 141087 145989
rect 141121 145961 141149 145989
rect 141183 145961 141211 145989
rect 127497 140147 127525 140175
rect 127559 140147 127587 140175
rect 127621 140147 127649 140175
rect 127683 140147 127711 140175
rect 127497 140085 127525 140113
rect 127559 140085 127587 140113
rect 127621 140085 127649 140113
rect 127683 140085 127711 140113
rect 127497 140023 127525 140051
rect 127559 140023 127587 140051
rect 127621 140023 127649 140051
rect 127683 140023 127711 140051
rect 127497 139961 127525 139989
rect 127559 139961 127587 139989
rect 127621 139961 127649 139989
rect 127683 139961 127711 139989
rect 138819 140147 138847 140175
rect 138881 140147 138909 140175
rect 138819 140085 138847 140113
rect 138881 140085 138909 140113
rect 138819 140023 138847 140051
rect 138881 140023 138909 140051
rect 138819 139961 138847 139989
rect 138881 139961 138909 139989
rect 131139 137147 131167 137175
rect 131201 137147 131229 137175
rect 131139 137085 131167 137113
rect 131201 137085 131229 137113
rect 131139 137023 131167 137051
rect 131201 137023 131229 137051
rect 131139 136961 131167 136989
rect 131201 136961 131229 136989
rect 140997 137147 141025 137175
rect 141059 137147 141087 137175
rect 141121 137147 141149 137175
rect 141183 137147 141211 137175
rect 140997 137085 141025 137113
rect 141059 137085 141087 137113
rect 141121 137085 141149 137113
rect 141183 137085 141211 137113
rect 140997 137023 141025 137051
rect 141059 137023 141087 137051
rect 141121 137023 141149 137051
rect 141183 137023 141211 137051
rect 140997 136961 141025 136989
rect 141059 136961 141087 136989
rect 141121 136961 141149 136989
rect 141183 136961 141211 136989
rect 127497 131147 127525 131175
rect 127559 131147 127587 131175
rect 127621 131147 127649 131175
rect 127683 131147 127711 131175
rect 127497 131085 127525 131113
rect 127559 131085 127587 131113
rect 127621 131085 127649 131113
rect 127683 131085 127711 131113
rect 127497 131023 127525 131051
rect 127559 131023 127587 131051
rect 127621 131023 127649 131051
rect 127683 131023 127711 131051
rect 127497 130961 127525 130989
rect 127559 130961 127587 130989
rect 127621 130961 127649 130989
rect 127683 130961 127711 130989
rect 138819 131147 138847 131175
rect 138881 131147 138909 131175
rect 138819 131085 138847 131113
rect 138881 131085 138909 131113
rect 138819 131023 138847 131051
rect 138881 131023 138909 131051
rect 138819 130961 138847 130989
rect 138881 130961 138909 130989
rect 131139 128147 131167 128175
rect 131201 128147 131229 128175
rect 131139 128085 131167 128113
rect 131201 128085 131229 128113
rect 131139 128023 131167 128051
rect 131201 128023 131229 128051
rect 131139 127961 131167 127989
rect 131201 127961 131229 127989
rect 140997 128147 141025 128175
rect 141059 128147 141087 128175
rect 141121 128147 141149 128175
rect 141183 128147 141211 128175
rect 140997 128085 141025 128113
rect 141059 128085 141087 128113
rect 141121 128085 141149 128113
rect 141183 128085 141211 128113
rect 140997 128023 141025 128051
rect 141059 128023 141087 128051
rect 141121 128023 141149 128051
rect 141183 128023 141211 128051
rect 140997 127961 141025 127989
rect 141059 127961 141087 127989
rect 141121 127961 141149 127989
rect 141183 127961 141211 127989
rect 127497 122147 127525 122175
rect 127559 122147 127587 122175
rect 127621 122147 127649 122175
rect 127683 122147 127711 122175
rect 127497 122085 127525 122113
rect 127559 122085 127587 122113
rect 127621 122085 127649 122113
rect 127683 122085 127711 122113
rect 127497 122023 127525 122051
rect 127559 122023 127587 122051
rect 127621 122023 127649 122051
rect 127683 122023 127711 122051
rect 127497 121961 127525 121989
rect 127559 121961 127587 121989
rect 127621 121961 127649 121989
rect 127683 121961 127711 121989
rect 138819 122147 138847 122175
rect 138881 122147 138909 122175
rect 138819 122085 138847 122113
rect 138881 122085 138909 122113
rect 138819 122023 138847 122051
rect 138881 122023 138909 122051
rect 138819 121961 138847 121989
rect 138881 121961 138909 121989
rect 131139 119147 131167 119175
rect 131201 119147 131229 119175
rect 131139 119085 131167 119113
rect 131201 119085 131229 119113
rect 131139 119023 131167 119051
rect 131201 119023 131229 119051
rect 131139 118961 131167 118989
rect 131201 118961 131229 118989
rect 140997 119147 141025 119175
rect 141059 119147 141087 119175
rect 141121 119147 141149 119175
rect 141183 119147 141211 119175
rect 140997 119085 141025 119113
rect 141059 119085 141087 119113
rect 141121 119085 141149 119113
rect 141183 119085 141211 119113
rect 140997 119023 141025 119051
rect 141059 119023 141087 119051
rect 141121 119023 141149 119051
rect 141183 119023 141211 119051
rect 140997 118961 141025 118989
rect 141059 118961 141087 118989
rect 141121 118961 141149 118989
rect 141183 118961 141211 118989
rect 127497 113147 127525 113175
rect 127559 113147 127587 113175
rect 127621 113147 127649 113175
rect 127683 113147 127711 113175
rect 127497 113085 127525 113113
rect 127559 113085 127587 113113
rect 127621 113085 127649 113113
rect 127683 113085 127711 113113
rect 127497 113023 127525 113051
rect 127559 113023 127587 113051
rect 127621 113023 127649 113051
rect 127683 113023 127711 113051
rect 127497 112961 127525 112989
rect 127559 112961 127587 112989
rect 127621 112961 127649 112989
rect 127683 112961 127711 112989
rect 138819 113147 138847 113175
rect 138881 113147 138909 113175
rect 138819 113085 138847 113113
rect 138881 113085 138909 113113
rect 138819 113023 138847 113051
rect 138881 113023 138909 113051
rect 138819 112961 138847 112989
rect 138881 112961 138909 112989
rect 131139 110147 131167 110175
rect 131201 110147 131229 110175
rect 131139 110085 131167 110113
rect 131201 110085 131229 110113
rect 131139 110023 131167 110051
rect 131201 110023 131229 110051
rect 131139 109961 131167 109989
rect 131201 109961 131229 109989
rect 140997 110147 141025 110175
rect 141059 110147 141087 110175
rect 141121 110147 141149 110175
rect 141183 110147 141211 110175
rect 140997 110085 141025 110113
rect 141059 110085 141087 110113
rect 141121 110085 141149 110113
rect 141183 110085 141211 110113
rect 140997 110023 141025 110051
rect 141059 110023 141087 110051
rect 141121 110023 141149 110051
rect 141183 110023 141211 110051
rect 140997 109961 141025 109989
rect 141059 109961 141087 109989
rect 141121 109961 141149 109989
rect 141183 109961 141211 109989
rect 127497 104147 127525 104175
rect 127559 104147 127587 104175
rect 127621 104147 127649 104175
rect 127683 104147 127711 104175
rect 127497 104085 127525 104113
rect 127559 104085 127587 104113
rect 127621 104085 127649 104113
rect 127683 104085 127711 104113
rect 127497 104023 127525 104051
rect 127559 104023 127587 104051
rect 127621 104023 127649 104051
rect 127683 104023 127711 104051
rect 127497 103961 127525 103989
rect 127559 103961 127587 103989
rect 127621 103961 127649 103989
rect 127683 103961 127711 103989
rect 138819 104147 138847 104175
rect 138881 104147 138909 104175
rect 138819 104085 138847 104113
rect 138881 104085 138909 104113
rect 138819 104023 138847 104051
rect 138881 104023 138909 104051
rect 138819 103961 138847 103989
rect 138881 103961 138909 103989
rect 131139 101147 131167 101175
rect 131201 101147 131229 101175
rect 131139 101085 131167 101113
rect 131201 101085 131229 101113
rect 131139 101023 131167 101051
rect 131201 101023 131229 101051
rect 131139 100961 131167 100989
rect 131201 100961 131229 100989
rect 140997 101147 141025 101175
rect 141059 101147 141087 101175
rect 141121 101147 141149 101175
rect 141183 101147 141211 101175
rect 140997 101085 141025 101113
rect 141059 101085 141087 101113
rect 141121 101085 141149 101113
rect 141183 101085 141211 101113
rect 140997 101023 141025 101051
rect 141059 101023 141087 101051
rect 141121 101023 141149 101051
rect 141183 101023 141211 101051
rect 140997 100961 141025 100989
rect 141059 100961 141087 100989
rect 141121 100961 141149 100989
rect 141183 100961 141211 100989
rect 127497 95147 127525 95175
rect 127559 95147 127587 95175
rect 127621 95147 127649 95175
rect 127683 95147 127711 95175
rect 127497 95085 127525 95113
rect 127559 95085 127587 95113
rect 127621 95085 127649 95113
rect 127683 95085 127711 95113
rect 127497 95023 127525 95051
rect 127559 95023 127587 95051
rect 127621 95023 127649 95051
rect 127683 95023 127711 95051
rect 127497 94961 127525 94989
rect 127559 94961 127587 94989
rect 127621 94961 127649 94989
rect 127683 94961 127711 94989
rect 138819 95147 138847 95175
rect 138881 95147 138909 95175
rect 138819 95085 138847 95113
rect 138881 95085 138909 95113
rect 138819 95023 138847 95051
rect 138881 95023 138909 95051
rect 138819 94961 138847 94989
rect 138881 94961 138909 94989
rect 131139 92147 131167 92175
rect 131201 92147 131229 92175
rect 131139 92085 131167 92113
rect 131201 92085 131229 92113
rect 131139 92023 131167 92051
rect 131201 92023 131229 92051
rect 131139 91961 131167 91989
rect 131201 91961 131229 91989
rect 140997 92147 141025 92175
rect 141059 92147 141087 92175
rect 141121 92147 141149 92175
rect 141183 92147 141211 92175
rect 140997 92085 141025 92113
rect 141059 92085 141087 92113
rect 141121 92085 141149 92113
rect 141183 92085 141211 92113
rect 140997 92023 141025 92051
rect 141059 92023 141087 92051
rect 141121 92023 141149 92051
rect 141183 92023 141211 92051
rect 140997 91961 141025 91989
rect 141059 91961 141087 91989
rect 141121 91961 141149 91989
rect 141183 91961 141211 91989
rect 127497 86147 127525 86175
rect 127559 86147 127587 86175
rect 127621 86147 127649 86175
rect 127683 86147 127711 86175
rect 127497 86085 127525 86113
rect 127559 86085 127587 86113
rect 127621 86085 127649 86113
rect 127683 86085 127711 86113
rect 127497 86023 127525 86051
rect 127559 86023 127587 86051
rect 127621 86023 127649 86051
rect 127683 86023 127711 86051
rect 127497 85961 127525 85989
rect 127559 85961 127587 85989
rect 127621 85961 127649 85989
rect 127683 85961 127711 85989
rect 138819 86147 138847 86175
rect 138881 86147 138909 86175
rect 138819 86085 138847 86113
rect 138881 86085 138909 86113
rect 138819 86023 138847 86051
rect 138881 86023 138909 86051
rect 138819 85961 138847 85989
rect 138881 85961 138909 85989
rect 131139 83147 131167 83175
rect 131201 83147 131229 83175
rect 131139 83085 131167 83113
rect 131201 83085 131229 83113
rect 131139 83023 131167 83051
rect 131201 83023 131229 83051
rect 131139 82961 131167 82989
rect 131201 82961 131229 82989
rect 140997 83147 141025 83175
rect 141059 83147 141087 83175
rect 141121 83147 141149 83175
rect 141183 83147 141211 83175
rect 140997 83085 141025 83113
rect 141059 83085 141087 83113
rect 141121 83085 141149 83113
rect 141183 83085 141211 83113
rect 140997 83023 141025 83051
rect 141059 83023 141087 83051
rect 141121 83023 141149 83051
rect 141183 83023 141211 83051
rect 140997 82961 141025 82989
rect 141059 82961 141087 82989
rect 141121 82961 141149 82989
rect 141183 82961 141211 82989
rect 127497 77147 127525 77175
rect 127559 77147 127587 77175
rect 127621 77147 127649 77175
rect 127683 77147 127711 77175
rect 127497 77085 127525 77113
rect 127559 77085 127587 77113
rect 127621 77085 127649 77113
rect 127683 77085 127711 77113
rect 127497 77023 127525 77051
rect 127559 77023 127587 77051
rect 127621 77023 127649 77051
rect 127683 77023 127711 77051
rect 127497 76961 127525 76989
rect 127559 76961 127587 76989
rect 127621 76961 127649 76989
rect 127683 76961 127711 76989
rect 138819 77147 138847 77175
rect 138881 77147 138909 77175
rect 138819 77085 138847 77113
rect 138881 77085 138909 77113
rect 138819 77023 138847 77051
rect 138881 77023 138909 77051
rect 138819 76961 138847 76989
rect 138881 76961 138909 76989
rect 131139 74147 131167 74175
rect 131201 74147 131229 74175
rect 131139 74085 131167 74113
rect 131201 74085 131229 74113
rect 131139 74023 131167 74051
rect 131201 74023 131229 74051
rect 131139 73961 131167 73989
rect 131201 73961 131229 73989
rect 140997 74147 141025 74175
rect 141059 74147 141087 74175
rect 141121 74147 141149 74175
rect 141183 74147 141211 74175
rect 140997 74085 141025 74113
rect 141059 74085 141087 74113
rect 141121 74085 141149 74113
rect 141183 74085 141211 74113
rect 140997 74023 141025 74051
rect 141059 74023 141087 74051
rect 141121 74023 141149 74051
rect 141183 74023 141211 74051
rect 140997 73961 141025 73989
rect 141059 73961 141087 73989
rect 141121 73961 141149 73989
rect 141183 73961 141211 73989
rect 127497 68147 127525 68175
rect 127559 68147 127587 68175
rect 127621 68147 127649 68175
rect 127683 68147 127711 68175
rect 127497 68085 127525 68113
rect 127559 68085 127587 68113
rect 127621 68085 127649 68113
rect 127683 68085 127711 68113
rect 127497 68023 127525 68051
rect 127559 68023 127587 68051
rect 127621 68023 127649 68051
rect 127683 68023 127711 68051
rect 127497 67961 127525 67989
rect 127559 67961 127587 67989
rect 127621 67961 127649 67989
rect 127683 67961 127711 67989
rect 138819 68147 138847 68175
rect 138881 68147 138909 68175
rect 138819 68085 138847 68113
rect 138881 68085 138909 68113
rect 138819 68023 138847 68051
rect 138881 68023 138909 68051
rect 138819 67961 138847 67989
rect 138881 67961 138909 67989
rect 131139 65147 131167 65175
rect 131201 65147 131229 65175
rect 131139 65085 131167 65113
rect 131201 65085 131229 65113
rect 131139 65023 131167 65051
rect 131201 65023 131229 65051
rect 131139 64961 131167 64989
rect 131201 64961 131229 64989
rect 140997 65147 141025 65175
rect 141059 65147 141087 65175
rect 141121 65147 141149 65175
rect 141183 65147 141211 65175
rect 140997 65085 141025 65113
rect 141059 65085 141087 65113
rect 141121 65085 141149 65113
rect 141183 65085 141211 65113
rect 140997 65023 141025 65051
rect 141059 65023 141087 65051
rect 141121 65023 141149 65051
rect 141183 65023 141211 65051
rect 140997 64961 141025 64989
rect 141059 64961 141087 64989
rect 141121 64961 141149 64989
rect 141183 64961 141211 64989
rect 127497 59147 127525 59175
rect 127559 59147 127587 59175
rect 127621 59147 127649 59175
rect 127683 59147 127711 59175
rect 127497 59085 127525 59113
rect 127559 59085 127587 59113
rect 127621 59085 127649 59113
rect 127683 59085 127711 59113
rect 127497 59023 127525 59051
rect 127559 59023 127587 59051
rect 127621 59023 127649 59051
rect 127683 59023 127711 59051
rect 127497 58961 127525 58989
rect 127559 58961 127587 58989
rect 127621 58961 127649 58989
rect 127683 58961 127711 58989
rect 138819 59147 138847 59175
rect 138881 59147 138909 59175
rect 138819 59085 138847 59113
rect 138881 59085 138909 59113
rect 138819 59023 138847 59051
rect 138881 59023 138909 59051
rect 138819 58961 138847 58989
rect 138881 58961 138909 58989
rect 131139 56147 131167 56175
rect 131201 56147 131229 56175
rect 131139 56085 131167 56113
rect 131201 56085 131229 56113
rect 131139 56023 131167 56051
rect 131201 56023 131229 56051
rect 131139 55961 131167 55989
rect 131201 55961 131229 55989
rect 140997 56147 141025 56175
rect 141059 56147 141087 56175
rect 141121 56147 141149 56175
rect 141183 56147 141211 56175
rect 140997 56085 141025 56113
rect 141059 56085 141087 56113
rect 141121 56085 141149 56113
rect 141183 56085 141211 56113
rect 140997 56023 141025 56051
rect 141059 56023 141087 56051
rect 141121 56023 141149 56051
rect 141183 56023 141211 56051
rect 140997 55961 141025 55989
rect 141059 55961 141087 55989
rect 141121 55961 141149 55989
rect 141183 55961 141211 55989
rect 127497 50147 127525 50175
rect 127559 50147 127587 50175
rect 127621 50147 127649 50175
rect 127683 50147 127711 50175
rect 127497 50085 127525 50113
rect 127559 50085 127587 50113
rect 127621 50085 127649 50113
rect 127683 50085 127711 50113
rect 127497 50023 127525 50051
rect 127559 50023 127587 50051
rect 127621 50023 127649 50051
rect 127683 50023 127711 50051
rect 127497 49961 127525 49989
rect 127559 49961 127587 49989
rect 127621 49961 127649 49989
rect 127683 49961 127711 49989
rect 138819 50147 138847 50175
rect 138881 50147 138909 50175
rect 138819 50085 138847 50113
rect 138881 50085 138909 50113
rect 138819 50023 138847 50051
rect 138881 50023 138909 50051
rect 138819 49961 138847 49989
rect 138881 49961 138909 49989
rect 131139 47147 131167 47175
rect 131201 47147 131229 47175
rect 131139 47085 131167 47113
rect 131201 47085 131229 47113
rect 131139 47023 131167 47051
rect 131201 47023 131229 47051
rect 131139 46961 131167 46989
rect 131201 46961 131229 46989
rect 140997 47147 141025 47175
rect 141059 47147 141087 47175
rect 141121 47147 141149 47175
rect 141183 47147 141211 47175
rect 140997 47085 141025 47113
rect 141059 47085 141087 47113
rect 141121 47085 141149 47113
rect 141183 47085 141211 47113
rect 140997 47023 141025 47051
rect 141059 47023 141087 47051
rect 141121 47023 141149 47051
rect 141183 47023 141211 47051
rect 140997 46961 141025 46989
rect 141059 46961 141087 46989
rect 141121 46961 141149 46989
rect 141183 46961 141211 46989
rect 127497 41147 127525 41175
rect 127559 41147 127587 41175
rect 127621 41147 127649 41175
rect 127683 41147 127711 41175
rect 127497 41085 127525 41113
rect 127559 41085 127587 41113
rect 127621 41085 127649 41113
rect 127683 41085 127711 41113
rect 127497 41023 127525 41051
rect 127559 41023 127587 41051
rect 127621 41023 127649 41051
rect 127683 41023 127711 41051
rect 127497 40961 127525 40989
rect 127559 40961 127587 40989
rect 127621 40961 127649 40989
rect 127683 40961 127711 40989
rect 138819 41147 138847 41175
rect 138881 41147 138909 41175
rect 138819 41085 138847 41113
rect 138881 41085 138909 41113
rect 138819 41023 138847 41051
rect 138881 41023 138909 41051
rect 138819 40961 138847 40989
rect 138881 40961 138909 40989
rect 131139 38147 131167 38175
rect 131201 38147 131229 38175
rect 131139 38085 131167 38113
rect 131201 38085 131229 38113
rect 131139 38023 131167 38051
rect 131201 38023 131229 38051
rect 131139 37961 131167 37989
rect 131201 37961 131229 37989
rect 140997 38147 141025 38175
rect 141059 38147 141087 38175
rect 141121 38147 141149 38175
rect 141183 38147 141211 38175
rect 140997 38085 141025 38113
rect 141059 38085 141087 38113
rect 141121 38085 141149 38113
rect 141183 38085 141211 38113
rect 140997 38023 141025 38051
rect 141059 38023 141087 38051
rect 141121 38023 141149 38051
rect 141183 38023 141211 38051
rect 140997 37961 141025 37989
rect 141059 37961 141087 37989
rect 141121 37961 141149 37989
rect 141183 37961 141211 37989
rect 127497 32147 127525 32175
rect 127559 32147 127587 32175
rect 127621 32147 127649 32175
rect 127683 32147 127711 32175
rect 127497 32085 127525 32113
rect 127559 32085 127587 32113
rect 127621 32085 127649 32113
rect 127683 32085 127711 32113
rect 127497 32023 127525 32051
rect 127559 32023 127587 32051
rect 127621 32023 127649 32051
rect 127683 32023 127711 32051
rect 127497 31961 127525 31989
rect 127559 31961 127587 31989
rect 127621 31961 127649 31989
rect 127683 31961 127711 31989
rect 138819 32147 138847 32175
rect 138881 32147 138909 32175
rect 138819 32085 138847 32113
rect 138881 32085 138909 32113
rect 138819 32023 138847 32051
rect 138881 32023 138909 32051
rect 138819 31961 138847 31989
rect 138881 31961 138909 31989
rect 131139 29147 131167 29175
rect 131201 29147 131229 29175
rect 131139 29085 131167 29113
rect 131201 29085 131229 29113
rect 131139 29023 131167 29051
rect 131201 29023 131229 29051
rect 131139 28961 131167 28989
rect 131201 28961 131229 28989
rect 140997 29147 141025 29175
rect 141059 29147 141087 29175
rect 141121 29147 141149 29175
rect 141183 29147 141211 29175
rect 140997 29085 141025 29113
rect 141059 29085 141087 29113
rect 141121 29085 141149 29113
rect 141183 29085 141211 29113
rect 140997 29023 141025 29051
rect 141059 29023 141087 29051
rect 141121 29023 141149 29051
rect 141183 29023 141211 29051
rect 140997 28961 141025 28989
rect 141059 28961 141087 28989
rect 141121 28961 141149 28989
rect 141183 28961 141211 28989
rect 127497 23147 127525 23175
rect 127559 23147 127587 23175
rect 127621 23147 127649 23175
rect 127683 23147 127711 23175
rect 127497 23085 127525 23113
rect 127559 23085 127587 23113
rect 127621 23085 127649 23113
rect 127683 23085 127711 23113
rect 127497 23023 127525 23051
rect 127559 23023 127587 23051
rect 127621 23023 127649 23051
rect 127683 23023 127711 23051
rect 127497 22961 127525 22989
rect 127559 22961 127587 22989
rect 127621 22961 127649 22989
rect 127683 22961 127711 22989
rect 138819 23147 138847 23175
rect 138881 23147 138909 23175
rect 138819 23085 138847 23113
rect 138881 23085 138909 23113
rect 138819 23023 138847 23051
rect 138881 23023 138909 23051
rect 138819 22961 138847 22989
rect 138881 22961 138909 22989
rect 131139 20147 131167 20175
rect 131201 20147 131229 20175
rect 131139 20085 131167 20113
rect 131201 20085 131229 20113
rect 131139 20023 131167 20051
rect 131201 20023 131229 20051
rect 131139 19961 131167 19989
rect 131201 19961 131229 19989
rect 140997 20147 141025 20175
rect 141059 20147 141087 20175
rect 141121 20147 141149 20175
rect 141183 20147 141211 20175
rect 140997 20085 141025 20113
rect 141059 20085 141087 20113
rect 141121 20085 141149 20113
rect 141183 20085 141211 20113
rect 140997 20023 141025 20051
rect 141059 20023 141087 20051
rect 141121 20023 141149 20051
rect 141183 20023 141211 20051
rect 140997 19961 141025 19989
rect 141059 19961 141087 19989
rect 141121 19961 141149 19989
rect 141183 19961 141211 19989
rect 127497 14147 127525 14175
rect 127559 14147 127587 14175
rect 127621 14147 127649 14175
rect 127683 14147 127711 14175
rect 127497 14085 127525 14113
rect 127559 14085 127587 14113
rect 127621 14085 127649 14113
rect 127683 14085 127711 14113
rect 127497 14023 127525 14051
rect 127559 14023 127587 14051
rect 127621 14023 127649 14051
rect 127683 14023 127711 14051
rect 127497 13961 127525 13989
rect 127559 13961 127587 13989
rect 127621 13961 127649 13989
rect 127683 13961 127711 13989
rect 138819 14147 138847 14175
rect 138881 14147 138909 14175
rect 138819 14085 138847 14113
rect 138881 14085 138909 14113
rect 138819 14023 138847 14051
rect 138881 14023 138909 14051
rect 138819 13961 138847 13989
rect 138881 13961 138909 13989
rect 131139 11147 131167 11175
rect 131201 11147 131229 11175
rect 131139 11085 131167 11113
rect 131201 11085 131229 11113
rect 131139 11023 131167 11051
rect 131201 11023 131229 11051
rect 131139 10961 131167 10989
rect 131201 10961 131229 10989
rect 140997 11147 141025 11175
rect 141059 11147 141087 11175
rect 141121 11147 141149 11175
rect 141183 11147 141211 11175
rect 140997 11085 141025 11113
rect 141059 11085 141087 11113
rect 141121 11085 141149 11113
rect 141183 11085 141211 11113
rect 140997 11023 141025 11051
rect 141059 11023 141087 11051
rect 141121 11023 141149 11051
rect 141183 11023 141211 11051
rect 140997 10961 141025 10989
rect 141059 10961 141087 10989
rect 141121 10961 141149 10989
rect 141183 10961 141211 10989
rect 127497 5147 127525 5175
rect 127559 5147 127587 5175
rect 127621 5147 127649 5175
rect 127683 5147 127711 5175
rect 127497 5085 127525 5113
rect 127559 5085 127587 5113
rect 127621 5085 127649 5113
rect 127683 5085 127711 5113
rect 127497 5023 127525 5051
rect 127559 5023 127587 5051
rect 127621 5023 127649 5051
rect 127683 5023 127711 5051
rect 127497 4961 127525 4989
rect 127559 4961 127587 4989
rect 127621 4961 127649 4989
rect 127683 4961 127711 4989
rect 138819 5147 138847 5175
rect 138881 5147 138909 5175
rect 138819 5085 138847 5113
rect 138881 5085 138909 5113
rect 138819 5023 138847 5051
rect 138881 5023 138909 5051
rect 138819 4961 138847 4989
rect 138881 4961 138909 4989
rect 127497 -588 127525 -560
rect 127559 -588 127587 -560
rect 127621 -588 127649 -560
rect 127683 -588 127711 -560
rect 127497 -650 127525 -622
rect 127559 -650 127587 -622
rect 127621 -650 127649 -622
rect 127683 -650 127711 -622
rect 127497 -712 127525 -684
rect 127559 -712 127587 -684
rect 127621 -712 127649 -684
rect 127683 -712 127711 -684
rect 127497 -774 127525 -746
rect 127559 -774 127587 -746
rect 127621 -774 127649 -746
rect 127683 -774 127711 -746
rect 140997 2147 141025 2175
rect 141059 2147 141087 2175
rect 141121 2147 141149 2175
rect 141183 2147 141211 2175
rect 140997 2085 141025 2113
rect 141059 2085 141087 2113
rect 141121 2085 141149 2113
rect 141183 2085 141211 2113
rect 140997 2023 141025 2051
rect 141059 2023 141087 2051
rect 141121 2023 141149 2051
rect 141183 2023 141211 2051
rect 140997 1961 141025 1989
rect 141059 1961 141087 1989
rect 141121 1961 141149 1989
rect 141183 1961 141211 1989
rect 140997 -108 141025 -80
rect 141059 -108 141087 -80
rect 141121 -108 141149 -80
rect 141183 -108 141211 -80
rect 140997 -170 141025 -142
rect 141059 -170 141087 -142
rect 141121 -170 141149 -142
rect 141183 -170 141211 -142
rect 140997 -232 141025 -204
rect 141059 -232 141087 -204
rect 141121 -232 141149 -204
rect 141183 -232 141211 -204
rect 140997 -294 141025 -266
rect 141059 -294 141087 -266
rect 141121 -294 141149 -266
rect 141183 -294 141211 -266
rect 142857 299058 142885 299086
rect 142919 299058 142947 299086
rect 142981 299058 143009 299086
rect 143043 299058 143071 299086
rect 142857 298996 142885 299024
rect 142919 298996 142947 299024
rect 142981 298996 143009 299024
rect 143043 298996 143071 299024
rect 142857 298934 142885 298962
rect 142919 298934 142947 298962
rect 142981 298934 143009 298962
rect 143043 298934 143071 298962
rect 142857 298872 142885 298900
rect 142919 298872 142947 298900
rect 142981 298872 143009 298900
rect 143043 298872 143071 298900
rect 142857 293147 142885 293175
rect 142919 293147 142947 293175
rect 142981 293147 143009 293175
rect 143043 293147 143071 293175
rect 142857 293085 142885 293113
rect 142919 293085 142947 293113
rect 142981 293085 143009 293113
rect 143043 293085 143071 293113
rect 142857 293023 142885 293051
rect 142919 293023 142947 293051
rect 142981 293023 143009 293051
rect 143043 293023 143071 293051
rect 142857 292961 142885 292989
rect 142919 292961 142947 292989
rect 142981 292961 143009 292989
rect 143043 292961 143071 292989
rect 142857 284147 142885 284175
rect 142919 284147 142947 284175
rect 142981 284147 143009 284175
rect 143043 284147 143071 284175
rect 142857 284085 142885 284113
rect 142919 284085 142947 284113
rect 142981 284085 143009 284113
rect 143043 284085 143071 284113
rect 142857 284023 142885 284051
rect 142919 284023 142947 284051
rect 142981 284023 143009 284051
rect 143043 284023 143071 284051
rect 142857 283961 142885 283989
rect 142919 283961 142947 283989
rect 142981 283961 143009 283989
rect 143043 283961 143071 283989
rect 142857 275147 142885 275175
rect 142919 275147 142947 275175
rect 142981 275147 143009 275175
rect 143043 275147 143071 275175
rect 142857 275085 142885 275113
rect 142919 275085 142947 275113
rect 142981 275085 143009 275113
rect 143043 275085 143071 275113
rect 142857 275023 142885 275051
rect 142919 275023 142947 275051
rect 142981 275023 143009 275051
rect 143043 275023 143071 275051
rect 142857 274961 142885 274989
rect 142919 274961 142947 274989
rect 142981 274961 143009 274989
rect 143043 274961 143071 274989
rect 142857 266147 142885 266175
rect 142919 266147 142947 266175
rect 142981 266147 143009 266175
rect 143043 266147 143071 266175
rect 142857 266085 142885 266113
rect 142919 266085 142947 266113
rect 142981 266085 143009 266113
rect 143043 266085 143071 266113
rect 142857 266023 142885 266051
rect 142919 266023 142947 266051
rect 142981 266023 143009 266051
rect 143043 266023 143071 266051
rect 142857 265961 142885 265989
rect 142919 265961 142947 265989
rect 142981 265961 143009 265989
rect 143043 265961 143071 265989
rect 142857 257147 142885 257175
rect 142919 257147 142947 257175
rect 142981 257147 143009 257175
rect 143043 257147 143071 257175
rect 142857 257085 142885 257113
rect 142919 257085 142947 257113
rect 142981 257085 143009 257113
rect 143043 257085 143071 257113
rect 142857 257023 142885 257051
rect 142919 257023 142947 257051
rect 142981 257023 143009 257051
rect 143043 257023 143071 257051
rect 142857 256961 142885 256989
rect 142919 256961 142947 256989
rect 142981 256961 143009 256989
rect 143043 256961 143071 256989
rect 142857 248147 142885 248175
rect 142919 248147 142947 248175
rect 142981 248147 143009 248175
rect 143043 248147 143071 248175
rect 142857 248085 142885 248113
rect 142919 248085 142947 248113
rect 142981 248085 143009 248113
rect 143043 248085 143071 248113
rect 142857 248023 142885 248051
rect 142919 248023 142947 248051
rect 142981 248023 143009 248051
rect 143043 248023 143071 248051
rect 142857 247961 142885 247989
rect 142919 247961 142947 247989
rect 142981 247961 143009 247989
rect 143043 247961 143071 247989
rect 142857 239147 142885 239175
rect 142919 239147 142947 239175
rect 142981 239147 143009 239175
rect 143043 239147 143071 239175
rect 142857 239085 142885 239113
rect 142919 239085 142947 239113
rect 142981 239085 143009 239113
rect 143043 239085 143071 239113
rect 142857 239023 142885 239051
rect 142919 239023 142947 239051
rect 142981 239023 143009 239051
rect 143043 239023 143071 239051
rect 142857 238961 142885 238989
rect 142919 238961 142947 238989
rect 142981 238961 143009 238989
rect 143043 238961 143071 238989
rect 142857 230147 142885 230175
rect 142919 230147 142947 230175
rect 142981 230147 143009 230175
rect 143043 230147 143071 230175
rect 142857 230085 142885 230113
rect 142919 230085 142947 230113
rect 142981 230085 143009 230113
rect 143043 230085 143071 230113
rect 142857 230023 142885 230051
rect 142919 230023 142947 230051
rect 142981 230023 143009 230051
rect 143043 230023 143071 230051
rect 142857 229961 142885 229989
rect 142919 229961 142947 229989
rect 142981 229961 143009 229989
rect 143043 229961 143071 229989
rect 142857 221147 142885 221175
rect 142919 221147 142947 221175
rect 142981 221147 143009 221175
rect 143043 221147 143071 221175
rect 142857 221085 142885 221113
rect 142919 221085 142947 221113
rect 142981 221085 143009 221113
rect 143043 221085 143071 221113
rect 142857 221023 142885 221051
rect 142919 221023 142947 221051
rect 142981 221023 143009 221051
rect 143043 221023 143071 221051
rect 142857 220961 142885 220989
rect 142919 220961 142947 220989
rect 142981 220961 143009 220989
rect 143043 220961 143071 220989
rect 142857 212147 142885 212175
rect 142919 212147 142947 212175
rect 142981 212147 143009 212175
rect 143043 212147 143071 212175
rect 142857 212085 142885 212113
rect 142919 212085 142947 212113
rect 142981 212085 143009 212113
rect 143043 212085 143071 212113
rect 142857 212023 142885 212051
rect 142919 212023 142947 212051
rect 142981 212023 143009 212051
rect 143043 212023 143071 212051
rect 142857 211961 142885 211989
rect 142919 211961 142947 211989
rect 142981 211961 143009 211989
rect 143043 211961 143071 211989
rect 142857 203147 142885 203175
rect 142919 203147 142947 203175
rect 142981 203147 143009 203175
rect 143043 203147 143071 203175
rect 142857 203085 142885 203113
rect 142919 203085 142947 203113
rect 142981 203085 143009 203113
rect 143043 203085 143071 203113
rect 142857 203023 142885 203051
rect 142919 203023 142947 203051
rect 142981 203023 143009 203051
rect 143043 203023 143071 203051
rect 142857 202961 142885 202989
rect 142919 202961 142947 202989
rect 142981 202961 143009 202989
rect 143043 202961 143071 202989
rect 142857 194147 142885 194175
rect 142919 194147 142947 194175
rect 142981 194147 143009 194175
rect 143043 194147 143071 194175
rect 142857 194085 142885 194113
rect 142919 194085 142947 194113
rect 142981 194085 143009 194113
rect 143043 194085 143071 194113
rect 142857 194023 142885 194051
rect 142919 194023 142947 194051
rect 142981 194023 143009 194051
rect 143043 194023 143071 194051
rect 142857 193961 142885 193989
rect 142919 193961 142947 193989
rect 142981 193961 143009 193989
rect 143043 193961 143071 193989
rect 142857 185147 142885 185175
rect 142919 185147 142947 185175
rect 142981 185147 143009 185175
rect 143043 185147 143071 185175
rect 142857 185085 142885 185113
rect 142919 185085 142947 185113
rect 142981 185085 143009 185113
rect 143043 185085 143071 185113
rect 142857 185023 142885 185051
rect 142919 185023 142947 185051
rect 142981 185023 143009 185051
rect 143043 185023 143071 185051
rect 142857 184961 142885 184989
rect 142919 184961 142947 184989
rect 142981 184961 143009 184989
rect 143043 184961 143071 184989
rect 142857 176147 142885 176175
rect 142919 176147 142947 176175
rect 142981 176147 143009 176175
rect 143043 176147 143071 176175
rect 142857 176085 142885 176113
rect 142919 176085 142947 176113
rect 142981 176085 143009 176113
rect 143043 176085 143071 176113
rect 142857 176023 142885 176051
rect 142919 176023 142947 176051
rect 142981 176023 143009 176051
rect 143043 176023 143071 176051
rect 142857 175961 142885 175989
rect 142919 175961 142947 175989
rect 142981 175961 143009 175989
rect 143043 175961 143071 175989
rect 156357 298578 156385 298606
rect 156419 298578 156447 298606
rect 156481 298578 156509 298606
rect 156543 298578 156571 298606
rect 156357 298516 156385 298544
rect 156419 298516 156447 298544
rect 156481 298516 156509 298544
rect 156543 298516 156571 298544
rect 156357 298454 156385 298482
rect 156419 298454 156447 298482
rect 156481 298454 156509 298482
rect 156543 298454 156571 298482
rect 156357 298392 156385 298420
rect 156419 298392 156447 298420
rect 156481 298392 156509 298420
rect 156543 298392 156571 298420
rect 156357 290147 156385 290175
rect 156419 290147 156447 290175
rect 156481 290147 156509 290175
rect 156543 290147 156571 290175
rect 156357 290085 156385 290113
rect 156419 290085 156447 290113
rect 156481 290085 156509 290113
rect 156543 290085 156571 290113
rect 156357 290023 156385 290051
rect 156419 290023 156447 290051
rect 156481 290023 156509 290051
rect 156543 290023 156571 290051
rect 156357 289961 156385 289989
rect 156419 289961 156447 289989
rect 156481 289961 156509 289989
rect 156543 289961 156571 289989
rect 156357 281147 156385 281175
rect 156419 281147 156447 281175
rect 156481 281147 156509 281175
rect 156543 281147 156571 281175
rect 156357 281085 156385 281113
rect 156419 281085 156447 281113
rect 156481 281085 156509 281113
rect 156543 281085 156571 281113
rect 156357 281023 156385 281051
rect 156419 281023 156447 281051
rect 156481 281023 156509 281051
rect 156543 281023 156571 281051
rect 156357 280961 156385 280989
rect 156419 280961 156447 280989
rect 156481 280961 156509 280989
rect 156543 280961 156571 280989
rect 156357 272147 156385 272175
rect 156419 272147 156447 272175
rect 156481 272147 156509 272175
rect 156543 272147 156571 272175
rect 156357 272085 156385 272113
rect 156419 272085 156447 272113
rect 156481 272085 156509 272113
rect 156543 272085 156571 272113
rect 156357 272023 156385 272051
rect 156419 272023 156447 272051
rect 156481 272023 156509 272051
rect 156543 272023 156571 272051
rect 156357 271961 156385 271989
rect 156419 271961 156447 271989
rect 156481 271961 156509 271989
rect 156543 271961 156571 271989
rect 156357 263147 156385 263175
rect 156419 263147 156447 263175
rect 156481 263147 156509 263175
rect 156543 263147 156571 263175
rect 156357 263085 156385 263113
rect 156419 263085 156447 263113
rect 156481 263085 156509 263113
rect 156543 263085 156571 263113
rect 156357 263023 156385 263051
rect 156419 263023 156447 263051
rect 156481 263023 156509 263051
rect 156543 263023 156571 263051
rect 156357 262961 156385 262989
rect 156419 262961 156447 262989
rect 156481 262961 156509 262989
rect 156543 262961 156571 262989
rect 156357 254147 156385 254175
rect 156419 254147 156447 254175
rect 156481 254147 156509 254175
rect 156543 254147 156571 254175
rect 156357 254085 156385 254113
rect 156419 254085 156447 254113
rect 156481 254085 156509 254113
rect 156543 254085 156571 254113
rect 156357 254023 156385 254051
rect 156419 254023 156447 254051
rect 156481 254023 156509 254051
rect 156543 254023 156571 254051
rect 156357 253961 156385 253989
rect 156419 253961 156447 253989
rect 156481 253961 156509 253989
rect 156543 253961 156571 253989
rect 156357 245147 156385 245175
rect 156419 245147 156447 245175
rect 156481 245147 156509 245175
rect 156543 245147 156571 245175
rect 156357 245085 156385 245113
rect 156419 245085 156447 245113
rect 156481 245085 156509 245113
rect 156543 245085 156571 245113
rect 156357 245023 156385 245051
rect 156419 245023 156447 245051
rect 156481 245023 156509 245051
rect 156543 245023 156571 245051
rect 156357 244961 156385 244989
rect 156419 244961 156447 244989
rect 156481 244961 156509 244989
rect 156543 244961 156571 244989
rect 156357 236147 156385 236175
rect 156419 236147 156447 236175
rect 156481 236147 156509 236175
rect 156543 236147 156571 236175
rect 156357 236085 156385 236113
rect 156419 236085 156447 236113
rect 156481 236085 156509 236113
rect 156543 236085 156571 236113
rect 156357 236023 156385 236051
rect 156419 236023 156447 236051
rect 156481 236023 156509 236051
rect 156543 236023 156571 236051
rect 156357 235961 156385 235989
rect 156419 235961 156447 235989
rect 156481 235961 156509 235989
rect 156543 235961 156571 235989
rect 156357 227147 156385 227175
rect 156419 227147 156447 227175
rect 156481 227147 156509 227175
rect 156543 227147 156571 227175
rect 156357 227085 156385 227113
rect 156419 227085 156447 227113
rect 156481 227085 156509 227113
rect 156543 227085 156571 227113
rect 156357 227023 156385 227051
rect 156419 227023 156447 227051
rect 156481 227023 156509 227051
rect 156543 227023 156571 227051
rect 156357 226961 156385 226989
rect 156419 226961 156447 226989
rect 156481 226961 156509 226989
rect 156543 226961 156571 226989
rect 156357 218147 156385 218175
rect 156419 218147 156447 218175
rect 156481 218147 156509 218175
rect 156543 218147 156571 218175
rect 156357 218085 156385 218113
rect 156419 218085 156447 218113
rect 156481 218085 156509 218113
rect 156543 218085 156571 218113
rect 156357 218023 156385 218051
rect 156419 218023 156447 218051
rect 156481 218023 156509 218051
rect 156543 218023 156571 218051
rect 156357 217961 156385 217989
rect 156419 217961 156447 217989
rect 156481 217961 156509 217989
rect 156543 217961 156571 217989
rect 156357 209147 156385 209175
rect 156419 209147 156447 209175
rect 156481 209147 156509 209175
rect 156543 209147 156571 209175
rect 156357 209085 156385 209113
rect 156419 209085 156447 209113
rect 156481 209085 156509 209113
rect 156543 209085 156571 209113
rect 156357 209023 156385 209051
rect 156419 209023 156447 209051
rect 156481 209023 156509 209051
rect 156543 209023 156571 209051
rect 156357 208961 156385 208989
rect 156419 208961 156447 208989
rect 156481 208961 156509 208989
rect 156543 208961 156571 208989
rect 156357 200147 156385 200175
rect 156419 200147 156447 200175
rect 156481 200147 156509 200175
rect 156543 200147 156571 200175
rect 156357 200085 156385 200113
rect 156419 200085 156447 200113
rect 156481 200085 156509 200113
rect 156543 200085 156571 200113
rect 156357 200023 156385 200051
rect 156419 200023 156447 200051
rect 156481 200023 156509 200051
rect 156543 200023 156571 200051
rect 156357 199961 156385 199989
rect 156419 199961 156447 199989
rect 156481 199961 156509 199989
rect 156543 199961 156571 199989
rect 156357 191147 156385 191175
rect 156419 191147 156447 191175
rect 156481 191147 156509 191175
rect 156543 191147 156571 191175
rect 156357 191085 156385 191113
rect 156419 191085 156447 191113
rect 156481 191085 156509 191113
rect 156543 191085 156571 191113
rect 156357 191023 156385 191051
rect 156419 191023 156447 191051
rect 156481 191023 156509 191051
rect 156543 191023 156571 191051
rect 156357 190961 156385 190989
rect 156419 190961 156447 190989
rect 156481 190961 156509 190989
rect 156543 190961 156571 190989
rect 156357 182147 156385 182175
rect 156419 182147 156447 182175
rect 156481 182147 156509 182175
rect 156543 182147 156571 182175
rect 156357 182085 156385 182113
rect 156419 182085 156447 182113
rect 156481 182085 156509 182113
rect 156543 182085 156571 182113
rect 156357 182023 156385 182051
rect 156419 182023 156447 182051
rect 156481 182023 156509 182051
rect 156543 182023 156571 182051
rect 156357 181961 156385 181989
rect 156419 181961 156447 181989
rect 156481 181961 156509 181989
rect 156543 181961 156571 181989
rect 146499 173147 146527 173175
rect 146561 173147 146589 173175
rect 146499 173085 146527 173113
rect 146561 173085 146589 173113
rect 146499 173023 146527 173051
rect 146561 173023 146589 173051
rect 146499 172961 146527 172989
rect 146561 172961 146589 172989
rect 156357 173147 156385 173175
rect 156419 173147 156447 173175
rect 156481 173147 156509 173175
rect 156543 173147 156571 173175
rect 156357 173085 156385 173113
rect 156419 173085 156447 173113
rect 156481 173085 156509 173113
rect 156543 173085 156571 173113
rect 156357 173023 156385 173051
rect 156419 173023 156447 173051
rect 156481 173023 156509 173051
rect 156543 173023 156571 173051
rect 156357 172961 156385 172989
rect 156419 172961 156447 172989
rect 156481 172961 156509 172989
rect 156543 172961 156571 172989
rect 142857 167147 142885 167175
rect 142919 167147 142947 167175
rect 142981 167147 143009 167175
rect 143043 167147 143071 167175
rect 142857 167085 142885 167113
rect 142919 167085 142947 167113
rect 142981 167085 143009 167113
rect 143043 167085 143071 167113
rect 142857 167023 142885 167051
rect 142919 167023 142947 167051
rect 142981 167023 143009 167051
rect 143043 167023 143071 167051
rect 142857 166961 142885 166989
rect 142919 166961 142947 166989
rect 142981 166961 143009 166989
rect 143043 166961 143071 166989
rect 154179 167147 154207 167175
rect 154241 167147 154269 167175
rect 154179 167085 154207 167113
rect 154241 167085 154269 167113
rect 154179 167023 154207 167051
rect 154241 167023 154269 167051
rect 154179 166961 154207 166989
rect 154241 166961 154269 166989
rect 146499 164147 146527 164175
rect 146561 164147 146589 164175
rect 146499 164085 146527 164113
rect 146561 164085 146589 164113
rect 146499 164023 146527 164051
rect 146561 164023 146589 164051
rect 146499 163961 146527 163989
rect 146561 163961 146589 163989
rect 156357 164147 156385 164175
rect 156419 164147 156447 164175
rect 156481 164147 156509 164175
rect 156543 164147 156571 164175
rect 156357 164085 156385 164113
rect 156419 164085 156447 164113
rect 156481 164085 156509 164113
rect 156543 164085 156571 164113
rect 156357 164023 156385 164051
rect 156419 164023 156447 164051
rect 156481 164023 156509 164051
rect 156543 164023 156571 164051
rect 156357 163961 156385 163989
rect 156419 163961 156447 163989
rect 156481 163961 156509 163989
rect 156543 163961 156571 163989
rect 142857 158147 142885 158175
rect 142919 158147 142947 158175
rect 142981 158147 143009 158175
rect 143043 158147 143071 158175
rect 142857 158085 142885 158113
rect 142919 158085 142947 158113
rect 142981 158085 143009 158113
rect 143043 158085 143071 158113
rect 142857 158023 142885 158051
rect 142919 158023 142947 158051
rect 142981 158023 143009 158051
rect 143043 158023 143071 158051
rect 142857 157961 142885 157989
rect 142919 157961 142947 157989
rect 142981 157961 143009 157989
rect 143043 157961 143071 157989
rect 154179 158147 154207 158175
rect 154241 158147 154269 158175
rect 154179 158085 154207 158113
rect 154241 158085 154269 158113
rect 154179 158023 154207 158051
rect 154241 158023 154269 158051
rect 154179 157961 154207 157989
rect 154241 157961 154269 157989
rect 146499 155147 146527 155175
rect 146561 155147 146589 155175
rect 146499 155085 146527 155113
rect 146561 155085 146589 155113
rect 146499 155023 146527 155051
rect 146561 155023 146589 155051
rect 146499 154961 146527 154989
rect 146561 154961 146589 154989
rect 156357 155147 156385 155175
rect 156419 155147 156447 155175
rect 156481 155147 156509 155175
rect 156543 155147 156571 155175
rect 156357 155085 156385 155113
rect 156419 155085 156447 155113
rect 156481 155085 156509 155113
rect 156543 155085 156571 155113
rect 156357 155023 156385 155051
rect 156419 155023 156447 155051
rect 156481 155023 156509 155051
rect 156543 155023 156571 155051
rect 156357 154961 156385 154989
rect 156419 154961 156447 154989
rect 156481 154961 156509 154989
rect 156543 154961 156571 154989
rect 142857 149147 142885 149175
rect 142919 149147 142947 149175
rect 142981 149147 143009 149175
rect 143043 149147 143071 149175
rect 142857 149085 142885 149113
rect 142919 149085 142947 149113
rect 142981 149085 143009 149113
rect 143043 149085 143071 149113
rect 142857 149023 142885 149051
rect 142919 149023 142947 149051
rect 142981 149023 143009 149051
rect 143043 149023 143071 149051
rect 142857 148961 142885 148989
rect 142919 148961 142947 148989
rect 142981 148961 143009 148989
rect 143043 148961 143071 148989
rect 154179 149147 154207 149175
rect 154241 149147 154269 149175
rect 154179 149085 154207 149113
rect 154241 149085 154269 149113
rect 154179 149023 154207 149051
rect 154241 149023 154269 149051
rect 154179 148961 154207 148989
rect 154241 148961 154269 148989
rect 146499 146147 146527 146175
rect 146561 146147 146589 146175
rect 146499 146085 146527 146113
rect 146561 146085 146589 146113
rect 146499 146023 146527 146051
rect 146561 146023 146589 146051
rect 146499 145961 146527 145989
rect 146561 145961 146589 145989
rect 156357 146147 156385 146175
rect 156419 146147 156447 146175
rect 156481 146147 156509 146175
rect 156543 146147 156571 146175
rect 156357 146085 156385 146113
rect 156419 146085 156447 146113
rect 156481 146085 156509 146113
rect 156543 146085 156571 146113
rect 156357 146023 156385 146051
rect 156419 146023 156447 146051
rect 156481 146023 156509 146051
rect 156543 146023 156571 146051
rect 156357 145961 156385 145989
rect 156419 145961 156447 145989
rect 156481 145961 156509 145989
rect 156543 145961 156571 145989
rect 142857 140147 142885 140175
rect 142919 140147 142947 140175
rect 142981 140147 143009 140175
rect 143043 140147 143071 140175
rect 142857 140085 142885 140113
rect 142919 140085 142947 140113
rect 142981 140085 143009 140113
rect 143043 140085 143071 140113
rect 142857 140023 142885 140051
rect 142919 140023 142947 140051
rect 142981 140023 143009 140051
rect 143043 140023 143071 140051
rect 142857 139961 142885 139989
rect 142919 139961 142947 139989
rect 142981 139961 143009 139989
rect 143043 139961 143071 139989
rect 154179 140147 154207 140175
rect 154241 140147 154269 140175
rect 154179 140085 154207 140113
rect 154241 140085 154269 140113
rect 154179 140023 154207 140051
rect 154241 140023 154269 140051
rect 154179 139961 154207 139989
rect 154241 139961 154269 139989
rect 146499 137147 146527 137175
rect 146561 137147 146589 137175
rect 146499 137085 146527 137113
rect 146561 137085 146589 137113
rect 146499 137023 146527 137051
rect 146561 137023 146589 137051
rect 146499 136961 146527 136989
rect 146561 136961 146589 136989
rect 156357 137147 156385 137175
rect 156419 137147 156447 137175
rect 156481 137147 156509 137175
rect 156543 137147 156571 137175
rect 156357 137085 156385 137113
rect 156419 137085 156447 137113
rect 156481 137085 156509 137113
rect 156543 137085 156571 137113
rect 156357 137023 156385 137051
rect 156419 137023 156447 137051
rect 156481 137023 156509 137051
rect 156543 137023 156571 137051
rect 156357 136961 156385 136989
rect 156419 136961 156447 136989
rect 156481 136961 156509 136989
rect 156543 136961 156571 136989
rect 142857 131147 142885 131175
rect 142919 131147 142947 131175
rect 142981 131147 143009 131175
rect 143043 131147 143071 131175
rect 142857 131085 142885 131113
rect 142919 131085 142947 131113
rect 142981 131085 143009 131113
rect 143043 131085 143071 131113
rect 142857 131023 142885 131051
rect 142919 131023 142947 131051
rect 142981 131023 143009 131051
rect 143043 131023 143071 131051
rect 142857 130961 142885 130989
rect 142919 130961 142947 130989
rect 142981 130961 143009 130989
rect 143043 130961 143071 130989
rect 154179 131147 154207 131175
rect 154241 131147 154269 131175
rect 154179 131085 154207 131113
rect 154241 131085 154269 131113
rect 154179 131023 154207 131051
rect 154241 131023 154269 131051
rect 154179 130961 154207 130989
rect 154241 130961 154269 130989
rect 146499 128147 146527 128175
rect 146561 128147 146589 128175
rect 146499 128085 146527 128113
rect 146561 128085 146589 128113
rect 146499 128023 146527 128051
rect 146561 128023 146589 128051
rect 146499 127961 146527 127989
rect 146561 127961 146589 127989
rect 156357 128147 156385 128175
rect 156419 128147 156447 128175
rect 156481 128147 156509 128175
rect 156543 128147 156571 128175
rect 156357 128085 156385 128113
rect 156419 128085 156447 128113
rect 156481 128085 156509 128113
rect 156543 128085 156571 128113
rect 156357 128023 156385 128051
rect 156419 128023 156447 128051
rect 156481 128023 156509 128051
rect 156543 128023 156571 128051
rect 156357 127961 156385 127989
rect 156419 127961 156447 127989
rect 156481 127961 156509 127989
rect 156543 127961 156571 127989
rect 142857 122147 142885 122175
rect 142919 122147 142947 122175
rect 142981 122147 143009 122175
rect 143043 122147 143071 122175
rect 142857 122085 142885 122113
rect 142919 122085 142947 122113
rect 142981 122085 143009 122113
rect 143043 122085 143071 122113
rect 142857 122023 142885 122051
rect 142919 122023 142947 122051
rect 142981 122023 143009 122051
rect 143043 122023 143071 122051
rect 142857 121961 142885 121989
rect 142919 121961 142947 121989
rect 142981 121961 143009 121989
rect 143043 121961 143071 121989
rect 154179 122147 154207 122175
rect 154241 122147 154269 122175
rect 154179 122085 154207 122113
rect 154241 122085 154269 122113
rect 154179 122023 154207 122051
rect 154241 122023 154269 122051
rect 154179 121961 154207 121989
rect 154241 121961 154269 121989
rect 146499 119147 146527 119175
rect 146561 119147 146589 119175
rect 146499 119085 146527 119113
rect 146561 119085 146589 119113
rect 146499 119023 146527 119051
rect 146561 119023 146589 119051
rect 146499 118961 146527 118989
rect 146561 118961 146589 118989
rect 156357 119147 156385 119175
rect 156419 119147 156447 119175
rect 156481 119147 156509 119175
rect 156543 119147 156571 119175
rect 156357 119085 156385 119113
rect 156419 119085 156447 119113
rect 156481 119085 156509 119113
rect 156543 119085 156571 119113
rect 156357 119023 156385 119051
rect 156419 119023 156447 119051
rect 156481 119023 156509 119051
rect 156543 119023 156571 119051
rect 156357 118961 156385 118989
rect 156419 118961 156447 118989
rect 156481 118961 156509 118989
rect 156543 118961 156571 118989
rect 142857 113147 142885 113175
rect 142919 113147 142947 113175
rect 142981 113147 143009 113175
rect 143043 113147 143071 113175
rect 142857 113085 142885 113113
rect 142919 113085 142947 113113
rect 142981 113085 143009 113113
rect 143043 113085 143071 113113
rect 142857 113023 142885 113051
rect 142919 113023 142947 113051
rect 142981 113023 143009 113051
rect 143043 113023 143071 113051
rect 142857 112961 142885 112989
rect 142919 112961 142947 112989
rect 142981 112961 143009 112989
rect 143043 112961 143071 112989
rect 154179 113147 154207 113175
rect 154241 113147 154269 113175
rect 154179 113085 154207 113113
rect 154241 113085 154269 113113
rect 154179 113023 154207 113051
rect 154241 113023 154269 113051
rect 154179 112961 154207 112989
rect 154241 112961 154269 112989
rect 146499 110147 146527 110175
rect 146561 110147 146589 110175
rect 146499 110085 146527 110113
rect 146561 110085 146589 110113
rect 146499 110023 146527 110051
rect 146561 110023 146589 110051
rect 146499 109961 146527 109989
rect 146561 109961 146589 109989
rect 156357 110147 156385 110175
rect 156419 110147 156447 110175
rect 156481 110147 156509 110175
rect 156543 110147 156571 110175
rect 156357 110085 156385 110113
rect 156419 110085 156447 110113
rect 156481 110085 156509 110113
rect 156543 110085 156571 110113
rect 156357 110023 156385 110051
rect 156419 110023 156447 110051
rect 156481 110023 156509 110051
rect 156543 110023 156571 110051
rect 156357 109961 156385 109989
rect 156419 109961 156447 109989
rect 156481 109961 156509 109989
rect 156543 109961 156571 109989
rect 142857 104147 142885 104175
rect 142919 104147 142947 104175
rect 142981 104147 143009 104175
rect 143043 104147 143071 104175
rect 142857 104085 142885 104113
rect 142919 104085 142947 104113
rect 142981 104085 143009 104113
rect 143043 104085 143071 104113
rect 142857 104023 142885 104051
rect 142919 104023 142947 104051
rect 142981 104023 143009 104051
rect 143043 104023 143071 104051
rect 142857 103961 142885 103989
rect 142919 103961 142947 103989
rect 142981 103961 143009 103989
rect 143043 103961 143071 103989
rect 154179 104147 154207 104175
rect 154241 104147 154269 104175
rect 154179 104085 154207 104113
rect 154241 104085 154269 104113
rect 154179 104023 154207 104051
rect 154241 104023 154269 104051
rect 154179 103961 154207 103989
rect 154241 103961 154269 103989
rect 146499 101147 146527 101175
rect 146561 101147 146589 101175
rect 146499 101085 146527 101113
rect 146561 101085 146589 101113
rect 146499 101023 146527 101051
rect 146561 101023 146589 101051
rect 146499 100961 146527 100989
rect 146561 100961 146589 100989
rect 156357 101147 156385 101175
rect 156419 101147 156447 101175
rect 156481 101147 156509 101175
rect 156543 101147 156571 101175
rect 156357 101085 156385 101113
rect 156419 101085 156447 101113
rect 156481 101085 156509 101113
rect 156543 101085 156571 101113
rect 156357 101023 156385 101051
rect 156419 101023 156447 101051
rect 156481 101023 156509 101051
rect 156543 101023 156571 101051
rect 156357 100961 156385 100989
rect 156419 100961 156447 100989
rect 156481 100961 156509 100989
rect 156543 100961 156571 100989
rect 142857 95147 142885 95175
rect 142919 95147 142947 95175
rect 142981 95147 143009 95175
rect 143043 95147 143071 95175
rect 142857 95085 142885 95113
rect 142919 95085 142947 95113
rect 142981 95085 143009 95113
rect 143043 95085 143071 95113
rect 142857 95023 142885 95051
rect 142919 95023 142947 95051
rect 142981 95023 143009 95051
rect 143043 95023 143071 95051
rect 142857 94961 142885 94989
rect 142919 94961 142947 94989
rect 142981 94961 143009 94989
rect 143043 94961 143071 94989
rect 154179 95147 154207 95175
rect 154241 95147 154269 95175
rect 154179 95085 154207 95113
rect 154241 95085 154269 95113
rect 154179 95023 154207 95051
rect 154241 95023 154269 95051
rect 154179 94961 154207 94989
rect 154241 94961 154269 94989
rect 146499 92147 146527 92175
rect 146561 92147 146589 92175
rect 146499 92085 146527 92113
rect 146561 92085 146589 92113
rect 146499 92023 146527 92051
rect 146561 92023 146589 92051
rect 146499 91961 146527 91989
rect 146561 91961 146589 91989
rect 156357 92147 156385 92175
rect 156419 92147 156447 92175
rect 156481 92147 156509 92175
rect 156543 92147 156571 92175
rect 156357 92085 156385 92113
rect 156419 92085 156447 92113
rect 156481 92085 156509 92113
rect 156543 92085 156571 92113
rect 156357 92023 156385 92051
rect 156419 92023 156447 92051
rect 156481 92023 156509 92051
rect 156543 92023 156571 92051
rect 156357 91961 156385 91989
rect 156419 91961 156447 91989
rect 156481 91961 156509 91989
rect 156543 91961 156571 91989
rect 142857 86147 142885 86175
rect 142919 86147 142947 86175
rect 142981 86147 143009 86175
rect 143043 86147 143071 86175
rect 142857 86085 142885 86113
rect 142919 86085 142947 86113
rect 142981 86085 143009 86113
rect 143043 86085 143071 86113
rect 142857 86023 142885 86051
rect 142919 86023 142947 86051
rect 142981 86023 143009 86051
rect 143043 86023 143071 86051
rect 142857 85961 142885 85989
rect 142919 85961 142947 85989
rect 142981 85961 143009 85989
rect 143043 85961 143071 85989
rect 154179 86147 154207 86175
rect 154241 86147 154269 86175
rect 154179 86085 154207 86113
rect 154241 86085 154269 86113
rect 154179 86023 154207 86051
rect 154241 86023 154269 86051
rect 154179 85961 154207 85989
rect 154241 85961 154269 85989
rect 146499 83147 146527 83175
rect 146561 83147 146589 83175
rect 146499 83085 146527 83113
rect 146561 83085 146589 83113
rect 146499 83023 146527 83051
rect 146561 83023 146589 83051
rect 146499 82961 146527 82989
rect 146561 82961 146589 82989
rect 156357 83147 156385 83175
rect 156419 83147 156447 83175
rect 156481 83147 156509 83175
rect 156543 83147 156571 83175
rect 156357 83085 156385 83113
rect 156419 83085 156447 83113
rect 156481 83085 156509 83113
rect 156543 83085 156571 83113
rect 156357 83023 156385 83051
rect 156419 83023 156447 83051
rect 156481 83023 156509 83051
rect 156543 83023 156571 83051
rect 156357 82961 156385 82989
rect 156419 82961 156447 82989
rect 156481 82961 156509 82989
rect 156543 82961 156571 82989
rect 142857 77147 142885 77175
rect 142919 77147 142947 77175
rect 142981 77147 143009 77175
rect 143043 77147 143071 77175
rect 142857 77085 142885 77113
rect 142919 77085 142947 77113
rect 142981 77085 143009 77113
rect 143043 77085 143071 77113
rect 142857 77023 142885 77051
rect 142919 77023 142947 77051
rect 142981 77023 143009 77051
rect 143043 77023 143071 77051
rect 142857 76961 142885 76989
rect 142919 76961 142947 76989
rect 142981 76961 143009 76989
rect 143043 76961 143071 76989
rect 154179 77147 154207 77175
rect 154241 77147 154269 77175
rect 154179 77085 154207 77113
rect 154241 77085 154269 77113
rect 154179 77023 154207 77051
rect 154241 77023 154269 77051
rect 154179 76961 154207 76989
rect 154241 76961 154269 76989
rect 146499 74147 146527 74175
rect 146561 74147 146589 74175
rect 146499 74085 146527 74113
rect 146561 74085 146589 74113
rect 146499 74023 146527 74051
rect 146561 74023 146589 74051
rect 146499 73961 146527 73989
rect 146561 73961 146589 73989
rect 156357 74147 156385 74175
rect 156419 74147 156447 74175
rect 156481 74147 156509 74175
rect 156543 74147 156571 74175
rect 156357 74085 156385 74113
rect 156419 74085 156447 74113
rect 156481 74085 156509 74113
rect 156543 74085 156571 74113
rect 156357 74023 156385 74051
rect 156419 74023 156447 74051
rect 156481 74023 156509 74051
rect 156543 74023 156571 74051
rect 156357 73961 156385 73989
rect 156419 73961 156447 73989
rect 156481 73961 156509 73989
rect 156543 73961 156571 73989
rect 142857 68147 142885 68175
rect 142919 68147 142947 68175
rect 142981 68147 143009 68175
rect 143043 68147 143071 68175
rect 142857 68085 142885 68113
rect 142919 68085 142947 68113
rect 142981 68085 143009 68113
rect 143043 68085 143071 68113
rect 142857 68023 142885 68051
rect 142919 68023 142947 68051
rect 142981 68023 143009 68051
rect 143043 68023 143071 68051
rect 142857 67961 142885 67989
rect 142919 67961 142947 67989
rect 142981 67961 143009 67989
rect 143043 67961 143071 67989
rect 154179 68147 154207 68175
rect 154241 68147 154269 68175
rect 154179 68085 154207 68113
rect 154241 68085 154269 68113
rect 154179 68023 154207 68051
rect 154241 68023 154269 68051
rect 154179 67961 154207 67989
rect 154241 67961 154269 67989
rect 146499 65147 146527 65175
rect 146561 65147 146589 65175
rect 146499 65085 146527 65113
rect 146561 65085 146589 65113
rect 146499 65023 146527 65051
rect 146561 65023 146589 65051
rect 146499 64961 146527 64989
rect 146561 64961 146589 64989
rect 156357 65147 156385 65175
rect 156419 65147 156447 65175
rect 156481 65147 156509 65175
rect 156543 65147 156571 65175
rect 156357 65085 156385 65113
rect 156419 65085 156447 65113
rect 156481 65085 156509 65113
rect 156543 65085 156571 65113
rect 156357 65023 156385 65051
rect 156419 65023 156447 65051
rect 156481 65023 156509 65051
rect 156543 65023 156571 65051
rect 156357 64961 156385 64989
rect 156419 64961 156447 64989
rect 156481 64961 156509 64989
rect 156543 64961 156571 64989
rect 142857 59147 142885 59175
rect 142919 59147 142947 59175
rect 142981 59147 143009 59175
rect 143043 59147 143071 59175
rect 142857 59085 142885 59113
rect 142919 59085 142947 59113
rect 142981 59085 143009 59113
rect 143043 59085 143071 59113
rect 142857 59023 142885 59051
rect 142919 59023 142947 59051
rect 142981 59023 143009 59051
rect 143043 59023 143071 59051
rect 142857 58961 142885 58989
rect 142919 58961 142947 58989
rect 142981 58961 143009 58989
rect 143043 58961 143071 58989
rect 154179 59147 154207 59175
rect 154241 59147 154269 59175
rect 154179 59085 154207 59113
rect 154241 59085 154269 59113
rect 154179 59023 154207 59051
rect 154241 59023 154269 59051
rect 154179 58961 154207 58989
rect 154241 58961 154269 58989
rect 146499 56147 146527 56175
rect 146561 56147 146589 56175
rect 146499 56085 146527 56113
rect 146561 56085 146589 56113
rect 146499 56023 146527 56051
rect 146561 56023 146589 56051
rect 146499 55961 146527 55989
rect 146561 55961 146589 55989
rect 156357 56147 156385 56175
rect 156419 56147 156447 56175
rect 156481 56147 156509 56175
rect 156543 56147 156571 56175
rect 156357 56085 156385 56113
rect 156419 56085 156447 56113
rect 156481 56085 156509 56113
rect 156543 56085 156571 56113
rect 156357 56023 156385 56051
rect 156419 56023 156447 56051
rect 156481 56023 156509 56051
rect 156543 56023 156571 56051
rect 156357 55961 156385 55989
rect 156419 55961 156447 55989
rect 156481 55961 156509 55989
rect 156543 55961 156571 55989
rect 142857 50147 142885 50175
rect 142919 50147 142947 50175
rect 142981 50147 143009 50175
rect 143043 50147 143071 50175
rect 142857 50085 142885 50113
rect 142919 50085 142947 50113
rect 142981 50085 143009 50113
rect 143043 50085 143071 50113
rect 142857 50023 142885 50051
rect 142919 50023 142947 50051
rect 142981 50023 143009 50051
rect 143043 50023 143071 50051
rect 142857 49961 142885 49989
rect 142919 49961 142947 49989
rect 142981 49961 143009 49989
rect 143043 49961 143071 49989
rect 154179 50147 154207 50175
rect 154241 50147 154269 50175
rect 154179 50085 154207 50113
rect 154241 50085 154269 50113
rect 154179 50023 154207 50051
rect 154241 50023 154269 50051
rect 154179 49961 154207 49989
rect 154241 49961 154269 49989
rect 146499 47147 146527 47175
rect 146561 47147 146589 47175
rect 146499 47085 146527 47113
rect 146561 47085 146589 47113
rect 146499 47023 146527 47051
rect 146561 47023 146589 47051
rect 146499 46961 146527 46989
rect 146561 46961 146589 46989
rect 156357 47147 156385 47175
rect 156419 47147 156447 47175
rect 156481 47147 156509 47175
rect 156543 47147 156571 47175
rect 156357 47085 156385 47113
rect 156419 47085 156447 47113
rect 156481 47085 156509 47113
rect 156543 47085 156571 47113
rect 156357 47023 156385 47051
rect 156419 47023 156447 47051
rect 156481 47023 156509 47051
rect 156543 47023 156571 47051
rect 156357 46961 156385 46989
rect 156419 46961 156447 46989
rect 156481 46961 156509 46989
rect 156543 46961 156571 46989
rect 142857 41147 142885 41175
rect 142919 41147 142947 41175
rect 142981 41147 143009 41175
rect 143043 41147 143071 41175
rect 142857 41085 142885 41113
rect 142919 41085 142947 41113
rect 142981 41085 143009 41113
rect 143043 41085 143071 41113
rect 142857 41023 142885 41051
rect 142919 41023 142947 41051
rect 142981 41023 143009 41051
rect 143043 41023 143071 41051
rect 142857 40961 142885 40989
rect 142919 40961 142947 40989
rect 142981 40961 143009 40989
rect 143043 40961 143071 40989
rect 154179 41147 154207 41175
rect 154241 41147 154269 41175
rect 154179 41085 154207 41113
rect 154241 41085 154269 41113
rect 154179 41023 154207 41051
rect 154241 41023 154269 41051
rect 154179 40961 154207 40989
rect 154241 40961 154269 40989
rect 146499 38147 146527 38175
rect 146561 38147 146589 38175
rect 146499 38085 146527 38113
rect 146561 38085 146589 38113
rect 146499 38023 146527 38051
rect 146561 38023 146589 38051
rect 146499 37961 146527 37989
rect 146561 37961 146589 37989
rect 156357 38147 156385 38175
rect 156419 38147 156447 38175
rect 156481 38147 156509 38175
rect 156543 38147 156571 38175
rect 156357 38085 156385 38113
rect 156419 38085 156447 38113
rect 156481 38085 156509 38113
rect 156543 38085 156571 38113
rect 156357 38023 156385 38051
rect 156419 38023 156447 38051
rect 156481 38023 156509 38051
rect 156543 38023 156571 38051
rect 156357 37961 156385 37989
rect 156419 37961 156447 37989
rect 156481 37961 156509 37989
rect 156543 37961 156571 37989
rect 142857 32147 142885 32175
rect 142919 32147 142947 32175
rect 142981 32147 143009 32175
rect 143043 32147 143071 32175
rect 142857 32085 142885 32113
rect 142919 32085 142947 32113
rect 142981 32085 143009 32113
rect 143043 32085 143071 32113
rect 142857 32023 142885 32051
rect 142919 32023 142947 32051
rect 142981 32023 143009 32051
rect 143043 32023 143071 32051
rect 142857 31961 142885 31989
rect 142919 31961 142947 31989
rect 142981 31961 143009 31989
rect 143043 31961 143071 31989
rect 154179 32147 154207 32175
rect 154241 32147 154269 32175
rect 154179 32085 154207 32113
rect 154241 32085 154269 32113
rect 154179 32023 154207 32051
rect 154241 32023 154269 32051
rect 154179 31961 154207 31989
rect 154241 31961 154269 31989
rect 146499 29147 146527 29175
rect 146561 29147 146589 29175
rect 146499 29085 146527 29113
rect 146561 29085 146589 29113
rect 146499 29023 146527 29051
rect 146561 29023 146589 29051
rect 146499 28961 146527 28989
rect 146561 28961 146589 28989
rect 156357 29147 156385 29175
rect 156419 29147 156447 29175
rect 156481 29147 156509 29175
rect 156543 29147 156571 29175
rect 156357 29085 156385 29113
rect 156419 29085 156447 29113
rect 156481 29085 156509 29113
rect 156543 29085 156571 29113
rect 156357 29023 156385 29051
rect 156419 29023 156447 29051
rect 156481 29023 156509 29051
rect 156543 29023 156571 29051
rect 156357 28961 156385 28989
rect 156419 28961 156447 28989
rect 156481 28961 156509 28989
rect 156543 28961 156571 28989
rect 142857 23147 142885 23175
rect 142919 23147 142947 23175
rect 142981 23147 143009 23175
rect 143043 23147 143071 23175
rect 142857 23085 142885 23113
rect 142919 23085 142947 23113
rect 142981 23085 143009 23113
rect 143043 23085 143071 23113
rect 142857 23023 142885 23051
rect 142919 23023 142947 23051
rect 142981 23023 143009 23051
rect 143043 23023 143071 23051
rect 142857 22961 142885 22989
rect 142919 22961 142947 22989
rect 142981 22961 143009 22989
rect 143043 22961 143071 22989
rect 154179 23147 154207 23175
rect 154241 23147 154269 23175
rect 154179 23085 154207 23113
rect 154241 23085 154269 23113
rect 154179 23023 154207 23051
rect 154241 23023 154269 23051
rect 154179 22961 154207 22989
rect 154241 22961 154269 22989
rect 146499 20147 146527 20175
rect 146561 20147 146589 20175
rect 146499 20085 146527 20113
rect 146561 20085 146589 20113
rect 146499 20023 146527 20051
rect 146561 20023 146589 20051
rect 146499 19961 146527 19989
rect 146561 19961 146589 19989
rect 156357 20147 156385 20175
rect 156419 20147 156447 20175
rect 156481 20147 156509 20175
rect 156543 20147 156571 20175
rect 156357 20085 156385 20113
rect 156419 20085 156447 20113
rect 156481 20085 156509 20113
rect 156543 20085 156571 20113
rect 156357 20023 156385 20051
rect 156419 20023 156447 20051
rect 156481 20023 156509 20051
rect 156543 20023 156571 20051
rect 156357 19961 156385 19989
rect 156419 19961 156447 19989
rect 156481 19961 156509 19989
rect 156543 19961 156571 19989
rect 142857 14147 142885 14175
rect 142919 14147 142947 14175
rect 142981 14147 143009 14175
rect 143043 14147 143071 14175
rect 142857 14085 142885 14113
rect 142919 14085 142947 14113
rect 142981 14085 143009 14113
rect 143043 14085 143071 14113
rect 142857 14023 142885 14051
rect 142919 14023 142947 14051
rect 142981 14023 143009 14051
rect 143043 14023 143071 14051
rect 142857 13961 142885 13989
rect 142919 13961 142947 13989
rect 142981 13961 143009 13989
rect 143043 13961 143071 13989
rect 154179 14147 154207 14175
rect 154241 14147 154269 14175
rect 154179 14085 154207 14113
rect 154241 14085 154269 14113
rect 154179 14023 154207 14051
rect 154241 14023 154269 14051
rect 154179 13961 154207 13989
rect 154241 13961 154269 13989
rect 146499 11147 146527 11175
rect 146561 11147 146589 11175
rect 146499 11085 146527 11113
rect 146561 11085 146589 11113
rect 146499 11023 146527 11051
rect 146561 11023 146589 11051
rect 146499 10961 146527 10989
rect 146561 10961 146589 10989
rect 156357 11147 156385 11175
rect 156419 11147 156447 11175
rect 156481 11147 156509 11175
rect 156543 11147 156571 11175
rect 156357 11085 156385 11113
rect 156419 11085 156447 11113
rect 156481 11085 156509 11113
rect 156543 11085 156571 11113
rect 156357 11023 156385 11051
rect 156419 11023 156447 11051
rect 156481 11023 156509 11051
rect 156543 11023 156571 11051
rect 156357 10961 156385 10989
rect 156419 10961 156447 10989
rect 156481 10961 156509 10989
rect 156543 10961 156571 10989
rect 142857 5147 142885 5175
rect 142919 5147 142947 5175
rect 142981 5147 143009 5175
rect 143043 5147 143071 5175
rect 142857 5085 142885 5113
rect 142919 5085 142947 5113
rect 142981 5085 143009 5113
rect 143043 5085 143071 5113
rect 142857 5023 142885 5051
rect 142919 5023 142947 5051
rect 142981 5023 143009 5051
rect 143043 5023 143071 5051
rect 142857 4961 142885 4989
rect 142919 4961 142947 4989
rect 142981 4961 143009 4989
rect 143043 4961 143071 4989
rect 154179 5147 154207 5175
rect 154241 5147 154269 5175
rect 154179 5085 154207 5113
rect 154241 5085 154269 5113
rect 154179 5023 154207 5051
rect 154241 5023 154269 5051
rect 154179 4961 154207 4989
rect 154241 4961 154269 4989
rect 142857 -588 142885 -560
rect 142919 -588 142947 -560
rect 142981 -588 143009 -560
rect 143043 -588 143071 -560
rect 142857 -650 142885 -622
rect 142919 -650 142947 -622
rect 142981 -650 143009 -622
rect 143043 -650 143071 -622
rect 142857 -712 142885 -684
rect 142919 -712 142947 -684
rect 142981 -712 143009 -684
rect 143043 -712 143071 -684
rect 142857 -774 142885 -746
rect 142919 -774 142947 -746
rect 142981 -774 143009 -746
rect 143043 -774 143071 -746
rect 156357 2147 156385 2175
rect 156419 2147 156447 2175
rect 156481 2147 156509 2175
rect 156543 2147 156571 2175
rect 156357 2085 156385 2113
rect 156419 2085 156447 2113
rect 156481 2085 156509 2113
rect 156543 2085 156571 2113
rect 156357 2023 156385 2051
rect 156419 2023 156447 2051
rect 156481 2023 156509 2051
rect 156543 2023 156571 2051
rect 156357 1961 156385 1989
rect 156419 1961 156447 1989
rect 156481 1961 156509 1989
rect 156543 1961 156571 1989
rect 156357 -108 156385 -80
rect 156419 -108 156447 -80
rect 156481 -108 156509 -80
rect 156543 -108 156571 -80
rect 156357 -170 156385 -142
rect 156419 -170 156447 -142
rect 156481 -170 156509 -142
rect 156543 -170 156571 -142
rect 156357 -232 156385 -204
rect 156419 -232 156447 -204
rect 156481 -232 156509 -204
rect 156543 -232 156571 -204
rect 156357 -294 156385 -266
rect 156419 -294 156447 -266
rect 156481 -294 156509 -266
rect 156543 -294 156571 -266
rect 158217 299058 158245 299086
rect 158279 299058 158307 299086
rect 158341 299058 158369 299086
rect 158403 299058 158431 299086
rect 158217 298996 158245 299024
rect 158279 298996 158307 299024
rect 158341 298996 158369 299024
rect 158403 298996 158431 299024
rect 158217 298934 158245 298962
rect 158279 298934 158307 298962
rect 158341 298934 158369 298962
rect 158403 298934 158431 298962
rect 158217 298872 158245 298900
rect 158279 298872 158307 298900
rect 158341 298872 158369 298900
rect 158403 298872 158431 298900
rect 158217 293147 158245 293175
rect 158279 293147 158307 293175
rect 158341 293147 158369 293175
rect 158403 293147 158431 293175
rect 158217 293085 158245 293113
rect 158279 293085 158307 293113
rect 158341 293085 158369 293113
rect 158403 293085 158431 293113
rect 158217 293023 158245 293051
rect 158279 293023 158307 293051
rect 158341 293023 158369 293051
rect 158403 293023 158431 293051
rect 158217 292961 158245 292989
rect 158279 292961 158307 292989
rect 158341 292961 158369 292989
rect 158403 292961 158431 292989
rect 158217 284147 158245 284175
rect 158279 284147 158307 284175
rect 158341 284147 158369 284175
rect 158403 284147 158431 284175
rect 158217 284085 158245 284113
rect 158279 284085 158307 284113
rect 158341 284085 158369 284113
rect 158403 284085 158431 284113
rect 158217 284023 158245 284051
rect 158279 284023 158307 284051
rect 158341 284023 158369 284051
rect 158403 284023 158431 284051
rect 158217 283961 158245 283989
rect 158279 283961 158307 283989
rect 158341 283961 158369 283989
rect 158403 283961 158431 283989
rect 158217 275147 158245 275175
rect 158279 275147 158307 275175
rect 158341 275147 158369 275175
rect 158403 275147 158431 275175
rect 158217 275085 158245 275113
rect 158279 275085 158307 275113
rect 158341 275085 158369 275113
rect 158403 275085 158431 275113
rect 158217 275023 158245 275051
rect 158279 275023 158307 275051
rect 158341 275023 158369 275051
rect 158403 275023 158431 275051
rect 158217 274961 158245 274989
rect 158279 274961 158307 274989
rect 158341 274961 158369 274989
rect 158403 274961 158431 274989
rect 158217 266147 158245 266175
rect 158279 266147 158307 266175
rect 158341 266147 158369 266175
rect 158403 266147 158431 266175
rect 158217 266085 158245 266113
rect 158279 266085 158307 266113
rect 158341 266085 158369 266113
rect 158403 266085 158431 266113
rect 158217 266023 158245 266051
rect 158279 266023 158307 266051
rect 158341 266023 158369 266051
rect 158403 266023 158431 266051
rect 158217 265961 158245 265989
rect 158279 265961 158307 265989
rect 158341 265961 158369 265989
rect 158403 265961 158431 265989
rect 158217 257147 158245 257175
rect 158279 257147 158307 257175
rect 158341 257147 158369 257175
rect 158403 257147 158431 257175
rect 158217 257085 158245 257113
rect 158279 257085 158307 257113
rect 158341 257085 158369 257113
rect 158403 257085 158431 257113
rect 158217 257023 158245 257051
rect 158279 257023 158307 257051
rect 158341 257023 158369 257051
rect 158403 257023 158431 257051
rect 158217 256961 158245 256989
rect 158279 256961 158307 256989
rect 158341 256961 158369 256989
rect 158403 256961 158431 256989
rect 158217 248147 158245 248175
rect 158279 248147 158307 248175
rect 158341 248147 158369 248175
rect 158403 248147 158431 248175
rect 158217 248085 158245 248113
rect 158279 248085 158307 248113
rect 158341 248085 158369 248113
rect 158403 248085 158431 248113
rect 158217 248023 158245 248051
rect 158279 248023 158307 248051
rect 158341 248023 158369 248051
rect 158403 248023 158431 248051
rect 158217 247961 158245 247989
rect 158279 247961 158307 247989
rect 158341 247961 158369 247989
rect 158403 247961 158431 247989
rect 158217 239147 158245 239175
rect 158279 239147 158307 239175
rect 158341 239147 158369 239175
rect 158403 239147 158431 239175
rect 158217 239085 158245 239113
rect 158279 239085 158307 239113
rect 158341 239085 158369 239113
rect 158403 239085 158431 239113
rect 158217 239023 158245 239051
rect 158279 239023 158307 239051
rect 158341 239023 158369 239051
rect 158403 239023 158431 239051
rect 158217 238961 158245 238989
rect 158279 238961 158307 238989
rect 158341 238961 158369 238989
rect 158403 238961 158431 238989
rect 158217 230147 158245 230175
rect 158279 230147 158307 230175
rect 158341 230147 158369 230175
rect 158403 230147 158431 230175
rect 158217 230085 158245 230113
rect 158279 230085 158307 230113
rect 158341 230085 158369 230113
rect 158403 230085 158431 230113
rect 158217 230023 158245 230051
rect 158279 230023 158307 230051
rect 158341 230023 158369 230051
rect 158403 230023 158431 230051
rect 158217 229961 158245 229989
rect 158279 229961 158307 229989
rect 158341 229961 158369 229989
rect 158403 229961 158431 229989
rect 158217 221147 158245 221175
rect 158279 221147 158307 221175
rect 158341 221147 158369 221175
rect 158403 221147 158431 221175
rect 158217 221085 158245 221113
rect 158279 221085 158307 221113
rect 158341 221085 158369 221113
rect 158403 221085 158431 221113
rect 158217 221023 158245 221051
rect 158279 221023 158307 221051
rect 158341 221023 158369 221051
rect 158403 221023 158431 221051
rect 158217 220961 158245 220989
rect 158279 220961 158307 220989
rect 158341 220961 158369 220989
rect 158403 220961 158431 220989
rect 158217 212147 158245 212175
rect 158279 212147 158307 212175
rect 158341 212147 158369 212175
rect 158403 212147 158431 212175
rect 158217 212085 158245 212113
rect 158279 212085 158307 212113
rect 158341 212085 158369 212113
rect 158403 212085 158431 212113
rect 158217 212023 158245 212051
rect 158279 212023 158307 212051
rect 158341 212023 158369 212051
rect 158403 212023 158431 212051
rect 158217 211961 158245 211989
rect 158279 211961 158307 211989
rect 158341 211961 158369 211989
rect 158403 211961 158431 211989
rect 158217 203147 158245 203175
rect 158279 203147 158307 203175
rect 158341 203147 158369 203175
rect 158403 203147 158431 203175
rect 158217 203085 158245 203113
rect 158279 203085 158307 203113
rect 158341 203085 158369 203113
rect 158403 203085 158431 203113
rect 158217 203023 158245 203051
rect 158279 203023 158307 203051
rect 158341 203023 158369 203051
rect 158403 203023 158431 203051
rect 158217 202961 158245 202989
rect 158279 202961 158307 202989
rect 158341 202961 158369 202989
rect 158403 202961 158431 202989
rect 158217 194147 158245 194175
rect 158279 194147 158307 194175
rect 158341 194147 158369 194175
rect 158403 194147 158431 194175
rect 158217 194085 158245 194113
rect 158279 194085 158307 194113
rect 158341 194085 158369 194113
rect 158403 194085 158431 194113
rect 158217 194023 158245 194051
rect 158279 194023 158307 194051
rect 158341 194023 158369 194051
rect 158403 194023 158431 194051
rect 158217 193961 158245 193989
rect 158279 193961 158307 193989
rect 158341 193961 158369 193989
rect 158403 193961 158431 193989
rect 158217 185147 158245 185175
rect 158279 185147 158307 185175
rect 158341 185147 158369 185175
rect 158403 185147 158431 185175
rect 158217 185085 158245 185113
rect 158279 185085 158307 185113
rect 158341 185085 158369 185113
rect 158403 185085 158431 185113
rect 158217 185023 158245 185051
rect 158279 185023 158307 185051
rect 158341 185023 158369 185051
rect 158403 185023 158431 185051
rect 158217 184961 158245 184989
rect 158279 184961 158307 184989
rect 158341 184961 158369 184989
rect 158403 184961 158431 184989
rect 158217 176147 158245 176175
rect 158279 176147 158307 176175
rect 158341 176147 158369 176175
rect 158403 176147 158431 176175
rect 158217 176085 158245 176113
rect 158279 176085 158307 176113
rect 158341 176085 158369 176113
rect 158403 176085 158431 176113
rect 158217 176023 158245 176051
rect 158279 176023 158307 176051
rect 158341 176023 158369 176051
rect 158403 176023 158431 176051
rect 158217 175961 158245 175989
rect 158279 175961 158307 175989
rect 158341 175961 158369 175989
rect 158403 175961 158431 175989
rect 171717 298578 171745 298606
rect 171779 298578 171807 298606
rect 171841 298578 171869 298606
rect 171903 298578 171931 298606
rect 171717 298516 171745 298544
rect 171779 298516 171807 298544
rect 171841 298516 171869 298544
rect 171903 298516 171931 298544
rect 171717 298454 171745 298482
rect 171779 298454 171807 298482
rect 171841 298454 171869 298482
rect 171903 298454 171931 298482
rect 171717 298392 171745 298420
rect 171779 298392 171807 298420
rect 171841 298392 171869 298420
rect 171903 298392 171931 298420
rect 171717 290147 171745 290175
rect 171779 290147 171807 290175
rect 171841 290147 171869 290175
rect 171903 290147 171931 290175
rect 171717 290085 171745 290113
rect 171779 290085 171807 290113
rect 171841 290085 171869 290113
rect 171903 290085 171931 290113
rect 171717 290023 171745 290051
rect 171779 290023 171807 290051
rect 171841 290023 171869 290051
rect 171903 290023 171931 290051
rect 171717 289961 171745 289989
rect 171779 289961 171807 289989
rect 171841 289961 171869 289989
rect 171903 289961 171931 289989
rect 171717 281147 171745 281175
rect 171779 281147 171807 281175
rect 171841 281147 171869 281175
rect 171903 281147 171931 281175
rect 171717 281085 171745 281113
rect 171779 281085 171807 281113
rect 171841 281085 171869 281113
rect 171903 281085 171931 281113
rect 171717 281023 171745 281051
rect 171779 281023 171807 281051
rect 171841 281023 171869 281051
rect 171903 281023 171931 281051
rect 171717 280961 171745 280989
rect 171779 280961 171807 280989
rect 171841 280961 171869 280989
rect 171903 280961 171931 280989
rect 171717 272147 171745 272175
rect 171779 272147 171807 272175
rect 171841 272147 171869 272175
rect 171903 272147 171931 272175
rect 171717 272085 171745 272113
rect 171779 272085 171807 272113
rect 171841 272085 171869 272113
rect 171903 272085 171931 272113
rect 171717 272023 171745 272051
rect 171779 272023 171807 272051
rect 171841 272023 171869 272051
rect 171903 272023 171931 272051
rect 171717 271961 171745 271989
rect 171779 271961 171807 271989
rect 171841 271961 171869 271989
rect 171903 271961 171931 271989
rect 171717 263147 171745 263175
rect 171779 263147 171807 263175
rect 171841 263147 171869 263175
rect 171903 263147 171931 263175
rect 171717 263085 171745 263113
rect 171779 263085 171807 263113
rect 171841 263085 171869 263113
rect 171903 263085 171931 263113
rect 171717 263023 171745 263051
rect 171779 263023 171807 263051
rect 171841 263023 171869 263051
rect 171903 263023 171931 263051
rect 171717 262961 171745 262989
rect 171779 262961 171807 262989
rect 171841 262961 171869 262989
rect 171903 262961 171931 262989
rect 171717 254147 171745 254175
rect 171779 254147 171807 254175
rect 171841 254147 171869 254175
rect 171903 254147 171931 254175
rect 171717 254085 171745 254113
rect 171779 254085 171807 254113
rect 171841 254085 171869 254113
rect 171903 254085 171931 254113
rect 171717 254023 171745 254051
rect 171779 254023 171807 254051
rect 171841 254023 171869 254051
rect 171903 254023 171931 254051
rect 171717 253961 171745 253989
rect 171779 253961 171807 253989
rect 171841 253961 171869 253989
rect 171903 253961 171931 253989
rect 171717 245147 171745 245175
rect 171779 245147 171807 245175
rect 171841 245147 171869 245175
rect 171903 245147 171931 245175
rect 171717 245085 171745 245113
rect 171779 245085 171807 245113
rect 171841 245085 171869 245113
rect 171903 245085 171931 245113
rect 171717 245023 171745 245051
rect 171779 245023 171807 245051
rect 171841 245023 171869 245051
rect 171903 245023 171931 245051
rect 171717 244961 171745 244989
rect 171779 244961 171807 244989
rect 171841 244961 171869 244989
rect 171903 244961 171931 244989
rect 171717 236147 171745 236175
rect 171779 236147 171807 236175
rect 171841 236147 171869 236175
rect 171903 236147 171931 236175
rect 171717 236085 171745 236113
rect 171779 236085 171807 236113
rect 171841 236085 171869 236113
rect 171903 236085 171931 236113
rect 171717 236023 171745 236051
rect 171779 236023 171807 236051
rect 171841 236023 171869 236051
rect 171903 236023 171931 236051
rect 171717 235961 171745 235989
rect 171779 235961 171807 235989
rect 171841 235961 171869 235989
rect 171903 235961 171931 235989
rect 171717 227147 171745 227175
rect 171779 227147 171807 227175
rect 171841 227147 171869 227175
rect 171903 227147 171931 227175
rect 171717 227085 171745 227113
rect 171779 227085 171807 227113
rect 171841 227085 171869 227113
rect 171903 227085 171931 227113
rect 171717 227023 171745 227051
rect 171779 227023 171807 227051
rect 171841 227023 171869 227051
rect 171903 227023 171931 227051
rect 171717 226961 171745 226989
rect 171779 226961 171807 226989
rect 171841 226961 171869 226989
rect 171903 226961 171931 226989
rect 171717 218147 171745 218175
rect 171779 218147 171807 218175
rect 171841 218147 171869 218175
rect 171903 218147 171931 218175
rect 171717 218085 171745 218113
rect 171779 218085 171807 218113
rect 171841 218085 171869 218113
rect 171903 218085 171931 218113
rect 171717 218023 171745 218051
rect 171779 218023 171807 218051
rect 171841 218023 171869 218051
rect 171903 218023 171931 218051
rect 171717 217961 171745 217989
rect 171779 217961 171807 217989
rect 171841 217961 171869 217989
rect 171903 217961 171931 217989
rect 171717 209147 171745 209175
rect 171779 209147 171807 209175
rect 171841 209147 171869 209175
rect 171903 209147 171931 209175
rect 171717 209085 171745 209113
rect 171779 209085 171807 209113
rect 171841 209085 171869 209113
rect 171903 209085 171931 209113
rect 171717 209023 171745 209051
rect 171779 209023 171807 209051
rect 171841 209023 171869 209051
rect 171903 209023 171931 209051
rect 171717 208961 171745 208989
rect 171779 208961 171807 208989
rect 171841 208961 171869 208989
rect 171903 208961 171931 208989
rect 171717 200147 171745 200175
rect 171779 200147 171807 200175
rect 171841 200147 171869 200175
rect 171903 200147 171931 200175
rect 171717 200085 171745 200113
rect 171779 200085 171807 200113
rect 171841 200085 171869 200113
rect 171903 200085 171931 200113
rect 171717 200023 171745 200051
rect 171779 200023 171807 200051
rect 171841 200023 171869 200051
rect 171903 200023 171931 200051
rect 171717 199961 171745 199989
rect 171779 199961 171807 199989
rect 171841 199961 171869 199989
rect 171903 199961 171931 199989
rect 171717 191147 171745 191175
rect 171779 191147 171807 191175
rect 171841 191147 171869 191175
rect 171903 191147 171931 191175
rect 171717 191085 171745 191113
rect 171779 191085 171807 191113
rect 171841 191085 171869 191113
rect 171903 191085 171931 191113
rect 171717 191023 171745 191051
rect 171779 191023 171807 191051
rect 171841 191023 171869 191051
rect 171903 191023 171931 191051
rect 171717 190961 171745 190989
rect 171779 190961 171807 190989
rect 171841 190961 171869 190989
rect 171903 190961 171931 190989
rect 171717 182147 171745 182175
rect 171779 182147 171807 182175
rect 171841 182147 171869 182175
rect 171903 182147 171931 182175
rect 171717 182085 171745 182113
rect 171779 182085 171807 182113
rect 171841 182085 171869 182113
rect 171903 182085 171931 182113
rect 171717 182023 171745 182051
rect 171779 182023 171807 182051
rect 171841 182023 171869 182051
rect 171903 182023 171931 182051
rect 171717 181961 171745 181989
rect 171779 181961 171807 181989
rect 171841 181961 171869 181989
rect 171903 181961 171931 181989
rect 161859 173147 161887 173175
rect 161921 173147 161949 173175
rect 161859 173085 161887 173113
rect 161921 173085 161949 173113
rect 161859 173023 161887 173051
rect 161921 173023 161949 173051
rect 161859 172961 161887 172989
rect 161921 172961 161949 172989
rect 171717 173147 171745 173175
rect 171779 173147 171807 173175
rect 171841 173147 171869 173175
rect 171903 173147 171931 173175
rect 171717 173085 171745 173113
rect 171779 173085 171807 173113
rect 171841 173085 171869 173113
rect 171903 173085 171931 173113
rect 171717 173023 171745 173051
rect 171779 173023 171807 173051
rect 171841 173023 171869 173051
rect 171903 173023 171931 173051
rect 171717 172961 171745 172989
rect 171779 172961 171807 172989
rect 171841 172961 171869 172989
rect 171903 172961 171931 172989
rect 158217 167147 158245 167175
rect 158279 167147 158307 167175
rect 158341 167147 158369 167175
rect 158403 167147 158431 167175
rect 158217 167085 158245 167113
rect 158279 167085 158307 167113
rect 158341 167085 158369 167113
rect 158403 167085 158431 167113
rect 158217 167023 158245 167051
rect 158279 167023 158307 167051
rect 158341 167023 158369 167051
rect 158403 167023 158431 167051
rect 158217 166961 158245 166989
rect 158279 166961 158307 166989
rect 158341 166961 158369 166989
rect 158403 166961 158431 166989
rect 169539 167147 169567 167175
rect 169601 167147 169629 167175
rect 169539 167085 169567 167113
rect 169601 167085 169629 167113
rect 169539 167023 169567 167051
rect 169601 167023 169629 167051
rect 169539 166961 169567 166989
rect 169601 166961 169629 166989
rect 161859 164147 161887 164175
rect 161921 164147 161949 164175
rect 161859 164085 161887 164113
rect 161921 164085 161949 164113
rect 161859 164023 161887 164051
rect 161921 164023 161949 164051
rect 161859 163961 161887 163989
rect 161921 163961 161949 163989
rect 171717 164147 171745 164175
rect 171779 164147 171807 164175
rect 171841 164147 171869 164175
rect 171903 164147 171931 164175
rect 171717 164085 171745 164113
rect 171779 164085 171807 164113
rect 171841 164085 171869 164113
rect 171903 164085 171931 164113
rect 171717 164023 171745 164051
rect 171779 164023 171807 164051
rect 171841 164023 171869 164051
rect 171903 164023 171931 164051
rect 171717 163961 171745 163989
rect 171779 163961 171807 163989
rect 171841 163961 171869 163989
rect 171903 163961 171931 163989
rect 158217 158147 158245 158175
rect 158279 158147 158307 158175
rect 158341 158147 158369 158175
rect 158403 158147 158431 158175
rect 158217 158085 158245 158113
rect 158279 158085 158307 158113
rect 158341 158085 158369 158113
rect 158403 158085 158431 158113
rect 158217 158023 158245 158051
rect 158279 158023 158307 158051
rect 158341 158023 158369 158051
rect 158403 158023 158431 158051
rect 158217 157961 158245 157989
rect 158279 157961 158307 157989
rect 158341 157961 158369 157989
rect 158403 157961 158431 157989
rect 169539 158147 169567 158175
rect 169601 158147 169629 158175
rect 169539 158085 169567 158113
rect 169601 158085 169629 158113
rect 169539 158023 169567 158051
rect 169601 158023 169629 158051
rect 169539 157961 169567 157989
rect 169601 157961 169629 157989
rect 161859 155147 161887 155175
rect 161921 155147 161949 155175
rect 161859 155085 161887 155113
rect 161921 155085 161949 155113
rect 161859 155023 161887 155051
rect 161921 155023 161949 155051
rect 161859 154961 161887 154989
rect 161921 154961 161949 154989
rect 171717 155147 171745 155175
rect 171779 155147 171807 155175
rect 171841 155147 171869 155175
rect 171903 155147 171931 155175
rect 171717 155085 171745 155113
rect 171779 155085 171807 155113
rect 171841 155085 171869 155113
rect 171903 155085 171931 155113
rect 171717 155023 171745 155051
rect 171779 155023 171807 155051
rect 171841 155023 171869 155051
rect 171903 155023 171931 155051
rect 171717 154961 171745 154989
rect 171779 154961 171807 154989
rect 171841 154961 171869 154989
rect 171903 154961 171931 154989
rect 158217 149147 158245 149175
rect 158279 149147 158307 149175
rect 158341 149147 158369 149175
rect 158403 149147 158431 149175
rect 158217 149085 158245 149113
rect 158279 149085 158307 149113
rect 158341 149085 158369 149113
rect 158403 149085 158431 149113
rect 158217 149023 158245 149051
rect 158279 149023 158307 149051
rect 158341 149023 158369 149051
rect 158403 149023 158431 149051
rect 158217 148961 158245 148989
rect 158279 148961 158307 148989
rect 158341 148961 158369 148989
rect 158403 148961 158431 148989
rect 169539 149147 169567 149175
rect 169601 149147 169629 149175
rect 169539 149085 169567 149113
rect 169601 149085 169629 149113
rect 169539 149023 169567 149051
rect 169601 149023 169629 149051
rect 169539 148961 169567 148989
rect 169601 148961 169629 148989
rect 161859 146147 161887 146175
rect 161921 146147 161949 146175
rect 161859 146085 161887 146113
rect 161921 146085 161949 146113
rect 161859 146023 161887 146051
rect 161921 146023 161949 146051
rect 161859 145961 161887 145989
rect 161921 145961 161949 145989
rect 171717 146147 171745 146175
rect 171779 146147 171807 146175
rect 171841 146147 171869 146175
rect 171903 146147 171931 146175
rect 171717 146085 171745 146113
rect 171779 146085 171807 146113
rect 171841 146085 171869 146113
rect 171903 146085 171931 146113
rect 171717 146023 171745 146051
rect 171779 146023 171807 146051
rect 171841 146023 171869 146051
rect 171903 146023 171931 146051
rect 171717 145961 171745 145989
rect 171779 145961 171807 145989
rect 171841 145961 171869 145989
rect 171903 145961 171931 145989
rect 158217 140147 158245 140175
rect 158279 140147 158307 140175
rect 158341 140147 158369 140175
rect 158403 140147 158431 140175
rect 158217 140085 158245 140113
rect 158279 140085 158307 140113
rect 158341 140085 158369 140113
rect 158403 140085 158431 140113
rect 158217 140023 158245 140051
rect 158279 140023 158307 140051
rect 158341 140023 158369 140051
rect 158403 140023 158431 140051
rect 158217 139961 158245 139989
rect 158279 139961 158307 139989
rect 158341 139961 158369 139989
rect 158403 139961 158431 139989
rect 169539 140147 169567 140175
rect 169601 140147 169629 140175
rect 169539 140085 169567 140113
rect 169601 140085 169629 140113
rect 169539 140023 169567 140051
rect 169601 140023 169629 140051
rect 169539 139961 169567 139989
rect 169601 139961 169629 139989
rect 161859 137147 161887 137175
rect 161921 137147 161949 137175
rect 161859 137085 161887 137113
rect 161921 137085 161949 137113
rect 161859 137023 161887 137051
rect 161921 137023 161949 137051
rect 161859 136961 161887 136989
rect 161921 136961 161949 136989
rect 171717 137147 171745 137175
rect 171779 137147 171807 137175
rect 171841 137147 171869 137175
rect 171903 137147 171931 137175
rect 171717 137085 171745 137113
rect 171779 137085 171807 137113
rect 171841 137085 171869 137113
rect 171903 137085 171931 137113
rect 171717 137023 171745 137051
rect 171779 137023 171807 137051
rect 171841 137023 171869 137051
rect 171903 137023 171931 137051
rect 171717 136961 171745 136989
rect 171779 136961 171807 136989
rect 171841 136961 171869 136989
rect 171903 136961 171931 136989
rect 158217 131147 158245 131175
rect 158279 131147 158307 131175
rect 158341 131147 158369 131175
rect 158403 131147 158431 131175
rect 158217 131085 158245 131113
rect 158279 131085 158307 131113
rect 158341 131085 158369 131113
rect 158403 131085 158431 131113
rect 158217 131023 158245 131051
rect 158279 131023 158307 131051
rect 158341 131023 158369 131051
rect 158403 131023 158431 131051
rect 158217 130961 158245 130989
rect 158279 130961 158307 130989
rect 158341 130961 158369 130989
rect 158403 130961 158431 130989
rect 169539 131147 169567 131175
rect 169601 131147 169629 131175
rect 169539 131085 169567 131113
rect 169601 131085 169629 131113
rect 169539 131023 169567 131051
rect 169601 131023 169629 131051
rect 169539 130961 169567 130989
rect 169601 130961 169629 130989
rect 161859 128147 161887 128175
rect 161921 128147 161949 128175
rect 161859 128085 161887 128113
rect 161921 128085 161949 128113
rect 161859 128023 161887 128051
rect 161921 128023 161949 128051
rect 161859 127961 161887 127989
rect 161921 127961 161949 127989
rect 171717 128147 171745 128175
rect 171779 128147 171807 128175
rect 171841 128147 171869 128175
rect 171903 128147 171931 128175
rect 171717 128085 171745 128113
rect 171779 128085 171807 128113
rect 171841 128085 171869 128113
rect 171903 128085 171931 128113
rect 171717 128023 171745 128051
rect 171779 128023 171807 128051
rect 171841 128023 171869 128051
rect 171903 128023 171931 128051
rect 171717 127961 171745 127989
rect 171779 127961 171807 127989
rect 171841 127961 171869 127989
rect 171903 127961 171931 127989
rect 158217 122147 158245 122175
rect 158279 122147 158307 122175
rect 158341 122147 158369 122175
rect 158403 122147 158431 122175
rect 158217 122085 158245 122113
rect 158279 122085 158307 122113
rect 158341 122085 158369 122113
rect 158403 122085 158431 122113
rect 158217 122023 158245 122051
rect 158279 122023 158307 122051
rect 158341 122023 158369 122051
rect 158403 122023 158431 122051
rect 158217 121961 158245 121989
rect 158279 121961 158307 121989
rect 158341 121961 158369 121989
rect 158403 121961 158431 121989
rect 169539 122147 169567 122175
rect 169601 122147 169629 122175
rect 169539 122085 169567 122113
rect 169601 122085 169629 122113
rect 169539 122023 169567 122051
rect 169601 122023 169629 122051
rect 169539 121961 169567 121989
rect 169601 121961 169629 121989
rect 161859 119147 161887 119175
rect 161921 119147 161949 119175
rect 161859 119085 161887 119113
rect 161921 119085 161949 119113
rect 161859 119023 161887 119051
rect 161921 119023 161949 119051
rect 161859 118961 161887 118989
rect 161921 118961 161949 118989
rect 171717 119147 171745 119175
rect 171779 119147 171807 119175
rect 171841 119147 171869 119175
rect 171903 119147 171931 119175
rect 171717 119085 171745 119113
rect 171779 119085 171807 119113
rect 171841 119085 171869 119113
rect 171903 119085 171931 119113
rect 171717 119023 171745 119051
rect 171779 119023 171807 119051
rect 171841 119023 171869 119051
rect 171903 119023 171931 119051
rect 171717 118961 171745 118989
rect 171779 118961 171807 118989
rect 171841 118961 171869 118989
rect 171903 118961 171931 118989
rect 158217 113147 158245 113175
rect 158279 113147 158307 113175
rect 158341 113147 158369 113175
rect 158403 113147 158431 113175
rect 158217 113085 158245 113113
rect 158279 113085 158307 113113
rect 158341 113085 158369 113113
rect 158403 113085 158431 113113
rect 158217 113023 158245 113051
rect 158279 113023 158307 113051
rect 158341 113023 158369 113051
rect 158403 113023 158431 113051
rect 158217 112961 158245 112989
rect 158279 112961 158307 112989
rect 158341 112961 158369 112989
rect 158403 112961 158431 112989
rect 169539 113147 169567 113175
rect 169601 113147 169629 113175
rect 169539 113085 169567 113113
rect 169601 113085 169629 113113
rect 169539 113023 169567 113051
rect 169601 113023 169629 113051
rect 169539 112961 169567 112989
rect 169601 112961 169629 112989
rect 161859 110147 161887 110175
rect 161921 110147 161949 110175
rect 161859 110085 161887 110113
rect 161921 110085 161949 110113
rect 161859 110023 161887 110051
rect 161921 110023 161949 110051
rect 161859 109961 161887 109989
rect 161921 109961 161949 109989
rect 171717 110147 171745 110175
rect 171779 110147 171807 110175
rect 171841 110147 171869 110175
rect 171903 110147 171931 110175
rect 171717 110085 171745 110113
rect 171779 110085 171807 110113
rect 171841 110085 171869 110113
rect 171903 110085 171931 110113
rect 171717 110023 171745 110051
rect 171779 110023 171807 110051
rect 171841 110023 171869 110051
rect 171903 110023 171931 110051
rect 171717 109961 171745 109989
rect 171779 109961 171807 109989
rect 171841 109961 171869 109989
rect 171903 109961 171931 109989
rect 158217 104147 158245 104175
rect 158279 104147 158307 104175
rect 158341 104147 158369 104175
rect 158403 104147 158431 104175
rect 158217 104085 158245 104113
rect 158279 104085 158307 104113
rect 158341 104085 158369 104113
rect 158403 104085 158431 104113
rect 158217 104023 158245 104051
rect 158279 104023 158307 104051
rect 158341 104023 158369 104051
rect 158403 104023 158431 104051
rect 158217 103961 158245 103989
rect 158279 103961 158307 103989
rect 158341 103961 158369 103989
rect 158403 103961 158431 103989
rect 169539 104147 169567 104175
rect 169601 104147 169629 104175
rect 169539 104085 169567 104113
rect 169601 104085 169629 104113
rect 169539 104023 169567 104051
rect 169601 104023 169629 104051
rect 169539 103961 169567 103989
rect 169601 103961 169629 103989
rect 161859 101147 161887 101175
rect 161921 101147 161949 101175
rect 161859 101085 161887 101113
rect 161921 101085 161949 101113
rect 161859 101023 161887 101051
rect 161921 101023 161949 101051
rect 161859 100961 161887 100989
rect 161921 100961 161949 100989
rect 171717 101147 171745 101175
rect 171779 101147 171807 101175
rect 171841 101147 171869 101175
rect 171903 101147 171931 101175
rect 171717 101085 171745 101113
rect 171779 101085 171807 101113
rect 171841 101085 171869 101113
rect 171903 101085 171931 101113
rect 171717 101023 171745 101051
rect 171779 101023 171807 101051
rect 171841 101023 171869 101051
rect 171903 101023 171931 101051
rect 171717 100961 171745 100989
rect 171779 100961 171807 100989
rect 171841 100961 171869 100989
rect 171903 100961 171931 100989
rect 158217 95147 158245 95175
rect 158279 95147 158307 95175
rect 158341 95147 158369 95175
rect 158403 95147 158431 95175
rect 158217 95085 158245 95113
rect 158279 95085 158307 95113
rect 158341 95085 158369 95113
rect 158403 95085 158431 95113
rect 158217 95023 158245 95051
rect 158279 95023 158307 95051
rect 158341 95023 158369 95051
rect 158403 95023 158431 95051
rect 158217 94961 158245 94989
rect 158279 94961 158307 94989
rect 158341 94961 158369 94989
rect 158403 94961 158431 94989
rect 169539 95147 169567 95175
rect 169601 95147 169629 95175
rect 169539 95085 169567 95113
rect 169601 95085 169629 95113
rect 169539 95023 169567 95051
rect 169601 95023 169629 95051
rect 169539 94961 169567 94989
rect 169601 94961 169629 94989
rect 161859 92147 161887 92175
rect 161921 92147 161949 92175
rect 161859 92085 161887 92113
rect 161921 92085 161949 92113
rect 161859 92023 161887 92051
rect 161921 92023 161949 92051
rect 161859 91961 161887 91989
rect 161921 91961 161949 91989
rect 171717 92147 171745 92175
rect 171779 92147 171807 92175
rect 171841 92147 171869 92175
rect 171903 92147 171931 92175
rect 171717 92085 171745 92113
rect 171779 92085 171807 92113
rect 171841 92085 171869 92113
rect 171903 92085 171931 92113
rect 171717 92023 171745 92051
rect 171779 92023 171807 92051
rect 171841 92023 171869 92051
rect 171903 92023 171931 92051
rect 171717 91961 171745 91989
rect 171779 91961 171807 91989
rect 171841 91961 171869 91989
rect 171903 91961 171931 91989
rect 158217 86147 158245 86175
rect 158279 86147 158307 86175
rect 158341 86147 158369 86175
rect 158403 86147 158431 86175
rect 158217 86085 158245 86113
rect 158279 86085 158307 86113
rect 158341 86085 158369 86113
rect 158403 86085 158431 86113
rect 158217 86023 158245 86051
rect 158279 86023 158307 86051
rect 158341 86023 158369 86051
rect 158403 86023 158431 86051
rect 158217 85961 158245 85989
rect 158279 85961 158307 85989
rect 158341 85961 158369 85989
rect 158403 85961 158431 85989
rect 169539 86147 169567 86175
rect 169601 86147 169629 86175
rect 169539 86085 169567 86113
rect 169601 86085 169629 86113
rect 169539 86023 169567 86051
rect 169601 86023 169629 86051
rect 169539 85961 169567 85989
rect 169601 85961 169629 85989
rect 161859 83147 161887 83175
rect 161921 83147 161949 83175
rect 161859 83085 161887 83113
rect 161921 83085 161949 83113
rect 161859 83023 161887 83051
rect 161921 83023 161949 83051
rect 161859 82961 161887 82989
rect 161921 82961 161949 82989
rect 171717 83147 171745 83175
rect 171779 83147 171807 83175
rect 171841 83147 171869 83175
rect 171903 83147 171931 83175
rect 171717 83085 171745 83113
rect 171779 83085 171807 83113
rect 171841 83085 171869 83113
rect 171903 83085 171931 83113
rect 171717 83023 171745 83051
rect 171779 83023 171807 83051
rect 171841 83023 171869 83051
rect 171903 83023 171931 83051
rect 171717 82961 171745 82989
rect 171779 82961 171807 82989
rect 171841 82961 171869 82989
rect 171903 82961 171931 82989
rect 158217 77147 158245 77175
rect 158279 77147 158307 77175
rect 158341 77147 158369 77175
rect 158403 77147 158431 77175
rect 158217 77085 158245 77113
rect 158279 77085 158307 77113
rect 158341 77085 158369 77113
rect 158403 77085 158431 77113
rect 158217 77023 158245 77051
rect 158279 77023 158307 77051
rect 158341 77023 158369 77051
rect 158403 77023 158431 77051
rect 158217 76961 158245 76989
rect 158279 76961 158307 76989
rect 158341 76961 158369 76989
rect 158403 76961 158431 76989
rect 169539 77147 169567 77175
rect 169601 77147 169629 77175
rect 169539 77085 169567 77113
rect 169601 77085 169629 77113
rect 169539 77023 169567 77051
rect 169601 77023 169629 77051
rect 169539 76961 169567 76989
rect 169601 76961 169629 76989
rect 161859 74147 161887 74175
rect 161921 74147 161949 74175
rect 161859 74085 161887 74113
rect 161921 74085 161949 74113
rect 161859 74023 161887 74051
rect 161921 74023 161949 74051
rect 161859 73961 161887 73989
rect 161921 73961 161949 73989
rect 171717 74147 171745 74175
rect 171779 74147 171807 74175
rect 171841 74147 171869 74175
rect 171903 74147 171931 74175
rect 171717 74085 171745 74113
rect 171779 74085 171807 74113
rect 171841 74085 171869 74113
rect 171903 74085 171931 74113
rect 171717 74023 171745 74051
rect 171779 74023 171807 74051
rect 171841 74023 171869 74051
rect 171903 74023 171931 74051
rect 171717 73961 171745 73989
rect 171779 73961 171807 73989
rect 171841 73961 171869 73989
rect 171903 73961 171931 73989
rect 158217 68147 158245 68175
rect 158279 68147 158307 68175
rect 158341 68147 158369 68175
rect 158403 68147 158431 68175
rect 158217 68085 158245 68113
rect 158279 68085 158307 68113
rect 158341 68085 158369 68113
rect 158403 68085 158431 68113
rect 158217 68023 158245 68051
rect 158279 68023 158307 68051
rect 158341 68023 158369 68051
rect 158403 68023 158431 68051
rect 158217 67961 158245 67989
rect 158279 67961 158307 67989
rect 158341 67961 158369 67989
rect 158403 67961 158431 67989
rect 169539 68147 169567 68175
rect 169601 68147 169629 68175
rect 169539 68085 169567 68113
rect 169601 68085 169629 68113
rect 169539 68023 169567 68051
rect 169601 68023 169629 68051
rect 169539 67961 169567 67989
rect 169601 67961 169629 67989
rect 161859 65147 161887 65175
rect 161921 65147 161949 65175
rect 161859 65085 161887 65113
rect 161921 65085 161949 65113
rect 161859 65023 161887 65051
rect 161921 65023 161949 65051
rect 161859 64961 161887 64989
rect 161921 64961 161949 64989
rect 171717 65147 171745 65175
rect 171779 65147 171807 65175
rect 171841 65147 171869 65175
rect 171903 65147 171931 65175
rect 171717 65085 171745 65113
rect 171779 65085 171807 65113
rect 171841 65085 171869 65113
rect 171903 65085 171931 65113
rect 171717 65023 171745 65051
rect 171779 65023 171807 65051
rect 171841 65023 171869 65051
rect 171903 65023 171931 65051
rect 171717 64961 171745 64989
rect 171779 64961 171807 64989
rect 171841 64961 171869 64989
rect 171903 64961 171931 64989
rect 158217 59147 158245 59175
rect 158279 59147 158307 59175
rect 158341 59147 158369 59175
rect 158403 59147 158431 59175
rect 158217 59085 158245 59113
rect 158279 59085 158307 59113
rect 158341 59085 158369 59113
rect 158403 59085 158431 59113
rect 158217 59023 158245 59051
rect 158279 59023 158307 59051
rect 158341 59023 158369 59051
rect 158403 59023 158431 59051
rect 158217 58961 158245 58989
rect 158279 58961 158307 58989
rect 158341 58961 158369 58989
rect 158403 58961 158431 58989
rect 169539 59147 169567 59175
rect 169601 59147 169629 59175
rect 169539 59085 169567 59113
rect 169601 59085 169629 59113
rect 169539 59023 169567 59051
rect 169601 59023 169629 59051
rect 169539 58961 169567 58989
rect 169601 58961 169629 58989
rect 161859 56147 161887 56175
rect 161921 56147 161949 56175
rect 161859 56085 161887 56113
rect 161921 56085 161949 56113
rect 161859 56023 161887 56051
rect 161921 56023 161949 56051
rect 161859 55961 161887 55989
rect 161921 55961 161949 55989
rect 171717 56147 171745 56175
rect 171779 56147 171807 56175
rect 171841 56147 171869 56175
rect 171903 56147 171931 56175
rect 171717 56085 171745 56113
rect 171779 56085 171807 56113
rect 171841 56085 171869 56113
rect 171903 56085 171931 56113
rect 171717 56023 171745 56051
rect 171779 56023 171807 56051
rect 171841 56023 171869 56051
rect 171903 56023 171931 56051
rect 171717 55961 171745 55989
rect 171779 55961 171807 55989
rect 171841 55961 171869 55989
rect 171903 55961 171931 55989
rect 158217 50147 158245 50175
rect 158279 50147 158307 50175
rect 158341 50147 158369 50175
rect 158403 50147 158431 50175
rect 158217 50085 158245 50113
rect 158279 50085 158307 50113
rect 158341 50085 158369 50113
rect 158403 50085 158431 50113
rect 158217 50023 158245 50051
rect 158279 50023 158307 50051
rect 158341 50023 158369 50051
rect 158403 50023 158431 50051
rect 158217 49961 158245 49989
rect 158279 49961 158307 49989
rect 158341 49961 158369 49989
rect 158403 49961 158431 49989
rect 169539 50147 169567 50175
rect 169601 50147 169629 50175
rect 169539 50085 169567 50113
rect 169601 50085 169629 50113
rect 169539 50023 169567 50051
rect 169601 50023 169629 50051
rect 169539 49961 169567 49989
rect 169601 49961 169629 49989
rect 161859 47147 161887 47175
rect 161921 47147 161949 47175
rect 161859 47085 161887 47113
rect 161921 47085 161949 47113
rect 161859 47023 161887 47051
rect 161921 47023 161949 47051
rect 161859 46961 161887 46989
rect 161921 46961 161949 46989
rect 171717 47147 171745 47175
rect 171779 47147 171807 47175
rect 171841 47147 171869 47175
rect 171903 47147 171931 47175
rect 171717 47085 171745 47113
rect 171779 47085 171807 47113
rect 171841 47085 171869 47113
rect 171903 47085 171931 47113
rect 171717 47023 171745 47051
rect 171779 47023 171807 47051
rect 171841 47023 171869 47051
rect 171903 47023 171931 47051
rect 171717 46961 171745 46989
rect 171779 46961 171807 46989
rect 171841 46961 171869 46989
rect 171903 46961 171931 46989
rect 158217 41147 158245 41175
rect 158279 41147 158307 41175
rect 158341 41147 158369 41175
rect 158403 41147 158431 41175
rect 158217 41085 158245 41113
rect 158279 41085 158307 41113
rect 158341 41085 158369 41113
rect 158403 41085 158431 41113
rect 158217 41023 158245 41051
rect 158279 41023 158307 41051
rect 158341 41023 158369 41051
rect 158403 41023 158431 41051
rect 158217 40961 158245 40989
rect 158279 40961 158307 40989
rect 158341 40961 158369 40989
rect 158403 40961 158431 40989
rect 169539 41147 169567 41175
rect 169601 41147 169629 41175
rect 169539 41085 169567 41113
rect 169601 41085 169629 41113
rect 169539 41023 169567 41051
rect 169601 41023 169629 41051
rect 169539 40961 169567 40989
rect 169601 40961 169629 40989
rect 161859 38147 161887 38175
rect 161921 38147 161949 38175
rect 161859 38085 161887 38113
rect 161921 38085 161949 38113
rect 161859 38023 161887 38051
rect 161921 38023 161949 38051
rect 161859 37961 161887 37989
rect 161921 37961 161949 37989
rect 171717 38147 171745 38175
rect 171779 38147 171807 38175
rect 171841 38147 171869 38175
rect 171903 38147 171931 38175
rect 171717 38085 171745 38113
rect 171779 38085 171807 38113
rect 171841 38085 171869 38113
rect 171903 38085 171931 38113
rect 171717 38023 171745 38051
rect 171779 38023 171807 38051
rect 171841 38023 171869 38051
rect 171903 38023 171931 38051
rect 171717 37961 171745 37989
rect 171779 37961 171807 37989
rect 171841 37961 171869 37989
rect 171903 37961 171931 37989
rect 158217 32147 158245 32175
rect 158279 32147 158307 32175
rect 158341 32147 158369 32175
rect 158403 32147 158431 32175
rect 158217 32085 158245 32113
rect 158279 32085 158307 32113
rect 158341 32085 158369 32113
rect 158403 32085 158431 32113
rect 158217 32023 158245 32051
rect 158279 32023 158307 32051
rect 158341 32023 158369 32051
rect 158403 32023 158431 32051
rect 158217 31961 158245 31989
rect 158279 31961 158307 31989
rect 158341 31961 158369 31989
rect 158403 31961 158431 31989
rect 169539 32147 169567 32175
rect 169601 32147 169629 32175
rect 169539 32085 169567 32113
rect 169601 32085 169629 32113
rect 169539 32023 169567 32051
rect 169601 32023 169629 32051
rect 169539 31961 169567 31989
rect 169601 31961 169629 31989
rect 161859 29147 161887 29175
rect 161921 29147 161949 29175
rect 161859 29085 161887 29113
rect 161921 29085 161949 29113
rect 161859 29023 161887 29051
rect 161921 29023 161949 29051
rect 161859 28961 161887 28989
rect 161921 28961 161949 28989
rect 171717 29147 171745 29175
rect 171779 29147 171807 29175
rect 171841 29147 171869 29175
rect 171903 29147 171931 29175
rect 171717 29085 171745 29113
rect 171779 29085 171807 29113
rect 171841 29085 171869 29113
rect 171903 29085 171931 29113
rect 171717 29023 171745 29051
rect 171779 29023 171807 29051
rect 171841 29023 171869 29051
rect 171903 29023 171931 29051
rect 171717 28961 171745 28989
rect 171779 28961 171807 28989
rect 171841 28961 171869 28989
rect 171903 28961 171931 28989
rect 158217 23147 158245 23175
rect 158279 23147 158307 23175
rect 158341 23147 158369 23175
rect 158403 23147 158431 23175
rect 158217 23085 158245 23113
rect 158279 23085 158307 23113
rect 158341 23085 158369 23113
rect 158403 23085 158431 23113
rect 158217 23023 158245 23051
rect 158279 23023 158307 23051
rect 158341 23023 158369 23051
rect 158403 23023 158431 23051
rect 158217 22961 158245 22989
rect 158279 22961 158307 22989
rect 158341 22961 158369 22989
rect 158403 22961 158431 22989
rect 169539 23147 169567 23175
rect 169601 23147 169629 23175
rect 169539 23085 169567 23113
rect 169601 23085 169629 23113
rect 169539 23023 169567 23051
rect 169601 23023 169629 23051
rect 169539 22961 169567 22989
rect 169601 22961 169629 22989
rect 161859 20147 161887 20175
rect 161921 20147 161949 20175
rect 161859 20085 161887 20113
rect 161921 20085 161949 20113
rect 161859 20023 161887 20051
rect 161921 20023 161949 20051
rect 161859 19961 161887 19989
rect 161921 19961 161949 19989
rect 171717 20147 171745 20175
rect 171779 20147 171807 20175
rect 171841 20147 171869 20175
rect 171903 20147 171931 20175
rect 171717 20085 171745 20113
rect 171779 20085 171807 20113
rect 171841 20085 171869 20113
rect 171903 20085 171931 20113
rect 171717 20023 171745 20051
rect 171779 20023 171807 20051
rect 171841 20023 171869 20051
rect 171903 20023 171931 20051
rect 171717 19961 171745 19989
rect 171779 19961 171807 19989
rect 171841 19961 171869 19989
rect 171903 19961 171931 19989
rect 158217 14147 158245 14175
rect 158279 14147 158307 14175
rect 158341 14147 158369 14175
rect 158403 14147 158431 14175
rect 158217 14085 158245 14113
rect 158279 14085 158307 14113
rect 158341 14085 158369 14113
rect 158403 14085 158431 14113
rect 158217 14023 158245 14051
rect 158279 14023 158307 14051
rect 158341 14023 158369 14051
rect 158403 14023 158431 14051
rect 158217 13961 158245 13989
rect 158279 13961 158307 13989
rect 158341 13961 158369 13989
rect 158403 13961 158431 13989
rect 169539 14147 169567 14175
rect 169601 14147 169629 14175
rect 169539 14085 169567 14113
rect 169601 14085 169629 14113
rect 169539 14023 169567 14051
rect 169601 14023 169629 14051
rect 169539 13961 169567 13989
rect 169601 13961 169629 13989
rect 161859 11147 161887 11175
rect 161921 11147 161949 11175
rect 161859 11085 161887 11113
rect 161921 11085 161949 11113
rect 161859 11023 161887 11051
rect 161921 11023 161949 11051
rect 161859 10961 161887 10989
rect 161921 10961 161949 10989
rect 171717 11147 171745 11175
rect 171779 11147 171807 11175
rect 171841 11147 171869 11175
rect 171903 11147 171931 11175
rect 171717 11085 171745 11113
rect 171779 11085 171807 11113
rect 171841 11085 171869 11113
rect 171903 11085 171931 11113
rect 171717 11023 171745 11051
rect 171779 11023 171807 11051
rect 171841 11023 171869 11051
rect 171903 11023 171931 11051
rect 171717 10961 171745 10989
rect 171779 10961 171807 10989
rect 171841 10961 171869 10989
rect 171903 10961 171931 10989
rect 158217 5147 158245 5175
rect 158279 5147 158307 5175
rect 158341 5147 158369 5175
rect 158403 5147 158431 5175
rect 158217 5085 158245 5113
rect 158279 5085 158307 5113
rect 158341 5085 158369 5113
rect 158403 5085 158431 5113
rect 158217 5023 158245 5051
rect 158279 5023 158307 5051
rect 158341 5023 158369 5051
rect 158403 5023 158431 5051
rect 158217 4961 158245 4989
rect 158279 4961 158307 4989
rect 158341 4961 158369 4989
rect 158403 4961 158431 4989
rect 169539 5147 169567 5175
rect 169601 5147 169629 5175
rect 169539 5085 169567 5113
rect 169601 5085 169629 5113
rect 169539 5023 169567 5051
rect 169601 5023 169629 5051
rect 169539 4961 169567 4989
rect 169601 4961 169629 4989
rect 158217 -588 158245 -560
rect 158279 -588 158307 -560
rect 158341 -588 158369 -560
rect 158403 -588 158431 -560
rect 158217 -650 158245 -622
rect 158279 -650 158307 -622
rect 158341 -650 158369 -622
rect 158403 -650 158431 -622
rect 158217 -712 158245 -684
rect 158279 -712 158307 -684
rect 158341 -712 158369 -684
rect 158403 -712 158431 -684
rect 158217 -774 158245 -746
rect 158279 -774 158307 -746
rect 158341 -774 158369 -746
rect 158403 -774 158431 -746
rect 171717 2147 171745 2175
rect 171779 2147 171807 2175
rect 171841 2147 171869 2175
rect 171903 2147 171931 2175
rect 171717 2085 171745 2113
rect 171779 2085 171807 2113
rect 171841 2085 171869 2113
rect 171903 2085 171931 2113
rect 171717 2023 171745 2051
rect 171779 2023 171807 2051
rect 171841 2023 171869 2051
rect 171903 2023 171931 2051
rect 171717 1961 171745 1989
rect 171779 1961 171807 1989
rect 171841 1961 171869 1989
rect 171903 1961 171931 1989
rect 171717 -108 171745 -80
rect 171779 -108 171807 -80
rect 171841 -108 171869 -80
rect 171903 -108 171931 -80
rect 171717 -170 171745 -142
rect 171779 -170 171807 -142
rect 171841 -170 171869 -142
rect 171903 -170 171931 -142
rect 171717 -232 171745 -204
rect 171779 -232 171807 -204
rect 171841 -232 171869 -204
rect 171903 -232 171931 -204
rect 171717 -294 171745 -266
rect 171779 -294 171807 -266
rect 171841 -294 171869 -266
rect 171903 -294 171931 -266
rect 173577 299058 173605 299086
rect 173639 299058 173667 299086
rect 173701 299058 173729 299086
rect 173763 299058 173791 299086
rect 173577 298996 173605 299024
rect 173639 298996 173667 299024
rect 173701 298996 173729 299024
rect 173763 298996 173791 299024
rect 173577 298934 173605 298962
rect 173639 298934 173667 298962
rect 173701 298934 173729 298962
rect 173763 298934 173791 298962
rect 173577 298872 173605 298900
rect 173639 298872 173667 298900
rect 173701 298872 173729 298900
rect 173763 298872 173791 298900
rect 173577 293147 173605 293175
rect 173639 293147 173667 293175
rect 173701 293147 173729 293175
rect 173763 293147 173791 293175
rect 173577 293085 173605 293113
rect 173639 293085 173667 293113
rect 173701 293085 173729 293113
rect 173763 293085 173791 293113
rect 173577 293023 173605 293051
rect 173639 293023 173667 293051
rect 173701 293023 173729 293051
rect 173763 293023 173791 293051
rect 173577 292961 173605 292989
rect 173639 292961 173667 292989
rect 173701 292961 173729 292989
rect 173763 292961 173791 292989
rect 173577 284147 173605 284175
rect 173639 284147 173667 284175
rect 173701 284147 173729 284175
rect 173763 284147 173791 284175
rect 173577 284085 173605 284113
rect 173639 284085 173667 284113
rect 173701 284085 173729 284113
rect 173763 284085 173791 284113
rect 173577 284023 173605 284051
rect 173639 284023 173667 284051
rect 173701 284023 173729 284051
rect 173763 284023 173791 284051
rect 173577 283961 173605 283989
rect 173639 283961 173667 283989
rect 173701 283961 173729 283989
rect 173763 283961 173791 283989
rect 173577 275147 173605 275175
rect 173639 275147 173667 275175
rect 173701 275147 173729 275175
rect 173763 275147 173791 275175
rect 173577 275085 173605 275113
rect 173639 275085 173667 275113
rect 173701 275085 173729 275113
rect 173763 275085 173791 275113
rect 173577 275023 173605 275051
rect 173639 275023 173667 275051
rect 173701 275023 173729 275051
rect 173763 275023 173791 275051
rect 173577 274961 173605 274989
rect 173639 274961 173667 274989
rect 173701 274961 173729 274989
rect 173763 274961 173791 274989
rect 173577 266147 173605 266175
rect 173639 266147 173667 266175
rect 173701 266147 173729 266175
rect 173763 266147 173791 266175
rect 173577 266085 173605 266113
rect 173639 266085 173667 266113
rect 173701 266085 173729 266113
rect 173763 266085 173791 266113
rect 173577 266023 173605 266051
rect 173639 266023 173667 266051
rect 173701 266023 173729 266051
rect 173763 266023 173791 266051
rect 173577 265961 173605 265989
rect 173639 265961 173667 265989
rect 173701 265961 173729 265989
rect 173763 265961 173791 265989
rect 173577 257147 173605 257175
rect 173639 257147 173667 257175
rect 173701 257147 173729 257175
rect 173763 257147 173791 257175
rect 173577 257085 173605 257113
rect 173639 257085 173667 257113
rect 173701 257085 173729 257113
rect 173763 257085 173791 257113
rect 173577 257023 173605 257051
rect 173639 257023 173667 257051
rect 173701 257023 173729 257051
rect 173763 257023 173791 257051
rect 173577 256961 173605 256989
rect 173639 256961 173667 256989
rect 173701 256961 173729 256989
rect 173763 256961 173791 256989
rect 173577 248147 173605 248175
rect 173639 248147 173667 248175
rect 173701 248147 173729 248175
rect 173763 248147 173791 248175
rect 173577 248085 173605 248113
rect 173639 248085 173667 248113
rect 173701 248085 173729 248113
rect 173763 248085 173791 248113
rect 173577 248023 173605 248051
rect 173639 248023 173667 248051
rect 173701 248023 173729 248051
rect 173763 248023 173791 248051
rect 173577 247961 173605 247989
rect 173639 247961 173667 247989
rect 173701 247961 173729 247989
rect 173763 247961 173791 247989
rect 173577 239147 173605 239175
rect 173639 239147 173667 239175
rect 173701 239147 173729 239175
rect 173763 239147 173791 239175
rect 173577 239085 173605 239113
rect 173639 239085 173667 239113
rect 173701 239085 173729 239113
rect 173763 239085 173791 239113
rect 173577 239023 173605 239051
rect 173639 239023 173667 239051
rect 173701 239023 173729 239051
rect 173763 239023 173791 239051
rect 173577 238961 173605 238989
rect 173639 238961 173667 238989
rect 173701 238961 173729 238989
rect 173763 238961 173791 238989
rect 173577 230147 173605 230175
rect 173639 230147 173667 230175
rect 173701 230147 173729 230175
rect 173763 230147 173791 230175
rect 173577 230085 173605 230113
rect 173639 230085 173667 230113
rect 173701 230085 173729 230113
rect 173763 230085 173791 230113
rect 173577 230023 173605 230051
rect 173639 230023 173667 230051
rect 173701 230023 173729 230051
rect 173763 230023 173791 230051
rect 173577 229961 173605 229989
rect 173639 229961 173667 229989
rect 173701 229961 173729 229989
rect 173763 229961 173791 229989
rect 173577 221147 173605 221175
rect 173639 221147 173667 221175
rect 173701 221147 173729 221175
rect 173763 221147 173791 221175
rect 173577 221085 173605 221113
rect 173639 221085 173667 221113
rect 173701 221085 173729 221113
rect 173763 221085 173791 221113
rect 173577 221023 173605 221051
rect 173639 221023 173667 221051
rect 173701 221023 173729 221051
rect 173763 221023 173791 221051
rect 173577 220961 173605 220989
rect 173639 220961 173667 220989
rect 173701 220961 173729 220989
rect 173763 220961 173791 220989
rect 173577 212147 173605 212175
rect 173639 212147 173667 212175
rect 173701 212147 173729 212175
rect 173763 212147 173791 212175
rect 173577 212085 173605 212113
rect 173639 212085 173667 212113
rect 173701 212085 173729 212113
rect 173763 212085 173791 212113
rect 173577 212023 173605 212051
rect 173639 212023 173667 212051
rect 173701 212023 173729 212051
rect 173763 212023 173791 212051
rect 173577 211961 173605 211989
rect 173639 211961 173667 211989
rect 173701 211961 173729 211989
rect 173763 211961 173791 211989
rect 173577 203147 173605 203175
rect 173639 203147 173667 203175
rect 173701 203147 173729 203175
rect 173763 203147 173791 203175
rect 173577 203085 173605 203113
rect 173639 203085 173667 203113
rect 173701 203085 173729 203113
rect 173763 203085 173791 203113
rect 173577 203023 173605 203051
rect 173639 203023 173667 203051
rect 173701 203023 173729 203051
rect 173763 203023 173791 203051
rect 173577 202961 173605 202989
rect 173639 202961 173667 202989
rect 173701 202961 173729 202989
rect 173763 202961 173791 202989
rect 173577 194147 173605 194175
rect 173639 194147 173667 194175
rect 173701 194147 173729 194175
rect 173763 194147 173791 194175
rect 173577 194085 173605 194113
rect 173639 194085 173667 194113
rect 173701 194085 173729 194113
rect 173763 194085 173791 194113
rect 173577 194023 173605 194051
rect 173639 194023 173667 194051
rect 173701 194023 173729 194051
rect 173763 194023 173791 194051
rect 173577 193961 173605 193989
rect 173639 193961 173667 193989
rect 173701 193961 173729 193989
rect 173763 193961 173791 193989
rect 173577 185147 173605 185175
rect 173639 185147 173667 185175
rect 173701 185147 173729 185175
rect 173763 185147 173791 185175
rect 173577 185085 173605 185113
rect 173639 185085 173667 185113
rect 173701 185085 173729 185113
rect 173763 185085 173791 185113
rect 173577 185023 173605 185051
rect 173639 185023 173667 185051
rect 173701 185023 173729 185051
rect 173763 185023 173791 185051
rect 173577 184961 173605 184989
rect 173639 184961 173667 184989
rect 173701 184961 173729 184989
rect 173763 184961 173791 184989
rect 173577 176147 173605 176175
rect 173639 176147 173667 176175
rect 173701 176147 173729 176175
rect 173763 176147 173791 176175
rect 173577 176085 173605 176113
rect 173639 176085 173667 176113
rect 173701 176085 173729 176113
rect 173763 176085 173791 176113
rect 173577 176023 173605 176051
rect 173639 176023 173667 176051
rect 173701 176023 173729 176051
rect 173763 176023 173791 176051
rect 173577 175961 173605 175989
rect 173639 175961 173667 175989
rect 173701 175961 173729 175989
rect 173763 175961 173791 175989
rect 187077 298578 187105 298606
rect 187139 298578 187167 298606
rect 187201 298578 187229 298606
rect 187263 298578 187291 298606
rect 187077 298516 187105 298544
rect 187139 298516 187167 298544
rect 187201 298516 187229 298544
rect 187263 298516 187291 298544
rect 187077 298454 187105 298482
rect 187139 298454 187167 298482
rect 187201 298454 187229 298482
rect 187263 298454 187291 298482
rect 187077 298392 187105 298420
rect 187139 298392 187167 298420
rect 187201 298392 187229 298420
rect 187263 298392 187291 298420
rect 187077 290147 187105 290175
rect 187139 290147 187167 290175
rect 187201 290147 187229 290175
rect 187263 290147 187291 290175
rect 187077 290085 187105 290113
rect 187139 290085 187167 290113
rect 187201 290085 187229 290113
rect 187263 290085 187291 290113
rect 187077 290023 187105 290051
rect 187139 290023 187167 290051
rect 187201 290023 187229 290051
rect 187263 290023 187291 290051
rect 187077 289961 187105 289989
rect 187139 289961 187167 289989
rect 187201 289961 187229 289989
rect 187263 289961 187291 289989
rect 187077 281147 187105 281175
rect 187139 281147 187167 281175
rect 187201 281147 187229 281175
rect 187263 281147 187291 281175
rect 187077 281085 187105 281113
rect 187139 281085 187167 281113
rect 187201 281085 187229 281113
rect 187263 281085 187291 281113
rect 187077 281023 187105 281051
rect 187139 281023 187167 281051
rect 187201 281023 187229 281051
rect 187263 281023 187291 281051
rect 187077 280961 187105 280989
rect 187139 280961 187167 280989
rect 187201 280961 187229 280989
rect 187263 280961 187291 280989
rect 187077 272147 187105 272175
rect 187139 272147 187167 272175
rect 187201 272147 187229 272175
rect 187263 272147 187291 272175
rect 187077 272085 187105 272113
rect 187139 272085 187167 272113
rect 187201 272085 187229 272113
rect 187263 272085 187291 272113
rect 187077 272023 187105 272051
rect 187139 272023 187167 272051
rect 187201 272023 187229 272051
rect 187263 272023 187291 272051
rect 187077 271961 187105 271989
rect 187139 271961 187167 271989
rect 187201 271961 187229 271989
rect 187263 271961 187291 271989
rect 187077 263147 187105 263175
rect 187139 263147 187167 263175
rect 187201 263147 187229 263175
rect 187263 263147 187291 263175
rect 187077 263085 187105 263113
rect 187139 263085 187167 263113
rect 187201 263085 187229 263113
rect 187263 263085 187291 263113
rect 187077 263023 187105 263051
rect 187139 263023 187167 263051
rect 187201 263023 187229 263051
rect 187263 263023 187291 263051
rect 187077 262961 187105 262989
rect 187139 262961 187167 262989
rect 187201 262961 187229 262989
rect 187263 262961 187291 262989
rect 187077 254147 187105 254175
rect 187139 254147 187167 254175
rect 187201 254147 187229 254175
rect 187263 254147 187291 254175
rect 187077 254085 187105 254113
rect 187139 254085 187167 254113
rect 187201 254085 187229 254113
rect 187263 254085 187291 254113
rect 187077 254023 187105 254051
rect 187139 254023 187167 254051
rect 187201 254023 187229 254051
rect 187263 254023 187291 254051
rect 187077 253961 187105 253989
rect 187139 253961 187167 253989
rect 187201 253961 187229 253989
rect 187263 253961 187291 253989
rect 187077 245147 187105 245175
rect 187139 245147 187167 245175
rect 187201 245147 187229 245175
rect 187263 245147 187291 245175
rect 187077 245085 187105 245113
rect 187139 245085 187167 245113
rect 187201 245085 187229 245113
rect 187263 245085 187291 245113
rect 187077 245023 187105 245051
rect 187139 245023 187167 245051
rect 187201 245023 187229 245051
rect 187263 245023 187291 245051
rect 187077 244961 187105 244989
rect 187139 244961 187167 244989
rect 187201 244961 187229 244989
rect 187263 244961 187291 244989
rect 187077 236147 187105 236175
rect 187139 236147 187167 236175
rect 187201 236147 187229 236175
rect 187263 236147 187291 236175
rect 187077 236085 187105 236113
rect 187139 236085 187167 236113
rect 187201 236085 187229 236113
rect 187263 236085 187291 236113
rect 187077 236023 187105 236051
rect 187139 236023 187167 236051
rect 187201 236023 187229 236051
rect 187263 236023 187291 236051
rect 187077 235961 187105 235989
rect 187139 235961 187167 235989
rect 187201 235961 187229 235989
rect 187263 235961 187291 235989
rect 187077 227147 187105 227175
rect 187139 227147 187167 227175
rect 187201 227147 187229 227175
rect 187263 227147 187291 227175
rect 187077 227085 187105 227113
rect 187139 227085 187167 227113
rect 187201 227085 187229 227113
rect 187263 227085 187291 227113
rect 187077 227023 187105 227051
rect 187139 227023 187167 227051
rect 187201 227023 187229 227051
rect 187263 227023 187291 227051
rect 187077 226961 187105 226989
rect 187139 226961 187167 226989
rect 187201 226961 187229 226989
rect 187263 226961 187291 226989
rect 187077 218147 187105 218175
rect 187139 218147 187167 218175
rect 187201 218147 187229 218175
rect 187263 218147 187291 218175
rect 187077 218085 187105 218113
rect 187139 218085 187167 218113
rect 187201 218085 187229 218113
rect 187263 218085 187291 218113
rect 187077 218023 187105 218051
rect 187139 218023 187167 218051
rect 187201 218023 187229 218051
rect 187263 218023 187291 218051
rect 187077 217961 187105 217989
rect 187139 217961 187167 217989
rect 187201 217961 187229 217989
rect 187263 217961 187291 217989
rect 187077 209147 187105 209175
rect 187139 209147 187167 209175
rect 187201 209147 187229 209175
rect 187263 209147 187291 209175
rect 187077 209085 187105 209113
rect 187139 209085 187167 209113
rect 187201 209085 187229 209113
rect 187263 209085 187291 209113
rect 187077 209023 187105 209051
rect 187139 209023 187167 209051
rect 187201 209023 187229 209051
rect 187263 209023 187291 209051
rect 187077 208961 187105 208989
rect 187139 208961 187167 208989
rect 187201 208961 187229 208989
rect 187263 208961 187291 208989
rect 187077 200147 187105 200175
rect 187139 200147 187167 200175
rect 187201 200147 187229 200175
rect 187263 200147 187291 200175
rect 187077 200085 187105 200113
rect 187139 200085 187167 200113
rect 187201 200085 187229 200113
rect 187263 200085 187291 200113
rect 187077 200023 187105 200051
rect 187139 200023 187167 200051
rect 187201 200023 187229 200051
rect 187263 200023 187291 200051
rect 187077 199961 187105 199989
rect 187139 199961 187167 199989
rect 187201 199961 187229 199989
rect 187263 199961 187291 199989
rect 187077 191147 187105 191175
rect 187139 191147 187167 191175
rect 187201 191147 187229 191175
rect 187263 191147 187291 191175
rect 187077 191085 187105 191113
rect 187139 191085 187167 191113
rect 187201 191085 187229 191113
rect 187263 191085 187291 191113
rect 187077 191023 187105 191051
rect 187139 191023 187167 191051
rect 187201 191023 187229 191051
rect 187263 191023 187291 191051
rect 187077 190961 187105 190989
rect 187139 190961 187167 190989
rect 187201 190961 187229 190989
rect 187263 190961 187291 190989
rect 187077 182147 187105 182175
rect 187139 182147 187167 182175
rect 187201 182147 187229 182175
rect 187263 182147 187291 182175
rect 187077 182085 187105 182113
rect 187139 182085 187167 182113
rect 187201 182085 187229 182113
rect 187263 182085 187291 182113
rect 187077 182023 187105 182051
rect 187139 182023 187167 182051
rect 187201 182023 187229 182051
rect 187263 182023 187291 182051
rect 187077 181961 187105 181989
rect 187139 181961 187167 181989
rect 187201 181961 187229 181989
rect 187263 181961 187291 181989
rect 177219 173147 177247 173175
rect 177281 173147 177309 173175
rect 177219 173085 177247 173113
rect 177281 173085 177309 173113
rect 177219 173023 177247 173051
rect 177281 173023 177309 173051
rect 177219 172961 177247 172989
rect 177281 172961 177309 172989
rect 187077 173147 187105 173175
rect 187139 173147 187167 173175
rect 187201 173147 187229 173175
rect 187263 173147 187291 173175
rect 187077 173085 187105 173113
rect 187139 173085 187167 173113
rect 187201 173085 187229 173113
rect 187263 173085 187291 173113
rect 187077 173023 187105 173051
rect 187139 173023 187167 173051
rect 187201 173023 187229 173051
rect 187263 173023 187291 173051
rect 187077 172961 187105 172989
rect 187139 172961 187167 172989
rect 187201 172961 187229 172989
rect 187263 172961 187291 172989
rect 173577 167147 173605 167175
rect 173639 167147 173667 167175
rect 173701 167147 173729 167175
rect 173763 167147 173791 167175
rect 173577 167085 173605 167113
rect 173639 167085 173667 167113
rect 173701 167085 173729 167113
rect 173763 167085 173791 167113
rect 173577 167023 173605 167051
rect 173639 167023 173667 167051
rect 173701 167023 173729 167051
rect 173763 167023 173791 167051
rect 173577 166961 173605 166989
rect 173639 166961 173667 166989
rect 173701 166961 173729 166989
rect 173763 166961 173791 166989
rect 184899 167147 184927 167175
rect 184961 167147 184989 167175
rect 184899 167085 184927 167113
rect 184961 167085 184989 167113
rect 184899 167023 184927 167051
rect 184961 167023 184989 167051
rect 184899 166961 184927 166989
rect 184961 166961 184989 166989
rect 177219 164147 177247 164175
rect 177281 164147 177309 164175
rect 177219 164085 177247 164113
rect 177281 164085 177309 164113
rect 177219 164023 177247 164051
rect 177281 164023 177309 164051
rect 177219 163961 177247 163989
rect 177281 163961 177309 163989
rect 187077 164147 187105 164175
rect 187139 164147 187167 164175
rect 187201 164147 187229 164175
rect 187263 164147 187291 164175
rect 187077 164085 187105 164113
rect 187139 164085 187167 164113
rect 187201 164085 187229 164113
rect 187263 164085 187291 164113
rect 187077 164023 187105 164051
rect 187139 164023 187167 164051
rect 187201 164023 187229 164051
rect 187263 164023 187291 164051
rect 187077 163961 187105 163989
rect 187139 163961 187167 163989
rect 187201 163961 187229 163989
rect 187263 163961 187291 163989
rect 173577 158147 173605 158175
rect 173639 158147 173667 158175
rect 173701 158147 173729 158175
rect 173763 158147 173791 158175
rect 173577 158085 173605 158113
rect 173639 158085 173667 158113
rect 173701 158085 173729 158113
rect 173763 158085 173791 158113
rect 173577 158023 173605 158051
rect 173639 158023 173667 158051
rect 173701 158023 173729 158051
rect 173763 158023 173791 158051
rect 173577 157961 173605 157989
rect 173639 157961 173667 157989
rect 173701 157961 173729 157989
rect 173763 157961 173791 157989
rect 184899 158147 184927 158175
rect 184961 158147 184989 158175
rect 184899 158085 184927 158113
rect 184961 158085 184989 158113
rect 184899 158023 184927 158051
rect 184961 158023 184989 158051
rect 184899 157961 184927 157989
rect 184961 157961 184989 157989
rect 177219 155147 177247 155175
rect 177281 155147 177309 155175
rect 177219 155085 177247 155113
rect 177281 155085 177309 155113
rect 177219 155023 177247 155051
rect 177281 155023 177309 155051
rect 177219 154961 177247 154989
rect 177281 154961 177309 154989
rect 187077 155147 187105 155175
rect 187139 155147 187167 155175
rect 187201 155147 187229 155175
rect 187263 155147 187291 155175
rect 187077 155085 187105 155113
rect 187139 155085 187167 155113
rect 187201 155085 187229 155113
rect 187263 155085 187291 155113
rect 187077 155023 187105 155051
rect 187139 155023 187167 155051
rect 187201 155023 187229 155051
rect 187263 155023 187291 155051
rect 187077 154961 187105 154989
rect 187139 154961 187167 154989
rect 187201 154961 187229 154989
rect 187263 154961 187291 154989
rect 173577 149147 173605 149175
rect 173639 149147 173667 149175
rect 173701 149147 173729 149175
rect 173763 149147 173791 149175
rect 173577 149085 173605 149113
rect 173639 149085 173667 149113
rect 173701 149085 173729 149113
rect 173763 149085 173791 149113
rect 173577 149023 173605 149051
rect 173639 149023 173667 149051
rect 173701 149023 173729 149051
rect 173763 149023 173791 149051
rect 173577 148961 173605 148989
rect 173639 148961 173667 148989
rect 173701 148961 173729 148989
rect 173763 148961 173791 148989
rect 184899 149147 184927 149175
rect 184961 149147 184989 149175
rect 184899 149085 184927 149113
rect 184961 149085 184989 149113
rect 184899 149023 184927 149051
rect 184961 149023 184989 149051
rect 184899 148961 184927 148989
rect 184961 148961 184989 148989
rect 177219 146147 177247 146175
rect 177281 146147 177309 146175
rect 177219 146085 177247 146113
rect 177281 146085 177309 146113
rect 177219 146023 177247 146051
rect 177281 146023 177309 146051
rect 177219 145961 177247 145989
rect 177281 145961 177309 145989
rect 187077 146147 187105 146175
rect 187139 146147 187167 146175
rect 187201 146147 187229 146175
rect 187263 146147 187291 146175
rect 187077 146085 187105 146113
rect 187139 146085 187167 146113
rect 187201 146085 187229 146113
rect 187263 146085 187291 146113
rect 187077 146023 187105 146051
rect 187139 146023 187167 146051
rect 187201 146023 187229 146051
rect 187263 146023 187291 146051
rect 187077 145961 187105 145989
rect 187139 145961 187167 145989
rect 187201 145961 187229 145989
rect 187263 145961 187291 145989
rect 173577 140147 173605 140175
rect 173639 140147 173667 140175
rect 173701 140147 173729 140175
rect 173763 140147 173791 140175
rect 173577 140085 173605 140113
rect 173639 140085 173667 140113
rect 173701 140085 173729 140113
rect 173763 140085 173791 140113
rect 173577 140023 173605 140051
rect 173639 140023 173667 140051
rect 173701 140023 173729 140051
rect 173763 140023 173791 140051
rect 173577 139961 173605 139989
rect 173639 139961 173667 139989
rect 173701 139961 173729 139989
rect 173763 139961 173791 139989
rect 184899 140147 184927 140175
rect 184961 140147 184989 140175
rect 184899 140085 184927 140113
rect 184961 140085 184989 140113
rect 184899 140023 184927 140051
rect 184961 140023 184989 140051
rect 184899 139961 184927 139989
rect 184961 139961 184989 139989
rect 177219 137147 177247 137175
rect 177281 137147 177309 137175
rect 177219 137085 177247 137113
rect 177281 137085 177309 137113
rect 177219 137023 177247 137051
rect 177281 137023 177309 137051
rect 177219 136961 177247 136989
rect 177281 136961 177309 136989
rect 187077 137147 187105 137175
rect 187139 137147 187167 137175
rect 187201 137147 187229 137175
rect 187263 137147 187291 137175
rect 187077 137085 187105 137113
rect 187139 137085 187167 137113
rect 187201 137085 187229 137113
rect 187263 137085 187291 137113
rect 187077 137023 187105 137051
rect 187139 137023 187167 137051
rect 187201 137023 187229 137051
rect 187263 137023 187291 137051
rect 187077 136961 187105 136989
rect 187139 136961 187167 136989
rect 187201 136961 187229 136989
rect 187263 136961 187291 136989
rect 173577 131147 173605 131175
rect 173639 131147 173667 131175
rect 173701 131147 173729 131175
rect 173763 131147 173791 131175
rect 173577 131085 173605 131113
rect 173639 131085 173667 131113
rect 173701 131085 173729 131113
rect 173763 131085 173791 131113
rect 173577 131023 173605 131051
rect 173639 131023 173667 131051
rect 173701 131023 173729 131051
rect 173763 131023 173791 131051
rect 173577 130961 173605 130989
rect 173639 130961 173667 130989
rect 173701 130961 173729 130989
rect 173763 130961 173791 130989
rect 184899 131147 184927 131175
rect 184961 131147 184989 131175
rect 184899 131085 184927 131113
rect 184961 131085 184989 131113
rect 184899 131023 184927 131051
rect 184961 131023 184989 131051
rect 184899 130961 184927 130989
rect 184961 130961 184989 130989
rect 177219 128147 177247 128175
rect 177281 128147 177309 128175
rect 177219 128085 177247 128113
rect 177281 128085 177309 128113
rect 177219 128023 177247 128051
rect 177281 128023 177309 128051
rect 177219 127961 177247 127989
rect 177281 127961 177309 127989
rect 187077 128147 187105 128175
rect 187139 128147 187167 128175
rect 187201 128147 187229 128175
rect 187263 128147 187291 128175
rect 187077 128085 187105 128113
rect 187139 128085 187167 128113
rect 187201 128085 187229 128113
rect 187263 128085 187291 128113
rect 187077 128023 187105 128051
rect 187139 128023 187167 128051
rect 187201 128023 187229 128051
rect 187263 128023 187291 128051
rect 187077 127961 187105 127989
rect 187139 127961 187167 127989
rect 187201 127961 187229 127989
rect 187263 127961 187291 127989
rect 173577 122147 173605 122175
rect 173639 122147 173667 122175
rect 173701 122147 173729 122175
rect 173763 122147 173791 122175
rect 173577 122085 173605 122113
rect 173639 122085 173667 122113
rect 173701 122085 173729 122113
rect 173763 122085 173791 122113
rect 173577 122023 173605 122051
rect 173639 122023 173667 122051
rect 173701 122023 173729 122051
rect 173763 122023 173791 122051
rect 173577 121961 173605 121989
rect 173639 121961 173667 121989
rect 173701 121961 173729 121989
rect 173763 121961 173791 121989
rect 184899 122147 184927 122175
rect 184961 122147 184989 122175
rect 184899 122085 184927 122113
rect 184961 122085 184989 122113
rect 184899 122023 184927 122051
rect 184961 122023 184989 122051
rect 184899 121961 184927 121989
rect 184961 121961 184989 121989
rect 177219 119147 177247 119175
rect 177281 119147 177309 119175
rect 177219 119085 177247 119113
rect 177281 119085 177309 119113
rect 177219 119023 177247 119051
rect 177281 119023 177309 119051
rect 177219 118961 177247 118989
rect 177281 118961 177309 118989
rect 187077 119147 187105 119175
rect 187139 119147 187167 119175
rect 187201 119147 187229 119175
rect 187263 119147 187291 119175
rect 187077 119085 187105 119113
rect 187139 119085 187167 119113
rect 187201 119085 187229 119113
rect 187263 119085 187291 119113
rect 187077 119023 187105 119051
rect 187139 119023 187167 119051
rect 187201 119023 187229 119051
rect 187263 119023 187291 119051
rect 187077 118961 187105 118989
rect 187139 118961 187167 118989
rect 187201 118961 187229 118989
rect 187263 118961 187291 118989
rect 173577 113147 173605 113175
rect 173639 113147 173667 113175
rect 173701 113147 173729 113175
rect 173763 113147 173791 113175
rect 173577 113085 173605 113113
rect 173639 113085 173667 113113
rect 173701 113085 173729 113113
rect 173763 113085 173791 113113
rect 173577 113023 173605 113051
rect 173639 113023 173667 113051
rect 173701 113023 173729 113051
rect 173763 113023 173791 113051
rect 173577 112961 173605 112989
rect 173639 112961 173667 112989
rect 173701 112961 173729 112989
rect 173763 112961 173791 112989
rect 184899 113147 184927 113175
rect 184961 113147 184989 113175
rect 184899 113085 184927 113113
rect 184961 113085 184989 113113
rect 184899 113023 184927 113051
rect 184961 113023 184989 113051
rect 184899 112961 184927 112989
rect 184961 112961 184989 112989
rect 177219 110147 177247 110175
rect 177281 110147 177309 110175
rect 177219 110085 177247 110113
rect 177281 110085 177309 110113
rect 177219 110023 177247 110051
rect 177281 110023 177309 110051
rect 177219 109961 177247 109989
rect 177281 109961 177309 109989
rect 187077 110147 187105 110175
rect 187139 110147 187167 110175
rect 187201 110147 187229 110175
rect 187263 110147 187291 110175
rect 187077 110085 187105 110113
rect 187139 110085 187167 110113
rect 187201 110085 187229 110113
rect 187263 110085 187291 110113
rect 187077 110023 187105 110051
rect 187139 110023 187167 110051
rect 187201 110023 187229 110051
rect 187263 110023 187291 110051
rect 187077 109961 187105 109989
rect 187139 109961 187167 109989
rect 187201 109961 187229 109989
rect 187263 109961 187291 109989
rect 173577 104147 173605 104175
rect 173639 104147 173667 104175
rect 173701 104147 173729 104175
rect 173763 104147 173791 104175
rect 173577 104085 173605 104113
rect 173639 104085 173667 104113
rect 173701 104085 173729 104113
rect 173763 104085 173791 104113
rect 173577 104023 173605 104051
rect 173639 104023 173667 104051
rect 173701 104023 173729 104051
rect 173763 104023 173791 104051
rect 173577 103961 173605 103989
rect 173639 103961 173667 103989
rect 173701 103961 173729 103989
rect 173763 103961 173791 103989
rect 184899 104147 184927 104175
rect 184961 104147 184989 104175
rect 184899 104085 184927 104113
rect 184961 104085 184989 104113
rect 184899 104023 184927 104051
rect 184961 104023 184989 104051
rect 184899 103961 184927 103989
rect 184961 103961 184989 103989
rect 177219 101147 177247 101175
rect 177281 101147 177309 101175
rect 177219 101085 177247 101113
rect 177281 101085 177309 101113
rect 177219 101023 177247 101051
rect 177281 101023 177309 101051
rect 177219 100961 177247 100989
rect 177281 100961 177309 100989
rect 187077 101147 187105 101175
rect 187139 101147 187167 101175
rect 187201 101147 187229 101175
rect 187263 101147 187291 101175
rect 187077 101085 187105 101113
rect 187139 101085 187167 101113
rect 187201 101085 187229 101113
rect 187263 101085 187291 101113
rect 187077 101023 187105 101051
rect 187139 101023 187167 101051
rect 187201 101023 187229 101051
rect 187263 101023 187291 101051
rect 187077 100961 187105 100989
rect 187139 100961 187167 100989
rect 187201 100961 187229 100989
rect 187263 100961 187291 100989
rect 173577 95147 173605 95175
rect 173639 95147 173667 95175
rect 173701 95147 173729 95175
rect 173763 95147 173791 95175
rect 173577 95085 173605 95113
rect 173639 95085 173667 95113
rect 173701 95085 173729 95113
rect 173763 95085 173791 95113
rect 173577 95023 173605 95051
rect 173639 95023 173667 95051
rect 173701 95023 173729 95051
rect 173763 95023 173791 95051
rect 173577 94961 173605 94989
rect 173639 94961 173667 94989
rect 173701 94961 173729 94989
rect 173763 94961 173791 94989
rect 184899 95147 184927 95175
rect 184961 95147 184989 95175
rect 184899 95085 184927 95113
rect 184961 95085 184989 95113
rect 184899 95023 184927 95051
rect 184961 95023 184989 95051
rect 184899 94961 184927 94989
rect 184961 94961 184989 94989
rect 177219 92147 177247 92175
rect 177281 92147 177309 92175
rect 177219 92085 177247 92113
rect 177281 92085 177309 92113
rect 177219 92023 177247 92051
rect 177281 92023 177309 92051
rect 177219 91961 177247 91989
rect 177281 91961 177309 91989
rect 187077 92147 187105 92175
rect 187139 92147 187167 92175
rect 187201 92147 187229 92175
rect 187263 92147 187291 92175
rect 187077 92085 187105 92113
rect 187139 92085 187167 92113
rect 187201 92085 187229 92113
rect 187263 92085 187291 92113
rect 187077 92023 187105 92051
rect 187139 92023 187167 92051
rect 187201 92023 187229 92051
rect 187263 92023 187291 92051
rect 187077 91961 187105 91989
rect 187139 91961 187167 91989
rect 187201 91961 187229 91989
rect 187263 91961 187291 91989
rect 173577 86147 173605 86175
rect 173639 86147 173667 86175
rect 173701 86147 173729 86175
rect 173763 86147 173791 86175
rect 173577 86085 173605 86113
rect 173639 86085 173667 86113
rect 173701 86085 173729 86113
rect 173763 86085 173791 86113
rect 173577 86023 173605 86051
rect 173639 86023 173667 86051
rect 173701 86023 173729 86051
rect 173763 86023 173791 86051
rect 173577 85961 173605 85989
rect 173639 85961 173667 85989
rect 173701 85961 173729 85989
rect 173763 85961 173791 85989
rect 184899 86147 184927 86175
rect 184961 86147 184989 86175
rect 184899 86085 184927 86113
rect 184961 86085 184989 86113
rect 184899 86023 184927 86051
rect 184961 86023 184989 86051
rect 184899 85961 184927 85989
rect 184961 85961 184989 85989
rect 177219 83147 177247 83175
rect 177281 83147 177309 83175
rect 177219 83085 177247 83113
rect 177281 83085 177309 83113
rect 177219 83023 177247 83051
rect 177281 83023 177309 83051
rect 177219 82961 177247 82989
rect 177281 82961 177309 82989
rect 187077 83147 187105 83175
rect 187139 83147 187167 83175
rect 187201 83147 187229 83175
rect 187263 83147 187291 83175
rect 187077 83085 187105 83113
rect 187139 83085 187167 83113
rect 187201 83085 187229 83113
rect 187263 83085 187291 83113
rect 187077 83023 187105 83051
rect 187139 83023 187167 83051
rect 187201 83023 187229 83051
rect 187263 83023 187291 83051
rect 187077 82961 187105 82989
rect 187139 82961 187167 82989
rect 187201 82961 187229 82989
rect 187263 82961 187291 82989
rect 173577 77147 173605 77175
rect 173639 77147 173667 77175
rect 173701 77147 173729 77175
rect 173763 77147 173791 77175
rect 173577 77085 173605 77113
rect 173639 77085 173667 77113
rect 173701 77085 173729 77113
rect 173763 77085 173791 77113
rect 173577 77023 173605 77051
rect 173639 77023 173667 77051
rect 173701 77023 173729 77051
rect 173763 77023 173791 77051
rect 173577 76961 173605 76989
rect 173639 76961 173667 76989
rect 173701 76961 173729 76989
rect 173763 76961 173791 76989
rect 184899 77147 184927 77175
rect 184961 77147 184989 77175
rect 184899 77085 184927 77113
rect 184961 77085 184989 77113
rect 184899 77023 184927 77051
rect 184961 77023 184989 77051
rect 184899 76961 184927 76989
rect 184961 76961 184989 76989
rect 177219 74147 177247 74175
rect 177281 74147 177309 74175
rect 177219 74085 177247 74113
rect 177281 74085 177309 74113
rect 177219 74023 177247 74051
rect 177281 74023 177309 74051
rect 177219 73961 177247 73989
rect 177281 73961 177309 73989
rect 187077 74147 187105 74175
rect 187139 74147 187167 74175
rect 187201 74147 187229 74175
rect 187263 74147 187291 74175
rect 187077 74085 187105 74113
rect 187139 74085 187167 74113
rect 187201 74085 187229 74113
rect 187263 74085 187291 74113
rect 187077 74023 187105 74051
rect 187139 74023 187167 74051
rect 187201 74023 187229 74051
rect 187263 74023 187291 74051
rect 187077 73961 187105 73989
rect 187139 73961 187167 73989
rect 187201 73961 187229 73989
rect 187263 73961 187291 73989
rect 173577 68147 173605 68175
rect 173639 68147 173667 68175
rect 173701 68147 173729 68175
rect 173763 68147 173791 68175
rect 173577 68085 173605 68113
rect 173639 68085 173667 68113
rect 173701 68085 173729 68113
rect 173763 68085 173791 68113
rect 173577 68023 173605 68051
rect 173639 68023 173667 68051
rect 173701 68023 173729 68051
rect 173763 68023 173791 68051
rect 173577 67961 173605 67989
rect 173639 67961 173667 67989
rect 173701 67961 173729 67989
rect 173763 67961 173791 67989
rect 184899 68147 184927 68175
rect 184961 68147 184989 68175
rect 184899 68085 184927 68113
rect 184961 68085 184989 68113
rect 184899 68023 184927 68051
rect 184961 68023 184989 68051
rect 184899 67961 184927 67989
rect 184961 67961 184989 67989
rect 177219 65147 177247 65175
rect 177281 65147 177309 65175
rect 177219 65085 177247 65113
rect 177281 65085 177309 65113
rect 177219 65023 177247 65051
rect 177281 65023 177309 65051
rect 177219 64961 177247 64989
rect 177281 64961 177309 64989
rect 187077 65147 187105 65175
rect 187139 65147 187167 65175
rect 187201 65147 187229 65175
rect 187263 65147 187291 65175
rect 187077 65085 187105 65113
rect 187139 65085 187167 65113
rect 187201 65085 187229 65113
rect 187263 65085 187291 65113
rect 187077 65023 187105 65051
rect 187139 65023 187167 65051
rect 187201 65023 187229 65051
rect 187263 65023 187291 65051
rect 187077 64961 187105 64989
rect 187139 64961 187167 64989
rect 187201 64961 187229 64989
rect 187263 64961 187291 64989
rect 173577 59147 173605 59175
rect 173639 59147 173667 59175
rect 173701 59147 173729 59175
rect 173763 59147 173791 59175
rect 173577 59085 173605 59113
rect 173639 59085 173667 59113
rect 173701 59085 173729 59113
rect 173763 59085 173791 59113
rect 173577 59023 173605 59051
rect 173639 59023 173667 59051
rect 173701 59023 173729 59051
rect 173763 59023 173791 59051
rect 173577 58961 173605 58989
rect 173639 58961 173667 58989
rect 173701 58961 173729 58989
rect 173763 58961 173791 58989
rect 184899 59147 184927 59175
rect 184961 59147 184989 59175
rect 184899 59085 184927 59113
rect 184961 59085 184989 59113
rect 184899 59023 184927 59051
rect 184961 59023 184989 59051
rect 184899 58961 184927 58989
rect 184961 58961 184989 58989
rect 177219 56147 177247 56175
rect 177281 56147 177309 56175
rect 177219 56085 177247 56113
rect 177281 56085 177309 56113
rect 177219 56023 177247 56051
rect 177281 56023 177309 56051
rect 177219 55961 177247 55989
rect 177281 55961 177309 55989
rect 187077 56147 187105 56175
rect 187139 56147 187167 56175
rect 187201 56147 187229 56175
rect 187263 56147 187291 56175
rect 187077 56085 187105 56113
rect 187139 56085 187167 56113
rect 187201 56085 187229 56113
rect 187263 56085 187291 56113
rect 187077 56023 187105 56051
rect 187139 56023 187167 56051
rect 187201 56023 187229 56051
rect 187263 56023 187291 56051
rect 187077 55961 187105 55989
rect 187139 55961 187167 55989
rect 187201 55961 187229 55989
rect 187263 55961 187291 55989
rect 173577 50147 173605 50175
rect 173639 50147 173667 50175
rect 173701 50147 173729 50175
rect 173763 50147 173791 50175
rect 173577 50085 173605 50113
rect 173639 50085 173667 50113
rect 173701 50085 173729 50113
rect 173763 50085 173791 50113
rect 173577 50023 173605 50051
rect 173639 50023 173667 50051
rect 173701 50023 173729 50051
rect 173763 50023 173791 50051
rect 173577 49961 173605 49989
rect 173639 49961 173667 49989
rect 173701 49961 173729 49989
rect 173763 49961 173791 49989
rect 184899 50147 184927 50175
rect 184961 50147 184989 50175
rect 184899 50085 184927 50113
rect 184961 50085 184989 50113
rect 184899 50023 184927 50051
rect 184961 50023 184989 50051
rect 184899 49961 184927 49989
rect 184961 49961 184989 49989
rect 177219 47147 177247 47175
rect 177281 47147 177309 47175
rect 177219 47085 177247 47113
rect 177281 47085 177309 47113
rect 177219 47023 177247 47051
rect 177281 47023 177309 47051
rect 177219 46961 177247 46989
rect 177281 46961 177309 46989
rect 187077 47147 187105 47175
rect 187139 47147 187167 47175
rect 187201 47147 187229 47175
rect 187263 47147 187291 47175
rect 187077 47085 187105 47113
rect 187139 47085 187167 47113
rect 187201 47085 187229 47113
rect 187263 47085 187291 47113
rect 187077 47023 187105 47051
rect 187139 47023 187167 47051
rect 187201 47023 187229 47051
rect 187263 47023 187291 47051
rect 187077 46961 187105 46989
rect 187139 46961 187167 46989
rect 187201 46961 187229 46989
rect 187263 46961 187291 46989
rect 173577 41147 173605 41175
rect 173639 41147 173667 41175
rect 173701 41147 173729 41175
rect 173763 41147 173791 41175
rect 173577 41085 173605 41113
rect 173639 41085 173667 41113
rect 173701 41085 173729 41113
rect 173763 41085 173791 41113
rect 173577 41023 173605 41051
rect 173639 41023 173667 41051
rect 173701 41023 173729 41051
rect 173763 41023 173791 41051
rect 173577 40961 173605 40989
rect 173639 40961 173667 40989
rect 173701 40961 173729 40989
rect 173763 40961 173791 40989
rect 184899 41147 184927 41175
rect 184961 41147 184989 41175
rect 184899 41085 184927 41113
rect 184961 41085 184989 41113
rect 184899 41023 184927 41051
rect 184961 41023 184989 41051
rect 184899 40961 184927 40989
rect 184961 40961 184989 40989
rect 177219 38147 177247 38175
rect 177281 38147 177309 38175
rect 177219 38085 177247 38113
rect 177281 38085 177309 38113
rect 177219 38023 177247 38051
rect 177281 38023 177309 38051
rect 177219 37961 177247 37989
rect 177281 37961 177309 37989
rect 187077 38147 187105 38175
rect 187139 38147 187167 38175
rect 187201 38147 187229 38175
rect 187263 38147 187291 38175
rect 187077 38085 187105 38113
rect 187139 38085 187167 38113
rect 187201 38085 187229 38113
rect 187263 38085 187291 38113
rect 187077 38023 187105 38051
rect 187139 38023 187167 38051
rect 187201 38023 187229 38051
rect 187263 38023 187291 38051
rect 187077 37961 187105 37989
rect 187139 37961 187167 37989
rect 187201 37961 187229 37989
rect 187263 37961 187291 37989
rect 173577 32147 173605 32175
rect 173639 32147 173667 32175
rect 173701 32147 173729 32175
rect 173763 32147 173791 32175
rect 173577 32085 173605 32113
rect 173639 32085 173667 32113
rect 173701 32085 173729 32113
rect 173763 32085 173791 32113
rect 173577 32023 173605 32051
rect 173639 32023 173667 32051
rect 173701 32023 173729 32051
rect 173763 32023 173791 32051
rect 173577 31961 173605 31989
rect 173639 31961 173667 31989
rect 173701 31961 173729 31989
rect 173763 31961 173791 31989
rect 184899 32147 184927 32175
rect 184961 32147 184989 32175
rect 184899 32085 184927 32113
rect 184961 32085 184989 32113
rect 184899 32023 184927 32051
rect 184961 32023 184989 32051
rect 184899 31961 184927 31989
rect 184961 31961 184989 31989
rect 177219 29147 177247 29175
rect 177281 29147 177309 29175
rect 177219 29085 177247 29113
rect 177281 29085 177309 29113
rect 177219 29023 177247 29051
rect 177281 29023 177309 29051
rect 177219 28961 177247 28989
rect 177281 28961 177309 28989
rect 187077 29147 187105 29175
rect 187139 29147 187167 29175
rect 187201 29147 187229 29175
rect 187263 29147 187291 29175
rect 187077 29085 187105 29113
rect 187139 29085 187167 29113
rect 187201 29085 187229 29113
rect 187263 29085 187291 29113
rect 187077 29023 187105 29051
rect 187139 29023 187167 29051
rect 187201 29023 187229 29051
rect 187263 29023 187291 29051
rect 187077 28961 187105 28989
rect 187139 28961 187167 28989
rect 187201 28961 187229 28989
rect 187263 28961 187291 28989
rect 173577 23147 173605 23175
rect 173639 23147 173667 23175
rect 173701 23147 173729 23175
rect 173763 23147 173791 23175
rect 173577 23085 173605 23113
rect 173639 23085 173667 23113
rect 173701 23085 173729 23113
rect 173763 23085 173791 23113
rect 173577 23023 173605 23051
rect 173639 23023 173667 23051
rect 173701 23023 173729 23051
rect 173763 23023 173791 23051
rect 173577 22961 173605 22989
rect 173639 22961 173667 22989
rect 173701 22961 173729 22989
rect 173763 22961 173791 22989
rect 184899 23147 184927 23175
rect 184961 23147 184989 23175
rect 184899 23085 184927 23113
rect 184961 23085 184989 23113
rect 184899 23023 184927 23051
rect 184961 23023 184989 23051
rect 184899 22961 184927 22989
rect 184961 22961 184989 22989
rect 177219 20147 177247 20175
rect 177281 20147 177309 20175
rect 177219 20085 177247 20113
rect 177281 20085 177309 20113
rect 177219 20023 177247 20051
rect 177281 20023 177309 20051
rect 177219 19961 177247 19989
rect 177281 19961 177309 19989
rect 187077 20147 187105 20175
rect 187139 20147 187167 20175
rect 187201 20147 187229 20175
rect 187263 20147 187291 20175
rect 187077 20085 187105 20113
rect 187139 20085 187167 20113
rect 187201 20085 187229 20113
rect 187263 20085 187291 20113
rect 187077 20023 187105 20051
rect 187139 20023 187167 20051
rect 187201 20023 187229 20051
rect 187263 20023 187291 20051
rect 187077 19961 187105 19989
rect 187139 19961 187167 19989
rect 187201 19961 187229 19989
rect 187263 19961 187291 19989
rect 173577 14147 173605 14175
rect 173639 14147 173667 14175
rect 173701 14147 173729 14175
rect 173763 14147 173791 14175
rect 173577 14085 173605 14113
rect 173639 14085 173667 14113
rect 173701 14085 173729 14113
rect 173763 14085 173791 14113
rect 173577 14023 173605 14051
rect 173639 14023 173667 14051
rect 173701 14023 173729 14051
rect 173763 14023 173791 14051
rect 173577 13961 173605 13989
rect 173639 13961 173667 13989
rect 173701 13961 173729 13989
rect 173763 13961 173791 13989
rect 184899 14147 184927 14175
rect 184961 14147 184989 14175
rect 184899 14085 184927 14113
rect 184961 14085 184989 14113
rect 184899 14023 184927 14051
rect 184961 14023 184989 14051
rect 184899 13961 184927 13989
rect 184961 13961 184989 13989
rect 177219 11147 177247 11175
rect 177281 11147 177309 11175
rect 177219 11085 177247 11113
rect 177281 11085 177309 11113
rect 177219 11023 177247 11051
rect 177281 11023 177309 11051
rect 177219 10961 177247 10989
rect 177281 10961 177309 10989
rect 187077 11147 187105 11175
rect 187139 11147 187167 11175
rect 187201 11147 187229 11175
rect 187263 11147 187291 11175
rect 187077 11085 187105 11113
rect 187139 11085 187167 11113
rect 187201 11085 187229 11113
rect 187263 11085 187291 11113
rect 187077 11023 187105 11051
rect 187139 11023 187167 11051
rect 187201 11023 187229 11051
rect 187263 11023 187291 11051
rect 187077 10961 187105 10989
rect 187139 10961 187167 10989
rect 187201 10961 187229 10989
rect 187263 10961 187291 10989
rect 173577 5147 173605 5175
rect 173639 5147 173667 5175
rect 173701 5147 173729 5175
rect 173763 5147 173791 5175
rect 173577 5085 173605 5113
rect 173639 5085 173667 5113
rect 173701 5085 173729 5113
rect 173763 5085 173791 5113
rect 173577 5023 173605 5051
rect 173639 5023 173667 5051
rect 173701 5023 173729 5051
rect 173763 5023 173791 5051
rect 173577 4961 173605 4989
rect 173639 4961 173667 4989
rect 173701 4961 173729 4989
rect 173763 4961 173791 4989
rect 184899 5147 184927 5175
rect 184961 5147 184989 5175
rect 184899 5085 184927 5113
rect 184961 5085 184989 5113
rect 184899 5023 184927 5051
rect 184961 5023 184989 5051
rect 184899 4961 184927 4989
rect 184961 4961 184989 4989
rect 173577 -588 173605 -560
rect 173639 -588 173667 -560
rect 173701 -588 173729 -560
rect 173763 -588 173791 -560
rect 173577 -650 173605 -622
rect 173639 -650 173667 -622
rect 173701 -650 173729 -622
rect 173763 -650 173791 -622
rect 173577 -712 173605 -684
rect 173639 -712 173667 -684
rect 173701 -712 173729 -684
rect 173763 -712 173791 -684
rect 173577 -774 173605 -746
rect 173639 -774 173667 -746
rect 173701 -774 173729 -746
rect 173763 -774 173791 -746
rect 187077 2147 187105 2175
rect 187139 2147 187167 2175
rect 187201 2147 187229 2175
rect 187263 2147 187291 2175
rect 187077 2085 187105 2113
rect 187139 2085 187167 2113
rect 187201 2085 187229 2113
rect 187263 2085 187291 2113
rect 187077 2023 187105 2051
rect 187139 2023 187167 2051
rect 187201 2023 187229 2051
rect 187263 2023 187291 2051
rect 187077 1961 187105 1989
rect 187139 1961 187167 1989
rect 187201 1961 187229 1989
rect 187263 1961 187291 1989
rect 187077 -108 187105 -80
rect 187139 -108 187167 -80
rect 187201 -108 187229 -80
rect 187263 -108 187291 -80
rect 187077 -170 187105 -142
rect 187139 -170 187167 -142
rect 187201 -170 187229 -142
rect 187263 -170 187291 -142
rect 187077 -232 187105 -204
rect 187139 -232 187167 -204
rect 187201 -232 187229 -204
rect 187263 -232 187291 -204
rect 187077 -294 187105 -266
rect 187139 -294 187167 -266
rect 187201 -294 187229 -266
rect 187263 -294 187291 -266
rect 188937 299058 188965 299086
rect 188999 299058 189027 299086
rect 189061 299058 189089 299086
rect 189123 299058 189151 299086
rect 188937 298996 188965 299024
rect 188999 298996 189027 299024
rect 189061 298996 189089 299024
rect 189123 298996 189151 299024
rect 188937 298934 188965 298962
rect 188999 298934 189027 298962
rect 189061 298934 189089 298962
rect 189123 298934 189151 298962
rect 188937 298872 188965 298900
rect 188999 298872 189027 298900
rect 189061 298872 189089 298900
rect 189123 298872 189151 298900
rect 188937 293147 188965 293175
rect 188999 293147 189027 293175
rect 189061 293147 189089 293175
rect 189123 293147 189151 293175
rect 188937 293085 188965 293113
rect 188999 293085 189027 293113
rect 189061 293085 189089 293113
rect 189123 293085 189151 293113
rect 188937 293023 188965 293051
rect 188999 293023 189027 293051
rect 189061 293023 189089 293051
rect 189123 293023 189151 293051
rect 188937 292961 188965 292989
rect 188999 292961 189027 292989
rect 189061 292961 189089 292989
rect 189123 292961 189151 292989
rect 188937 284147 188965 284175
rect 188999 284147 189027 284175
rect 189061 284147 189089 284175
rect 189123 284147 189151 284175
rect 188937 284085 188965 284113
rect 188999 284085 189027 284113
rect 189061 284085 189089 284113
rect 189123 284085 189151 284113
rect 188937 284023 188965 284051
rect 188999 284023 189027 284051
rect 189061 284023 189089 284051
rect 189123 284023 189151 284051
rect 188937 283961 188965 283989
rect 188999 283961 189027 283989
rect 189061 283961 189089 283989
rect 189123 283961 189151 283989
rect 188937 275147 188965 275175
rect 188999 275147 189027 275175
rect 189061 275147 189089 275175
rect 189123 275147 189151 275175
rect 188937 275085 188965 275113
rect 188999 275085 189027 275113
rect 189061 275085 189089 275113
rect 189123 275085 189151 275113
rect 188937 275023 188965 275051
rect 188999 275023 189027 275051
rect 189061 275023 189089 275051
rect 189123 275023 189151 275051
rect 188937 274961 188965 274989
rect 188999 274961 189027 274989
rect 189061 274961 189089 274989
rect 189123 274961 189151 274989
rect 188937 266147 188965 266175
rect 188999 266147 189027 266175
rect 189061 266147 189089 266175
rect 189123 266147 189151 266175
rect 188937 266085 188965 266113
rect 188999 266085 189027 266113
rect 189061 266085 189089 266113
rect 189123 266085 189151 266113
rect 188937 266023 188965 266051
rect 188999 266023 189027 266051
rect 189061 266023 189089 266051
rect 189123 266023 189151 266051
rect 188937 265961 188965 265989
rect 188999 265961 189027 265989
rect 189061 265961 189089 265989
rect 189123 265961 189151 265989
rect 188937 257147 188965 257175
rect 188999 257147 189027 257175
rect 189061 257147 189089 257175
rect 189123 257147 189151 257175
rect 188937 257085 188965 257113
rect 188999 257085 189027 257113
rect 189061 257085 189089 257113
rect 189123 257085 189151 257113
rect 188937 257023 188965 257051
rect 188999 257023 189027 257051
rect 189061 257023 189089 257051
rect 189123 257023 189151 257051
rect 188937 256961 188965 256989
rect 188999 256961 189027 256989
rect 189061 256961 189089 256989
rect 189123 256961 189151 256989
rect 188937 248147 188965 248175
rect 188999 248147 189027 248175
rect 189061 248147 189089 248175
rect 189123 248147 189151 248175
rect 188937 248085 188965 248113
rect 188999 248085 189027 248113
rect 189061 248085 189089 248113
rect 189123 248085 189151 248113
rect 188937 248023 188965 248051
rect 188999 248023 189027 248051
rect 189061 248023 189089 248051
rect 189123 248023 189151 248051
rect 188937 247961 188965 247989
rect 188999 247961 189027 247989
rect 189061 247961 189089 247989
rect 189123 247961 189151 247989
rect 188937 239147 188965 239175
rect 188999 239147 189027 239175
rect 189061 239147 189089 239175
rect 189123 239147 189151 239175
rect 188937 239085 188965 239113
rect 188999 239085 189027 239113
rect 189061 239085 189089 239113
rect 189123 239085 189151 239113
rect 188937 239023 188965 239051
rect 188999 239023 189027 239051
rect 189061 239023 189089 239051
rect 189123 239023 189151 239051
rect 188937 238961 188965 238989
rect 188999 238961 189027 238989
rect 189061 238961 189089 238989
rect 189123 238961 189151 238989
rect 188937 230147 188965 230175
rect 188999 230147 189027 230175
rect 189061 230147 189089 230175
rect 189123 230147 189151 230175
rect 188937 230085 188965 230113
rect 188999 230085 189027 230113
rect 189061 230085 189089 230113
rect 189123 230085 189151 230113
rect 188937 230023 188965 230051
rect 188999 230023 189027 230051
rect 189061 230023 189089 230051
rect 189123 230023 189151 230051
rect 188937 229961 188965 229989
rect 188999 229961 189027 229989
rect 189061 229961 189089 229989
rect 189123 229961 189151 229989
rect 188937 221147 188965 221175
rect 188999 221147 189027 221175
rect 189061 221147 189089 221175
rect 189123 221147 189151 221175
rect 188937 221085 188965 221113
rect 188999 221085 189027 221113
rect 189061 221085 189089 221113
rect 189123 221085 189151 221113
rect 188937 221023 188965 221051
rect 188999 221023 189027 221051
rect 189061 221023 189089 221051
rect 189123 221023 189151 221051
rect 188937 220961 188965 220989
rect 188999 220961 189027 220989
rect 189061 220961 189089 220989
rect 189123 220961 189151 220989
rect 188937 212147 188965 212175
rect 188999 212147 189027 212175
rect 189061 212147 189089 212175
rect 189123 212147 189151 212175
rect 188937 212085 188965 212113
rect 188999 212085 189027 212113
rect 189061 212085 189089 212113
rect 189123 212085 189151 212113
rect 188937 212023 188965 212051
rect 188999 212023 189027 212051
rect 189061 212023 189089 212051
rect 189123 212023 189151 212051
rect 188937 211961 188965 211989
rect 188999 211961 189027 211989
rect 189061 211961 189089 211989
rect 189123 211961 189151 211989
rect 188937 203147 188965 203175
rect 188999 203147 189027 203175
rect 189061 203147 189089 203175
rect 189123 203147 189151 203175
rect 188937 203085 188965 203113
rect 188999 203085 189027 203113
rect 189061 203085 189089 203113
rect 189123 203085 189151 203113
rect 188937 203023 188965 203051
rect 188999 203023 189027 203051
rect 189061 203023 189089 203051
rect 189123 203023 189151 203051
rect 188937 202961 188965 202989
rect 188999 202961 189027 202989
rect 189061 202961 189089 202989
rect 189123 202961 189151 202989
rect 188937 194147 188965 194175
rect 188999 194147 189027 194175
rect 189061 194147 189089 194175
rect 189123 194147 189151 194175
rect 188937 194085 188965 194113
rect 188999 194085 189027 194113
rect 189061 194085 189089 194113
rect 189123 194085 189151 194113
rect 188937 194023 188965 194051
rect 188999 194023 189027 194051
rect 189061 194023 189089 194051
rect 189123 194023 189151 194051
rect 188937 193961 188965 193989
rect 188999 193961 189027 193989
rect 189061 193961 189089 193989
rect 189123 193961 189151 193989
rect 188937 185147 188965 185175
rect 188999 185147 189027 185175
rect 189061 185147 189089 185175
rect 189123 185147 189151 185175
rect 188937 185085 188965 185113
rect 188999 185085 189027 185113
rect 189061 185085 189089 185113
rect 189123 185085 189151 185113
rect 188937 185023 188965 185051
rect 188999 185023 189027 185051
rect 189061 185023 189089 185051
rect 189123 185023 189151 185051
rect 188937 184961 188965 184989
rect 188999 184961 189027 184989
rect 189061 184961 189089 184989
rect 189123 184961 189151 184989
rect 188937 176147 188965 176175
rect 188999 176147 189027 176175
rect 189061 176147 189089 176175
rect 189123 176147 189151 176175
rect 188937 176085 188965 176113
rect 188999 176085 189027 176113
rect 189061 176085 189089 176113
rect 189123 176085 189151 176113
rect 188937 176023 188965 176051
rect 188999 176023 189027 176051
rect 189061 176023 189089 176051
rect 189123 176023 189151 176051
rect 188937 175961 188965 175989
rect 188999 175961 189027 175989
rect 189061 175961 189089 175989
rect 189123 175961 189151 175989
rect 202437 298578 202465 298606
rect 202499 298578 202527 298606
rect 202561 298578 202589 298606
rect 202623 298578 202651 298606
rect 202437 298516 202465 298544
rect 202499 298516 202527 298544
rect 202561 298516 202589 298544
rect 202623 298516 202651 298544
rect 202437 298454 202465 298482
rect 202499 298454 202527 298482
rect 202561 298454 202589 298482
rect 202623 298454 202651 298482
rect 202437 298392 202465 298420
rect 202499 298392 202527 298420
rect 202561 298392 202589 298420
rect 202623 298392 202651 298420
rect 202437 290147 202465 290175
rect 202499 290147 202527 290175
rect 202561 290147 202589 290175
rect 202623 290147 202651 290175
rect 202437 290085 202465 290113
rect 202499 290085 202527 290113
rect 202561 290085 202589 290113
rect 202623 290085 202651 290113
rect 202437 290023 202465 290051
rect 202499 290023 202527 290051
rect 202561 290023 202589 290051
rect 202623 290023 202651 290051
rect 202437 289961 202465 289989
rect 202499 289961 202527 289989
rect 202561 289961 202589 289989
rect 202623 289961 202651 289989
rect 202437 281147 202465 281175
rect 202499 281147 202527 281175
rect 202561 281147 202589 281175
rect 202623 281147 202651 281175
rect 202437 281085 202465 281113
rect 202499 281085 202527 281113
rect 202561 281085 202589 281113
rect 202623 281085 202651 281113
rect 202437 281023 202465 281051
rect 202499 281023 202527 281051
rect 202561 281023 202589 281051
rect 202623 281023 202651 281051
rect 202437 280961 202465 280989
rect 202499 280961 202527 280989
rect 202561 280961 202589 280989
rect 202623 280961 202651 280989
rect 202437 272147 202465 272175
rect 202499 272147 202527 272175
rect 202561 272147 202589 272175
rect 202623 272147 202651 272175
rect 202437 272085 202465 272113
rect 202499 272085 202527 272113
rect 202561 272085 202589 272113
rect 202623 272085 202651 272113
rect 202437 272023 202465 272051
rect 202499 272023 202527 272051
rect 202561 272023 202589 272051
rect 202623 272023 202651 272051
rect 202437 271961 202465 271989
rect 202499 271961 202527 271989
rect 202561 271961 202589 271989
rect 202623 271961 202651 271989
rect 202437 263147 202465 263175
rect 202499 263147 202527 263175
rect 202561 263147 202589 263175
rect 202623 263147 202651 263175
rect 202437 263085 202465 263113
rect 202499 263085 202527 263113
rect 202561 263085 202589 263113
rect 202623 263085 202651 263113
rect 202437 263023 202465 263051
rect 202499 263023 202527 263051
rect 202561 263023 202589 263051
rect 202623 263023 202651 263051
rect 202437 262961 202465 262989
rect 202499 262961 202527 262989
rect 202561 262961 202589 262989
rect 202623 262961 202651 262989
rect 202437 254147 202465 254175
rect 202499 254147 202527 254175
rect 202561 254147 202589 254175
rect 202623 254147 202651 254175
rect 202437 254085 202465 254113
rect 202499 254085 202527 254113
rect 202561 254085 202589 254113
rect 202623 254085 202651 254113
rect 202437 254023 202465 254051
rect 202499 254023 202527 254051
rect 202561 254023 202589 254051
rect 202623 254023 202651 254051
rect 202437 253961 202465 253989
rect 202499 253961 202527 253989
rect 202561 253961 202589 253989
rect 202623 253961 202651 253989
rect 202437 245147 202465 245175
rect 202499 245147 202527 245175
rect 202561 245147 202589 245175
rect 202623 245147 202651 245175
rect 202437 245085 202465 245113
rect 202499 245085 202527 245113
rect 202561 245085 202589 245113
rect 202623 245085 202651 245113
rect 202437 245023 202465 245051
rect 202499 245023 202527 245051
rect 202561 245023 202589 245051
rect 202623 245023 202651 245051
rect 202437 244961 202465 244989
rect 202499 244961 202527 244989
rect 202561 244961 202589 244989
rect 202623 244961 202651 244989
rect 202437 236147 202465 236175
rect 202499 236147 202527 236175
rect 202561 236147 202589 236175
rect 202623 236147 202651 236175
rect 202437 236085 202465 236113
rect 202499 236085 202527 236113
rect 202561 236085 202589 236113
rect 202623 236085 202651 236113
rect 202437 236023 202465 236051
rect 202499 236023 202527 236051
rect 202561 236023 202589 236051
rect 202623 236023 202651 236051
rect 202437 235961 202465 235989
rect 202499 235961 202527 235989
rect 202561 235961 202589 235989
rect 202623 235961 202651 235989
rect 202437 227147 202465 227175
rect 202499 227147 202527 227175
rect 202561 227147 202589 227175
rect 202623 227147 202651 227175
rect 202437 227085 202465 227113
rect 202499 227085 202527 227113
rect 202561 227085 202589 227113
rect 202623 227085 202651 227113
rect 202437 227023 202465 227051
rect 202499 227023 202527 227051
rect 202561 227023 202589 227051
rect 202623 227023 202651 227051
rect 202437 226961 202465 226989
rect 202499 226961 202527 226989
rect 202561 226961 202589 226989
rect 202623 226961 202651 226989
rect 202437 218147 202465 218175
rect 202499 218147 202527 218175
rect 202561 218147 202589 218175
rect 202623 218147 202651 218175
rect 202437 218085 202465 218113
rect 202499 218085 202527 218113
rect 202561 218085 202589 218113
rect 202623 218085 202651 218113
rect 202437 218023 202465 218051
rect 202499 218023 202527 218051
rect 202561 218023 202589 218051
rect 202623 218023 202651 218051
rect 202437 217961 202465 217989
rect 202499 217961 202527 217989
rect 202561 217961 202589 217989
rect 202623 217961 202651 217989
rect 202437 209147 202465 209175
rect 202499 209147 202527 209175
rect 202561 209147 202589 209175
rect 202623 209147 202651 209175
rect 202437 209085 202465 209113
rect 202499 209085 202527 209113
rect 202561 209085 202589 209113
rect 202623 209085 202651 209113
rect 202437 209023 202465 209051
rect 202499 209023 202527 209051
rect 202561 209023 202589 209051
rect 202623 209023 202651 209051
rect 202437 208961 202465 208989
rect 202499 208961 202527 208989
rect 202561 208961 202589 208989
rect 202623 208961 202651 208989
rect 202437 200147 202465 200175
rect 202499 200147 202527 200175
rect 202561 200147 202589 200175
rect 202623 200147 202651 200175
rect 202437 200085 202465 200113
rect 202499 200085 202527 200113
rect 202561 200085 202589 200113
rect 202623 200085 202651 200113
rect 202437 200023 202465 200051
rect 202499 200023 202527 200051
rect 202561 200023 202589 200051
rect 202623 200023 202651 200051
rect 202437 199961 202465 199989
rect 202499 199961 202527 199989
rect 202561 199961 202589 199989
rect 202623 199961 202651 199989
rect 202437 191147 202465 191175
rect 202499 191147 202527 191175
rect 202561 191147 202589 191175
rect 202623 191147 202651 191175
rect 202437 191085 202465 191113
rect 202499 191085 202527 191113
rect 202561 191085 202589 191113
rect 202623 191085 202651 191113
rect 202437 191023 202465 191051
rect 202499 191023 202527 191051
rect 202561 191023 202589 191051
rect 202623 191023 202651 191051
rect 202437 190961 202465 190989
rect 202499 190961 202527 190989
rect 202561 190961 202589 190989
rect 202623 190961 202651 190989
rect 202437 182147 202465 182175
rect 202499 182147 202527 182175
rect 202561 182147 202589 182175
rect 202623 182147 202651 182175
rect 202437 182085 202465 182113
rect 202499 182085 202527 182113
rect 202561 182085 202589 182113
rect 202623 182085 202651 182113
rect 202437 182023 202465 182051
rect 202499 182023 202527 182051
rect 202561 182023 202589 182051
rect 202623 182023 202651 182051
rect 202437 181961 202465 181989
rect 202499 181961 202527 181989
rect 202561 181961 202589 181989
rect 202623 181961 202651 181989
rect 192579 173147 192607 173175
rect 192641 173147 192669 173175
rect 192579 173085 192607 173113
rect 192641 173085 192669 173113
rect 192579 173023 192607 173051
rect 192641 173023 192669 173051
rect 192579 172961 192607 172989
rect 192641 172961 192669 172989
rect 202437 173147 202465 173175
rect 202499 173147 202527 173175
rect 202561 173147 202589 173175
rect 202623 173147 202651 173175
rect 202437 173085 202465 173113
rect 202499 173085 202527 173113
rect 202561 173085 202589 173113
rect 202623 173085 202651 173113
rect 202437 173023 202465 173051
rect 202499 173023 202527 173051
rect 202561 173023 202589 173051
rect 202623 173023 202651 173051
rect 202437 172961 202465 172989
rect 202499 172961 202527 172989
rect 202561 172961 202589 172989
rect 202623 172961 202651 172989
rect 188937 167147 188965 167175
rect 188999 167147 189027 167175
rect 189061 167147 189089 167175
rect 189123 167147 189151 167175
rect 188937 167085 188965 167113
rect 188999 167085 189027 167113
rect 189061 167085 189089 167113
rect 189123 167085 189151 167113
rect 188937 167023 188965 167051
rect 188999 167023 189027 167051
rect 189061 167023 189089 167051
rect 189123 167023 189151 167051
rect 188937 166961 188965 166989
rect 188999 166961 189027 166989
rect 189061 166961 189089 166989
rect 189123 166961 189151 166989
rect 200259 167147 200287 167175
rect 200321 167147 200349 167175
rect 200259 167085 200287 167113
rect 200321 167085 200349 167113
rect 200259 167023 200287 167051
rect 200321 167023 200349 167051
rect 200259 166961 200287 166989
rect 200321 166961 200349 166989
rect 192579 164147 192607 164175
rect 192641 164147 192669 164175
rect 192579 164085 192607 164113
rect 192641 164085 192669 164113
rect 192579 164023 192607 164051
rect 192641 164023 192669 164051
rect 192579 163961 192607 163989
rect 192641 163961 192669 163989
rect 202437 164147 202465 164175
rect 202499 164147 202527 164175
rect 202561 164147 202589 164175
rect 202623 164147 202651 164175
rect 202437 164085 202465 164113
rect 202499 164085 202527 164113
rect 202561 164085 202589 164113
rect 202623 164085 202651 164113
rect 202437 164023 202465 164051
rect 202499 164023 202527 164051
rect 202561 164023 202589 164051
rect 202623 164023 202651 164051
rect 202437 163961 202465 163989
rect 202499 163961 202527 163989
rect 202561 163961 202589 163989
rect 202623 163961 202651 163989
rect 188937 158147 188965 158175
rect 188999 158147 189027 158175
rect 189061 158147 189089 158175
rect 189123 158147 189151 158175
rect 188937 158085 188965 158113
rect 188999 158085 189027 158113
rect 189061 158085 189089 158113
rect 189123 158085 189151 158113
rect 188937 158023 188965 158051
rect 188999 158023 189027 158051
rect 189061 158023 189089 158051
rect 189123 158023 189151 158051
rect 188937 157961 188965 157989
rect 188999 157961 189027 157989
rect 189061 157961 189089 157989
rect 189123 157961 189151 157989
rect 200259 158147 200287 158175
rect 200321 158147 200349 158175
rect 200259 158085 200287 158113
rect 200321 158085 200349 158113
rect 200259 158023 200287 158051
rect 200321 158023 200349 158051
rect 200259 157961 200287 157989
rect 200321 157961 200349 157989
rect 192579 155147 192607 155175
rect 192641 155147 192669 155175
rect 192579 155085 192607 155113
rect 192641 155085 192669 155113
rect 192579 155023 192607 155051
rect 192641 155023 192669 155051
rect 192579 154961 192607 154989
rect 192641 154961 192669 154989
rect 202437 155147 202465 155175
rect 202499 155147 202527 155175
rect 202561 155147 202589 155175
rect 202623 155147 202651 155175
rect 202437 155085 202465 155113
rect 202499 155085 202527 155113
rect 202561 155085 202589 155113
rect 202623 155085 202651 155113
rect 202437 155023 202465 155051
rect 202499 155023 202527 155051
rect 202561 155023 202589 155051
rect 202623 155023 202651 155051
rect 202437 154961 202465 154989
rect 202499 154961 202527 154989
rect 202561 154961 202589 154989
rect 202623 154961 202651 154989
rect 188937 149147 188965 149175
rect 188999 149147 189027 149175
rect 189061 149147 189089 149175
rect 189123 149147 189151 149175
rect 188937 149085 188965 149113
rect 188999 149085 189027 149113
rect 189061 149085 189089 149113
rect 189123 149085 189151 149113
rect 188937 149023 188965 149051
rect 188999 149023 189027 149051
rect 189061 149023 189089 149051
rect 189123 149023 189151 149051
rect 188937 148961 188965 148989
rect 188999 148961 189027 148989
rect 189061 148961 189089 148989
rect 189123 148961 189151 148989
rect 200259 149147 200287 149175
rect 200321 149147 200349 149175
rect 200259 149085 200287 149113
rect 200321 149085 200349 149113
rect 200259 149023 200287 149051
rect 200321 149023 200349 149051
rect 200259 148961 200287 148989
rect 200321 148961 200349 148989
rect 192579 146147 192607 146175
rect 192641 146147 192669 146175
rect 192579 146085 192607 146113
rect 192641 146085 192669 146113
rect 192579 146023 192607 146051
rect 192641 146023 192669 146051
rect 192579 145961 192607 145989
rect 192641 145961 192669 145989
rect 202437 146147 202465 146175
rect 202499 146147 202527 146175
rect 202561 146147 202589 146175
rect 202623 146147 202651 146175
rect 202437 146085 202465 146113
rect 202499 146085 202527 146113
rect 202561 146085 202589 146113
rect 202623 146085 202651 146113
rect 202437 146023 202465 146051
rect 202499 146023 202527 146051
rect 202561 146023 202589 146051
rect 202623 146023 202651 146051
rect 202437 145961 202465 145989
rect 202499 145961 202527 145989
rect 202561 145961 202589 145989
rect 202623 145961 202651 145989
rect 188937 140147 188965 140175
rect 188999 140147 189027 140175
rect 189061 140147 189089 140175
rect 189123 140147 189151 140175
rect 188937 140085 188965 140113
rect 188999 140085 189027 140113
rect 189061 140085 189089 140113
rect 189123 140085 189151 140113
rect 188937 140023 188965 140051
rect 188999 140023 189027 140051
rect 189061 140023 189089 140051
rect 189123 140023 189151 140051
rect 188937 139961 188965 139989
rect 188999 139961 189027 139989
rect 189061 139961 189089 139989
rect 189123 139961 189151 139989
rect 200259 140147 200287 140175
rect 200321 140147 200349 140175
rect 200259 140085 200287 140113
rect 200321 140085 200349 140113
rect 200259 140023 200287 140051
rect 200321 140023 200349 140051
rect 200259 139961 200287 139989
rect 200321 139961 200349 139989
rect 192579 137147 192607 137175
rect 192641 137147 192669 137175
rect 192579 137085 192607 137113
rect 192641 137085 192669 137113
rect 192579 137023 192607 137051
rect 192641 137023 192669 137051
rect 192579 136961 192607 136989
rect 192641 136961 192669 136989
rect 202437 137147 202465 137175
rect 202499 137147 202527 137175
rect 202561 137147 202589 137175
rect 202623 137147 202651 137175
rect 202437 137085 202465 137113
rect 202499 137085 202527 137113
rect 202561 137085 202589 137113
rect 202623 137085 202651 137113
rect 202437 137023 202465 137051
rect 202499 137023 202527 137051
rect 202561 137023 202589 137051
rect 202623 137023 202651 137051
rect 202437 136961 202465 136989
rect 202499 136961 202527 136989
rect 202561 136961 202589 136989
rect 202623 136961 202651 136989
rect 188937 131147 188965 131175
rect 188999 131147 189027 131175
rect 189061 131147 189089 131175
rect 189123 131147 189151 131175
rect 188937 131085 188965 131113
rect 188999 131085 189027 131113
rect 189061 131085 189089 131113
rect 189123 131085 189151 131113
rect 188937 131023 188965 131051
rect 188999 131023 189027 131051
rect 189061 131023 189089 131051
rect 189123 131023 189151 131051
rect 188937 130961 188965 130989
rect 188999 130961 189027 130989
rect 189061 130961 189089 130989
rect 189123 130961 189151 130989
rect 200259 131147 200287 131175
rect 200321 131147 200349 131175
rect 200259 131085 200287 131113
rect 200321 131085 200349 131113
rect 200259 131023 200287 131051
rect 200321 131023 200349 131051
rect 200259 130961 200287 130989
rect 200321 130961 200349 130989
rect 192579 128147 192607 128175
rect 192641 128147 192669 128175
rect 192579 128085 192607 128113
rect 192641 128085 192669 128113
rect 192579 128023 192607 128051
rect 192641 128023 192669 128051
rect 192579 127961 192607 127989
rect 192641 127961 192669 127989
rect 202437 128147 202465 128175
rect 202499 128147 202527 128175
rect 202561 128147 202589 128175
rect 202623 128147 202651 128175
rect 202437 128085 202465 128113
rect 202499 128085 202527 128113
rect 202561 128085 202589 128113
rect 202623 128085 202651 128113
rect 202437 128023 202465 128051
rect 202499 128023 202527 128051
rect 202561 128023 202589 128051
rect 202623 128023 202651 128051
rect 202437 127961 202465 127989
rect 202499 127961 202527 127989
rect 202561 127961 202589 127989
rect 202623 127961 202651 127989
rect 188937 122147 188965 122175
rect 188999 122147 189027 122175
rect 189061 122147 189089 122175
rect 189123 122147 189151 122175
rect 188937 122085 188965 122113
rect 188999 122085 189027 122113
rect 189061 122085 189089 122113
rect 189123 122085 189151 122113
rect 188937 122023 188965 122051
rect 188999 122023 189027 122051
rect 189061 122023 189089 122051
rect 189123 122023 189151 122051
rect 188937 121961 188965 121989
rect 188999 121961 189027 121989
rect 189061 121961 189089 121989
rect 189123 121961 189151 121989
rect 200259 122147 200287 122175
rect 200321 122147 200349 122175
rect 200259 122085 200287 122113
rect 200321 122085 200349 122113
rect 200259 122023 200287 122051
rect 200321 122023 200349 122051
rect 200259 121961 200287 121989
rect 200321 121961 200349 121989
rect 192579 119147 192607 119175
rect 192641 119147 192669 119175
rect 192579 119085 192607 119113
rect 192641 119085 192669 119113
rect 192579 119023 192607 119051
rect 192641 119023 192669 119051
rect 192579 118961 192607 118989
rect 192641 118961 192669 118989
rect 202437 119147 202465 119175
rect 202499 119147 202527 119175
rect 202561 119147 202589 119175
rect 202623 119147 202651 119175
rect 202437 119085 202465 119113
rect 202499 119085 202527 119113
rect 202561 119085 202589 119113
rect 202623 119085 202651 119113
rect 202437 119023 202465 119051
rect 202499 119023 202527 119051
rect 202561 119023 202589 119051
rect 202623 119023 202651 119051
rect 202437 118961 202465 118989
rect 202499 118961 202527 118989
rect 202561 118961 202589 118989
rect 202623 118961 202651 118989
rect 188937 113147 188965 113175
rect 188999 113147 189027 113175
rect 189061 113147 189089 113175
rect 189123 113147 189151 113175
rect 188937 113085 188965 113113
rect 188999 113085 189027 113113
rect 189061 113085 189089 113113
rect 189123 113085 189151 113113
rect 188937 113023 188965 113051
rect 188999 113023 189027 113051
rect 189061 113023 189089 113051
rect 189123 113023 189151 113051
rect 188937 112961 188965 112989
rect 188999 112961 189027 112989
rect 189061 112961 189089 112989
rect 189123 112961 189151 112989
rect 200259 113147 200287 113175
rect 200321 113147 200349 113175
rect 200259 113085 200287 113113
rect 200321 113085 200349 113113
rect 200259 113023 200287 113051
rect 200321 113023 200349 113051
rect 200259 112961 200287 112989
rect 200321 112961 200349 112989
rect 192579 110147 192607 110175
rect 192641 110147 192669 110175
rect 192579 110085 192607 110113
rect 192641 110085 192669 110113
rect 192579 110023 192607 110051
rect 192641 110023 192669 110051
rect 192579 109961 192607 109989
rect 192641 109961 192669 109989
rect 202437 110147 202465 110175
rect 202499 110147 202527 110175
rect 202561 110147 202589 110175
rect 202623 110147 202651 110175
rect 202437 110085 202465 110113
rect 202499 110085 202527 110113
rect 202561 110085 202589 110113
rect 202623 110085 202651 110113
rect 202437 110023 202465 110051
rect 202499 110023 202527 110051
rect 202561 110023 202589 110051
rect 202623 110023 202651 110051
rect 202437 109961 202465 109989
rect 202499 109961 202527 109989
rect 202561 109961 202589 109989
rect 202623 109961 202651 109989
rect 188937 104147 188965 104175
rect 188999 104147 189027 104175
rect 189061 104147 189089 104175
rect 189123 104147 189151 104175
rect 188937 104085 188965 104113
rect 188999 104085 189027 104113
rect 189061 104085 189089 104113
rect 189123 104085 189151 104113
rect 188937 104023 188965 104051
rect 188999 104023 189027 104051
rect 189061 104023 189089 104051
rect 189123 104023 189151 104051
rect 188937 103961 188965 103989
rect 188999 103961 189027 103989
rect 189061 103961 189089 103989
rect 189123 103961 189151 103989
rect 200259 104147 200287 104175
rect 200321 104147 200349 104175
rect 200259 104085 200287 104113
rect 200321 104085 200349 104113
rect 200259 104023 200287 104051
rect 200321 104023 200349 104051
rect 200259 103961 200287 103989
rect 200321 103961 200349 103989
rect 192579 101147 192607 101175
rect 192641 101147 192669 101175
rect 192579 101085 192607 101113
rect 192641 101085 192669 101113
rect 192579 101023 192607 101051
rect 192641 101023 192669 101051
rect 192579 100961 192607 100989
rect 192641 100961 192669 100989
rect 202437 101147 202465 101175
rect 202499 101147 202527 101175
rect 202561 101147 202589 101175
rect 202623 101147 202651 101175
rect 202437 101085 202465 101113
rect 202499 101085 202527 101113
rect 202561 101085 202589 101113
rect 202623 101085 202651 101113
rect 202437 101023 202465 101051
rect 202499 101023 202527 101051
rect 202561 101023 202589 101051
rect 202623 101023 202651 101051
rect 202437 100961 202465 100989
rect 202499 100961 202527 100989
rect 202561 100961 202589 100989
rect 202623 100961 202651 100989
rect 188937 95147 188965 95175
rect 188999 95147 189027 95175
rect 189061 95147 189089 95175
rect 189123 95147 189151 95175
rect 188937 95085 188965 95113
rect 188999 95085 189027 95113
rect 189061 95085 189089 95113
rect 189123 95085 189151 95113
rect 188937 95023 188965 95051
rect 188999 95023 189027 95051
rect 189061 95023 189089 95051
rect 189123 95023 189151 95051
rect 188937 94961 188965 94989
rect 188999 94961 189027 94989
rect 189061 94961 189089 94989
rect 189123 94961 189151 94989
rect 200259 95147 200287 95175
rect 200321 95147 200349 95175
rect 200259 95085 200287 95113
rect 200321 95085 200349 95113
rect 200259 95023 200287 95051
rect 200321 95023 200349 95051
rect 200259 94961 200287 94989
rect 200321 94961 200349 94989
rect 192579 92147 192607 92175
rect 192641 92147 192669 92175
rect 192579 92085 192607 92113
rect 192641 92085 192669 92113
rect 192579 92023 192607 92051
rect 192641 92023 192669 92051
rect 192579 91961 192607 91989
rect 192641 91961 192669 91989
rect 202437 92147 202465 92175
rect 202499 92147 202527 92175
rect 202561 92147 202589 92175
rect 202623 92147 202651 92175
rect 202437 92085 202465 92113
rect 202499 92085 202527 92113
rect 202561 92085 202589 92113
rect 202623 92085 202651 92113
rect 202437 92023 202465 92051
rect 202499 92023 202527 92051
rect 202561 92023 202589 92051
rect 202623 92023 202651 92051
rect 202437 91961 202465 91989
rect 202499 91961 202527 91989
rect 202561 91961 202589 91989
rect 202623 91961 202651 91989
rect 188937 86147 188965 86175
rect 188999 86147 189027 86175
rect 189061 86147 189089 86175
rect 189123 86147 189151 86175
rect 188937 86085 188965 86113
rect 188999 86085 189027 86113
rect 189061 86085 189089 86113
rect 189123 86085 189151 86113
rect 188937 86023 188965 86051
rect 188999 86023 189027 86051
rect 189061 86023 189089 86051
rect 189123 86023 189151 86051
rect 188937 85961 188965 85989
rect 188999 85961 189027 85989
rect 189061 85961 189089 85989
rect 189123 85961 189151 85989
rect 200259 86147 200287 86175
rect 200321 86147 200349 86175
rect 200259 86085 200287 86113
rect 200321 86085 200349 86113
rect 200259 86023 200287 86051
rect 200321 86023 200349 86051
rect 200259 85961 200287 85989
rect 200321 85961 200349 85989
rect 192579 83147 192607 83175
rect 192641 83147 192669 83175
rect 192579 83085 192607 83113
rect 192641 83085 192669 83113
rect 192579 83023 192607 83051
rect 192641 83023 192669 83051
rect 192579 82961 192607 82989
rect 192641 82961 192669 82989
rect 202437 83147 202465 83175
rect 202499 83147 202527 83175
rect 202561 83147 202589 83175
rect 202623 83147 202651 83175
rect 202437 83085 202465 83113
rect 202499 83085 202527 83113
rect 202561 83085 202589 83113
rect 202623 83085 202651 83113
rect 202437 83023 202465 83051
rect 202499 83023 202527 83051
rect 202561 83023 202589 83051
rect 202623 83023 202651 83051
rect 202437 82961 202465 82989
rect 202499 82961 202527 82989
rect 202561 82961 202589 82989
rect 202623 82961 202651 82989
rect 188937 77147 188965 77175
rect 188999 77147 189027 77175
rect 189061 77147 189089 77175
rect 189123 77147 189151 77175
rect 188937 77085 188965 77113
rect 188999 77085 189027 77113
rect 189061 77085 189089 77113
rect 189123 77085 189151 77113
rect 188937 77023 188965 77051
rect 188999 77023 189027 77051
rect 189061 77023 189089 77051
rect 189123 77023 189151 77051
rect 188937 76961 188965 76989
rect 188999 76961 189027 76989
rect 189061 76961 189089 76989
rect 189123 76961 189151 76989
rect 200259 77147 200287 77175
rect 200321 77147 200349 77175
rect 200259 77085 200287 77113
rect 200321 77085 200349 77113
rect 200259 77023 200287 77051
rect 200321 77023 200349 77051
rect 200259 76961 200287 76989
rect 200321 76961 200349 76989
rect 192579 74147 192607 74175
rect 192641 74147 192669 74175
rect 192579 74085 192607 74113
rect 192641 74085 192669 74113
rect 192579 74023 192607 74051
rect 192641 74023 192669 74051
rect 192579 73961 192607 73989
rect 192641 73961 192669 73989
rect 202437 74147 202465 74175
rect 202499 74147 202527 74175
rect 202561 74147 202589 74175
rect 202623 74147 202651 74175
rect 202437 74085 202465 74113
rect 202499 74085 202527 74113
rect 202561 74085 202589 74113
rect 202623 74085 202651 74113
rect 202437 74023 202465 74051
rect 202499 74023 202527 74051
rect 202561 74023 202589 74051
rect 202623 74023 202651 74051
rect 202437 73961 202465 73989
rect 202499 73961 202527 73989
rect 202561 73961 202589 73989
rect 202623 73961 202651 73989
rect 188937 68147 188965 68175
rect 188999 68147 189027 68175
rect 189061 68147 189089 68175
rect 189123 68147 189151 68175
rect 188937 68085 188965 68113
rect 188999 68085 189027 68113
rect 189061 68085 189089 68113
rect 189123 68085 189151 68113
rect 188937 68023 188965 68051
rect 188999 68023 189027 68051
rect 189061 68023 189089 68051
rect 189123 68023 189151 68051
rect 188937 67961 188965 67989
rect 188999 67961 189027 67989
rect 189061 67961 189089 67989
rect 189123 67961 189151 67989
rect 200259 68147 200287 68175
rect 200321 68147 200349 68175
rect 200259 68085 200287 68113
rect 200321 68085 200349 68113
rect 200259 68023 200287 68051
rect 200321 68023 200349 68051
rect 200259 67961 200287 67989
rect 200321 67961 200349 67989
rect 192579 65147 192607 65175
rect 192641 65147 192669 65175
rect 192579 65085 192607 65113
rect 192641 65085 192669 65113
rect 192579 65023 192607 65051
rect 192641 65023 192669 65051
rect 192579 64961 192607 64989
rect 192641 64961 192669 64989
rect 202437 65147 202465 65175
rect 202499 65147 202527 65175
rect 202561 65147 202589 65175
rect 202623 65147 202651 65175
rect 202437 65085 202465 65113
rect 202499 65085 202527 65113
rect 202561 65085 202589 65113
rect 202623 65085 202651 65113
rect 202437 65023 202465 65051
rect 202499 65023 202527 65051
rect 202561 65023 202589 65051
rect 202623 65023 202651 65051
rect 202437 64961 202465 64989
rect 202499 64961 202527 64989
rect 202561 64961 202589 64989
rect 202623 64961 202651 64989
rect 188937 59147 188965 59175
rect 188999 59147 189027 59175
rect 189061 59147 189089 59175
rect 189123 59147 189151 59175
rect 188937 59085 188965 59113
rect 188999 59085 189027 59113
rect 189061 59085 189089 59113
rect 189123 59085 189151 59113
rect 188937 59023 188965 59051
rect 188999 59023 189027 59051
rect 189061 59023 189089 59051
rect 189123 59023 189151 59051
rect 188937 58961 188965 58989
rect 188999 58961 189027 58989
rect 189061 58961 189089 58989
rect 189123 58961 189151 58989
rect 200259 59147 200287 59175
rect 200321 59147 200349 59175
rect 200259 59085 200287 59113
rect 200321 59085 200349 59113
rect 200259 59023 200287 59051
rect 200321 59023 200349 59051
rect 200259 58961 200287 58989
rect 200321 58961 200349 58989
rect 192579 56147 192607 56175
rect 192641 56147 192669 56175
rect 192579 56085 192607 56113
rect 192641 56085 192669 56113
rect 192579 56023 192607 56051
rect 192641 56023 192669 56051
rect 192579 55961 192607 55989
rect 192641 55961 192669 55989
rect 202437 56147 202465 56175
rect 202499 56147 202527 56175
rect 202561 56147 202589 56175
rect 202623 56147 202651 56175
rect 202437 56085 202465 56113
rect 202499 56085 202527 56113
rect 202561 56085 202589 56113
rect 202623 56085 202651 56113
rect 202437 56023 202465 56051
rect 202499 56023 202527 56051
rect 202561 56023 202589 56051
rect 202623 56023 202651 56051
rect 202437 55961 202465 55989
rect 202499 55961 202527 55989
rect 202561 55961 202589 55989
rect 202623 55961 202651 55989
rect 188937 50147 188965 50175
rect 188999 50147 189027 50175
rect 189061 50147 189089 50175
rect 189123 50147 189151 50175
rect 188937 50085 188965 50113
rect 188999 50085 189027 50113
rect 189061 50085 189089 50113
rect 189123 50085 189151 50113
rect 188937 50023 188965 50051
rect 188999 50023 189027 50051
rect 189061 50023 189089 50051
rect 189123 50023 189151 50051
rect 188937 49961 188965 49989
rect 188999 49961 189027 49989
rect 189061 49961 189089 49989
rect 189123 49961 189151 49989
rect 200259 50147 200287 50175
rect 200321 50147 200349 50175
rect 200259 50085 200287 50113
rect 200321 50085 200349 50113
rect 200259 50023 200287 50051
rect 200321 50023 200349 50051
rect 200259 49961 200287 49989
rect 200321 49961 200349 49989
rect 192579 47147 192607 47175
rect 192641 47147 192669 47175
rect 192579 47085 192607 47113
rect 192641 47085 192669 47113
rect 192579 47023 192607 47051
rect 192641 47023 192669 47051
rect 192579 46961 192607 46989
rect 192641 46961 192669 46989
rect 202437 47147 202465 47175
rect 202499 47147 202527 47175
rect 202561 47147 202589 47175
rect 202623 47147 202651 47175
rect 202437 47085 202465 47113
rect 202499 47085 202527 47113
rect 202561 47085 202589 47113
rect 202623 47085 202651 47113
rect 202437 47023 202465 47051
rect 202499 47023 202527 47051
rect 202561 47023 202589 47051
rect 202623 47023 202651 47051
rect 202437 46961 202465 46989
rect 202499 46961 202527 46989
rect 202561 46961 202589 46989
rect 202623 46961 202651 46989
rect 188937 41147 188965 41175
rect 188999 41147 189027 41175
rect 189061 41147 189089 41175
rect 189123 41147 189151 41175
rect 188937 41085 188965 41113
rect 188999 41085 189027 41113
rect 189061 41085 189089 41113
rect 189123 41085 189151 41113
rect 188937 41023 188965 41051
rect 188999 41023 189027 41051
rect 189061 41023 189089 41051
rect 189123 41023 189151 41051
rect 188937 40961 188965 40989
rect 188999 40961 189027 40989
rect 189061 40961 189089 40989
rect 189123 40961 189151 40989
rect 200259 41147 200287 41175
rect 200321 41147 200349 41175
rect 200259 41085 200287 41113
rect 200321 41085 200349 41113
rect 200259 41023 200287 41051
rect 200321 41023 200349 41051
rect 200259 40961 200287 40989
rect 200321 40961 200349 40989
rect 192579 38147 192607 38175
rect 192641 38147 192669 38175
rect 192579 38085 192607 38113
rect 192641 38085 192669 38113
rect 192579 38023 192607 38051
rect 192641 38023 192669 38051
rect 192579 37961 192607 37989
rect 192641 37961 192669 37989
rect 202437 38147 202465 38175
rect 202499 38147 202527 38175
rect 202561 38147 202589 38175
rect 202623 38147 202651 38175
rect 202437 38085 202465 38113
rect 202499 38085 202527 38113
rect 202561 38085 202589 38113
rect 202623 38085 202651 38113
rect 202437 38023 202465 38051
rect 202499 38023 202527 38051
rect 202561 38023 202589 38051
rect 202623 38023 202651 38051
rect 202437 37961 202465 37989
rect 202499 37961 202527 37989
rect 202561 37961 202589 37989
rect 202623 37961 202651 37989
rect 188937 32147 188965 32175
rect 188999 32147 189027 32175
rect 189061 32147 189089 32175
rect 189123 32147 189151 32175
rect 188937 32085 188965 32113
rect 188999 32085 189027 32113
rect 189061 32085 189089 32113
rect 189123 32085 189151 32113
rect 188937 32023 188965 32051
rect 188999 32023 189027 32051
rect 189061 32023 189089 32051
rect 189123 32023 189151 32051
rect 188937 31961 188965 31989
rect 188999 31961 189027 31989
rect 189061 31961 189089 31989
rect 189123 31961 189151 31989
rect 200259 32147 200287 32175
rect 200321 32147 200349 32175
rect 200259 32085 200287 32113
rect 200321 32085 200349 32113
rect 200259 32023 200287 32051
rect 200321 32023 200349 32051
rect 200259 31961 200287 31989
rect 200321 31961 200349 31989
rect 192579 29147 192607 29175
rect 192641 29147 192669 29175
rect 192579 29085 192607 29113
rect 192641 29085 192669 29113
rect 192579 29023 192607 29051
rect 192641 29023 192669 29051
rect 192579 28961 192607 28989
rect 192641 28961 192669 28989
rect 202437 29147 202465 29175
rect 202499 29147 202527 29175
rect 202561 29147 202589 29175
rect 202623 29147 202651 29175
rect 202437 29085 202465 29113
rect 202499 29085 202527 29113
rect 202561 29085 202589 29113
rect 202623 29085 202651 29113
rect 202437 29023 202465 29051
rect 202499 29023 202527 29051
rect 202561 29023 202589 29051
rect 202623 29023 202651 29051
rect 202437 28961 202465 28989
rect 202499 28961 202527 28989
rect 202561 28961 202589 28989
rect 202623 28961 202651 28989
rect 188937 23147 188965 23175
rect 188999 23147 189027 23175
rect 189061 23147 189089 23175
rect 189123 23147 189151 23175
rect 188937 23085 188965 23113
rect 188999 23085 189027 23113
rect 189061 23085 189089 23113
rect 189123 23085 189151 23113
rect 188937 23023 188965 23051
rect 188999 23023 189027 23051
rect 189061 23023 189089 23051
rect 189123 23023 189151 23051
rect 188937 22961 188965 22989
rect 188999 22961 189027 22989
rect 189061 22961 189089 22989
rect 189123 22961 189151 22989
rect 200259 23147 200287 23175
rect 200321 23147 200349 23175
rect 200259 23085 200287 23113
rect 200321 23085 200349 23113
rect 200259 23023 200287 23051
rect 200321 23023 200349 23051
rect 200259 22961 200287 22989
rect 200321 22961 200349 22989
rect 192579 20147 192607 20175
rect 192641 20147 192669 20175
rect 192579 20085 192607 20113
rect 192641 20085 192669 20113
rect 192579 20023 192607 20051
rect 192641 20023 192669 20051
rect 192579 19961 192607 19989
rect 192641 19961 192669 19989
rect 202437 20147 202465 20175
rect 202499 20147 202527 20175
rect 202561 20147 202589 20175
rect 202623 20147 202651 20175
rect 202437 20085 202465 20113
rect 202499 20085 202527 20113
rect 202561 20085 202589 20113
rect 202623 20085 202651 20113
rect 202437 20023 202465 20051
rect 202499 20023 202527 20051
rect 202561 20023 202589 20051
rect 202623 20023 202651 20051
rect 202437 19961 202465 19989
rect 202499 19961 202527 19989
rect 202561 19961 202589 19989
rect 202623 19961 202651 19989
rect 188937 14147 188965 14175
rect 188999 14147 189027 14175
rect 189061 14147 189089 14175
rect 189123 14147 189151 14175
rect 188937 14085 188965 14113
rect 188999 14085 189027 14113
rect 189061 14085 189089 14113
rect 189123 14085 189151 14113
rect 188937 14023 188965 14051
rect 188999 14023 189027 14051
rect 189061 14023 189089 14051
rect 189123 14023 189151 14051
rect 188937 13961 188965 13989
rect 188999 13961 189027 13989
rect 189061 13961 189089 13989
rect 189123 13961 189151 13989
rect 200259 14147 200287 14175
rect 200321 14147 200349 14175
rect 200259 14085 200287 14113
rect 200321 14085 200349 14113
rect 200259 14023 200287 14051
rect 200321 14023 200349 14051
rect 200259 13961 200287 13989
rect 200321 13961 200349 13989
rect 192579 11147 192607 11175
rect 192641 11147 192669 11175
rect 192579 11085 192607 11113
rect 192641 11085 192669 11113
rect 192579 11023 192607 11051
rect 192641 11023 192669 11051
rect 192579 10961 192607 10989
rect 192641 10961 192669 10989
rect 202437 11147 202465 11175
rect 202499 11147 202527 11175
rect 202561 11147 202589 11175
rect 202623 11147 202651 11175
rect 202437 11085 202465 11113
rect 202499 11085 202527 11113
rect 202561 11085 202589 11113
rect 202623 11085 202651 11113
rect 202437 11023 202465 11051
rect 202499 11023 202527 11051
rect 202561 11023 202589 11051
rect 202623 11023 202651 11051
rect 202437 10961 202465 10989
rect 202499 10961 202527 10989
rect 202561 10961 202589 10989
rect 202623 10961 202651 10989
rect 188937 5147 188965 5175
rect 188999 5147 189027 5175
rect 189061 5147 189089 5175
rect 189123 5147 189151 5175
rect 188937 5085 188965 5113
rect 188999 5085 189027 5113
rect 189061 5085 189089 5113
rect 189123 5085 189151 5113
rect 188937 5023 188965 5051
rect 188999 5023 189027 5051
rect 189061 5023 189089 5051
rect 189123 5023 189151 5051
rect 188937 4961 188965 4989
rect 188999 4961 189027 4989
rect 189061 4961 189089 4989
rect 189123 4961 189151 4989
rect 200259 5147 200287 5175
rect 200321 5147 200349 5175
rect 200259 5085 200287 5113
rect 200321 5085 200349 5113
rect 200259 5023 200287 5051
rect 200321 5023 200349 5051
rect 200259 4961 200287 4989
rect 200321 4961 200349 4989
rect 188937 -588 188965 -560
rect 188999 -588 189027 -560
rect 189061 -588 189089 -560
rect 189123 -588 189151 -560
rect 188937 -650 188965 -622
rect 188999 -650 189027 -622
rect 189061 -650 189089 -622
rect 189123 -650 189151 -622
rect 188937 -712 188965 -684
rect 188999 -712 189027 -684
rect 189061 -712 189089 -684
rect 189123 -712 189151 -684
rect 188937 -774 188965 -746
rect 188999 -774 189027 -746
rect 189061 -774 189089 -746
rect 189123 -774 189151 -746
rect 202437 2147 202465 2175
rect 202499 2147 202527 2175
rect 202561 2147 202589 2175
rect 202623 2147 202651 2175
rect 202437 2085 202465 2113
rect 202499 2085 202527 2113
rect 202561 2085 202589 2113
rect 202623 2085 202651 2113
rect 202437 2023 202465 2051
rect 202499 2023 202527 2051
rect 202561 2023 202589 2051
rect 202623 2023 202651 2051
rect 202437 1961 202465 1989
rect 202499 1961 202527 1989
rect 202561 1961 202589 1989
rect 202623 1961 202651 1989
rect 202437 -108 202465 -80
rect 202499 -108 202527 -80
rect 202561 -108 202589 -80
rect 202623 -108 202651 -80
rect 202437 -170 202465 -142
rect 202499 -170 202527 -142
rect 202561 -170 202589 -142
rect 202623 -170 202651 -142
rect 202437 -232 202465 -204
rect 202499 -232 202527 -204
rect 202561 -232 202589 -204
rect 202623 -232 202651 -204
rect 202437 -294 202465 -266
rect 202499 -294 202527 -266
rect 202561 -294 202589 -266
rect 202623 -294 202651 -266
rect 204297 299058 204325 299086
rect 204359 299058 204387 299086
rect 204421 299058 204449 299086
rect 204483 299058 204511 299086
rect 204297 298996 204325 299024
rect 204359 298996 204387 299024
rect 204421 298996 204449 299024
rect 204483 298996 204511 299024
rect 204297 298934 204325 298962
rect 204359 298934 204387 298962
rect 204421 298934 204449 298962
rect 204483 298934 204511 298962
rect 204297 298872 204325 298900
rect 204359 298872 204387 298900
rect 204421 298872 204449 298900
rect 204483 298872 204511 298900
rect 204297 293147 204325 293175
rect 204359 293147 204387 293175
rect 204421 293147 204449 293175
rect 204483 293147 204511 293175
rect 204297 293085 204325 293113
rect 204359 293085 204387 293113
rect 204421 293085 204449 293113
rect 204483 293085 204511 293113
rect 204297 293023 204325 293051
rect 204359 293023 204387 293051
rect 204421 293023 204449 293051
rect 204483 293023 204511 293051
rect 204297 292961 204325 292989
rect 204359 292961 204387 292989
rect 204421 292961 204449 292989
rect 204483 292961 204511 292989
rect 204297 284147 204325 284175
rect 204359 284147 204387 284175
rect 204421 284147 204449 284175
rect 204483 284147 204511 284175
rect 204297 284085 204325 284113
rect 204359 284085 204387 284113
rect 204421 284085 204449 284113
rect 204483 284085 204511 284113
rect 204297 284023 204325 284051
rect 204359 284023 204387 284051
rect 204421 284023 204449 284051
rect 204483 284023 204511 284051
rect 204297 283961 204325 283989
rect 204359 283961 204387 283989
rect 204421 283961 204449 283989
rect 204483 283961 204511 283989
rect 204297 275147 204325 275175
rect 204359 275147 204387 275175
rect 204421 275147 204449 275175
rect 204483 275147 204511 275175
rect 204297 275085 204325 275113
rect 204359 275085 204387 275113
rect 204421 275085 204449 275113
rect 204483 275085 204511 275113
rect 204297 275023 204325 275051
rect 204359 275023 204387 275051
rect 204421 275023 204449 275051
rect 204483 275023 204511 275051
rect 204297 274961 204325 274989
rect 204359 274961 204387 274989
rect 204421 274961 204449 274989
rect 204483 274961 204511 274989
rect 204297 266147 204325 266175
rect 204359 266147 204387 266175
rect 204421 266147 204449 266175
rect 204483 266147 204511 266175
rect 204297 266085 204325 266113
rect 204359 266085 204387 266113
rect 204421 266085 204449 266113
rect 204483 266085 204511 266113
rect 204297 266023 204325 266051
rect 204359 266023 204387 266051
rect 204421 266023 204449 266051
rect 204483 266023 204511 266051
rect 204297 265961 204325 265989
rect 204359 265961 204387 265989
rect 204421 265961 204449 265989
rect 204483 265961 204511 265989
rect 204297 257147 204325 257175
rect 204359 257147 204387 257175
rect 204421 257147 204449 257175
rect 204483 257147 204511 257175
rect 204297 257085 204325 257113
rect 204359 257085 204387 257113
rect 204421 257085 204449 257113
rect 204483 257085 204511 257113
rect 204297 257023 204325 257051
rect 204359 257023 204387 257051
rect 204421 257023 204449 257051
rect 204483 257023 204511 257051
rect 204297 256961 204325 256989
rect 204359 256961 204387 256989
rect 204421 256961 204449 256989
rect 204483 256961 204511 256989
rect 204297 248147 204325 248175
rect 204359 248147 204387 248175
rect 204421 248147 204449 248175
rect 204483 248147 204511 248175
rect 204297 248085 204325 248113
rect 204359 248085 204387 248113
rect 204421 248085 204449 248113
rect 204483 248085 204511 248113
rect 204297 248023 204325 248051
rect 204359 248023 204387 248051
rect 204421 248023 204449 248051
rect 204483 248023 204511 248051
rect 204297 247961 204325 247989
rect 204359 247961 204387 247989
rect 204421 247961 204449 247989
rect 204483 247961 204511 247989
rect 204297 239147 204325 239175
rect 204359 239147 204387 239175
rect 204421 239147 204449 239175
rect 204483 239147 204511 239175
rect 204297 239085 204325 239113
rect 204359 239085 204387 239113
rect 204421 239085 204449 239113
rect 204483 239085 204511 239113
rect 204297 239023 204325 239051
rect 204359 239023 204387 239051
rect 204421 239023 204449 239051
rect 204483 239023 204511 239051
rect 204297 238961 204325 238989
rect 204359 238961 204387 238989
rect 204421 238961 204449 238989
rect 204483 238961 204511 238989
rect 204297 230147 204325 230175
rect 204359 230147 204387 230175
rect 204421 230147 204449 230175
rect 204483 230147 204511 230175
rect 204297 230085 204325 230113
rect 204359 230085 204387 230113
rect 204421 230085 204449 230113
rect 204483 230085 204511 230113
rect 204297 230023 204325 230051
rect 204359 230023 204387 230051
rect 204421 230023 204449 230051
rect 204483 230023 204511 230051
rect 204297 229961 204325 229989
rect 204359 229961 204387 229989
rect 204421 229961 204449 229989
rect 204483 229961 204511 229989
rect 204297 221147 204325 221175
rect 204359 221147 204387 221175
rect 204421 221147 204449 221175
rect 204483 221147 204511 221175
rect 204297 221085 204325 221113
rect 204359 221085 204387 221113
rect 204421 221085 204449 221113
rect 204483 221085 204511 221113
rect 204297 221023 204325 221051
rect 204359 221023 204387 221051
rect 204421 221023 204449 221051
rect 204483 221023 204511 221051
rect 204297 220961 204325 220989
rect 204359 220961 204387 220989
rect 204421 220961 204449 220989
rect 204483 220961 204511 220989
rect 204297 212147 204325 212175
rect 204359 212147 204387 212175
rect 204421 212147 204449 212175
rect 204483 212147 204511 212175
rect 204297 212085 204325 212113
rect 204359 212085 204387 212113
rect 204421 212085 204449 212113
rect 204483 212085 204511 212113
rect 204297 212023 204325 212051
rect 204359 212023 204387 212051
rect 204421 212023 204449 212051
rect 204483 212023 204511 212051
rect 204297 211961 204325 211989
rect 204359 211961 204387 211989
rect 204421 211961 204449 211989
rect 204483 211961 204511 211989
rect 204297 203147 204325 203175
rect 204359 203147 204387 203175
rect 204421 203147 204449 203175
rect 204483 203147 204511 203175
rect 204297 203085 204325 203113
rect 204359 203085 204387 203113
rect 204421 203085 204449 203113
rect 204483 203085 204511 203113
rect 204297 203023 204325 203051
rect 204359 203023 204387 203051
rect 204421 203023 204449 203051
rect 204483 203023 204511 203051
rect 204297 202961 204325 202989
rect 204359 202961 204387 202989
rect 204421 202961 204449 202989
rect 204483 202961 204511 202989
rect 204297 194147 204325 194175
rect 204359 194147 204387 194175
rect 204421 194147 204449 194175
rect 204483 194147 204511 194175
rect 204297 194085 204325 194113
rect 204359 194085 204387 194113
rect 204421 194085 204449 194113
rect 204483 194085 204511 194113
rect 204297 194023 204325 194051
rect 204359 194023 204387 194051
rect 204421 194023 204449 194051
rect 204483 194023 204511 194051
rect 204297 193961 204325 193989
rect 204359 193961 204387 193989
rect 204421 193961 204449 193989
rect 204483 193961 204511 193989
rect 204297 185147 204325 185175
rect 204359 185147 204387 185175
rect 204421 185147 204449 185175
rect 204483 185147 204511 185175
rect 204297 185085 204325 185113
rect 204359 185085 204387 185113
rect 204421 185085 204449 185113
rect 204483 185085 204511 185113
rect 204297 185023 204325 185051
rect 204359 185023 204387 185051
rect 204421 185023 204449 185051
rect 204483 185023 204511 185051
rect 204297 184961 204325 184989
rect 204359 184961 204387 184989
rect 204421 184961 204449 184989
rect 204483 184961 204511 184989
rect 204297 176147 204325 176175
rect 204359 176147 204387 176175
rect 204421 176147 204449 176175
rect 204483 176147 204511 176175
rect 204297 176085 204325 176113
rect 204359 176085 204387 176113
rect 204421 176085 204449 176113
rect 204483 176085 204511 176113
rect 204297 176023 204325 176051
rect 204359 176023 204387 176051
rect 204421 176023 204449 176051
rect 204483 176023 204511 176051
rect 204297 175961 204325 175989
rect 204359 175961 204387 175989
rect 204421 175961 204449 175989
rect 204483 175961 204511 175989
rect 217797 298578 217825 298606
rect 217859 298578 217887 298606
rect 217921 298578 217949 298606
rect 217983 298578 218011 298606
rect 217797 298516 217825 298544
rect 217859 298516 217887 298544
rect 217921 298516 217949 298544
rect 217983 298516 218011 298544
rect 217797 298454 217825 298482
rect 217859 298454 217887 298482
rect 217921 298454 217949 298482
rect 217983 298454 218011 298482
rect 217797 298392 217825 298420
rect 217859 298392 217887 298420
rect 217921 298392 217949 298420
rect 217983 298392 218011 298420
rect 217797 290147 217825 290175
rect 217859 290147 217887 290175
rect 217921 290147 217949 290175
rect 217983 290147 218011 290175
rect 217797 290085 217825 290113
rect 217859 290085 217887 290113
rect 217921 290085 217949 290113
rect 217983 290085 218011 290113
rect 217797 290023 217825 290051
rect 217859 290023 217887 290051
rect 217921 290023 217949 290051
rect 217983 290023 218011 290051
rect 217797 289961 217825 289989
rect 217859 289961 217887 289989
rect 217921 289961 217949 289989
rect 217983 289961 218011 289989
rect 217797 281147 217825 281175
rect 217859 281147 217887 281175
rect 217921 281147 217949 281175
rect 217983 281147 218011 281175
rect 217797 281085 217825 281113
rect 217859 281085 217887 281113
rect 217921 281085 217949 281113
rect 217983 281085 218011 281113
rect 217797 281023 217825 281051
rect 217859 281023 217887 281051
rect 217921 281023 217949 281051
rect 217983 281023 218011 281051
rect 217797 280961 217825 280989
rect 217859 280961 217887 280989
rect 217921 280961 217949 280989
rect 217983 280961 218011 280989
rect 217797 272147 217825 272175
rect 217859 272147 217887 272175
rect 217921 272147 217949 272175
rect 217983 272147 218011 272175
rect 217797 272085 217825 272113
rect 217859 272085 217887 272113
rect 217921 272085 217949 272113
rect 217983 272085 218011 272113
rect 217797 272023 217825 272051
rect 217859 272023 217887 272051
rect 217921 272023 217949 272051
rect 217983 272023 218011 272051
rect 217797 271961 217825 271989
rect 217859 271961 217887 271989
rect 217921 271961 217949 271989
rect 217983 271961 218011 271989
rect 217797 263147 217825 263175
rect 217859 263147 217887 263175
rect 217921 263147 217949 263175
rect 217983 263147 218011 263175
rect 217797 263085 217825 263113
rect 217859 263085 217887 263113
rect 217921 263085 217949 263113
rect 217983 263085 218011 263113
rect 217797 263023 217825 263051
rect 217859 263023 217887 263051
rect 217921 263023 217949 263051
rect 217983 263023 218011 263051
rect 217797 262961 217825 262989
rect 217859 262961 217887 262989
rect 217921 262961 217949 262989
rect 217983 262961 218011 262989
rect 217797 254147 217825 254175
rect 217859 254147 217887 254175
rect 217921 254147 217949 254175
rect 217983 254147 218011 254175
rect 217797 254085 217825 254113
rect 217859 254085 217887 254113
rect 217921 254085 217949 254113
rect 217983 254085 218011 254113
rect 217797 254023 217825 254051
rect 217859 254023 217887 254051
rect 217921 254023 217949 254051
rect 217983 254023 218011 254051
rect 217797 253961 217825 253989
rect 217859 253961 217887 253989
rect 217921 253961 217949 253989
rect 217983 253961 218011 253989
rect 217797 245147 217825 245175
rect 217859 245147 217887 245175
rect 217921 245147 217949 245175
rect 217983 245147 218011 245175
rect 217797 245085 217825 245113
rect 217859 245085 217887 245113
rect 217921 245085 217949 245113
rect 217983 245085 218011 245113
rect 217797 245023 217825 245051
rect 217859 245023 217887 245051
rect 217921 245023 217949 245051
rect 217983 245023 218011 245051
rect 217797 244961 217825 244989
rect 217859 244961 217887 244989
rect 217921 244961 217949 244989
rect 217983 244961 218011 244989
rect 217797 236147 217825 236175
rect 217859 236147 217887 236175
rect 217921 236147 217949 236175
rect 217983 236147 218011 236175
rect 217797 236085 217825 236113
rect 217859 236085 217887 236113
rect 217921 236085 217949 236113
rect 217983 236085 218011 236113
rect 217797 236023 217825 236051
rect 217859 236023 217887 236051
rect 217921 236023 217949 236051
rect 217983 236023 218011 236051
rect 217797 235961 217825 235989
rect 217859 235961 217887 235989
rect 217921 235961 217949 235989
rect 217983 235961 218011 235989
rect 217797 227147 217825 227175
rect 217859 227147 217887 227175
rect 217921 227147 217949 227175
rect 217983 227147 218011 227175
rect 217797 227085 217825 227113
rect 217859 227085 217887 227113
rect 217921 227085 217949 227113
rect 217983 227085 218011 227113
rect 217797 227023 217825 227051
rect 217859 227023 217887 227051
rect 217921 227023 217949 227051
rect 217983 227023 218011 227051
rect 217797 226961 217825 226989
rect 217859 226961 217887 226989
rect 217921 226961 217949 226989
rect 217983 226961 218011 226989
rect 217797 218147 217825 218175
rect 217859 218147 217887 218175
rect 217921 218147 217949 218175
rect 217983 218147 218011 218175
rect 217797 218085 217825 218113
rect 217859 218085 217887 218113
rect 217921 218085 217949 218113
rect 217983 218085 218011 218113
rect 217797 218023 217825 218051
rect 217859 218023 217887 218051
rect 217921 218023 217949 218051
rect 217983 218023 218011 218051
rect 217797 217961 217825 217989
rect 217859 217961 217887 217989
rect 217921 217961 217949 217989
rect 217983 217961 218011 217989
rect 217797 209147 217825 209175
rect 217859 209147 217887 209175
rect 217921 209147 217949 209175
rect 217983 209147 218011 209175
rect 217797 209085 217825 209113
rect 217859 209085 217887 209113
rect 217921 209085 217949 209113
rect 217983 209085 218011 209113
rect 217797 209023 217825 209051
rect 217859 209023 217887 209051
rect 217921 209023 217949 209051
rect 217983 209023 218011 209051
rect 217797 208961 217825 208989
rect 217859 208961 217887 208989
rect 217921 208961 217949 208989
rect 217983 208961 218011 208989
rect 217797 200147 217825 200175
rect 217859 200147 217887 200175
rect 217921 200147 217949 200175
rect 217983 200147 218011 200175
rect 217797 200085 217825 200113
rect 217859 200085 217887 200113
rect 217921 200085 217949 200113
rect 217983 200085 218011 200113
rect 217797 200023 217825 200051
rect 217859 200023 217887 200051
rect 217921 200023 217949 200051
rect 217983 200023 218011 200051
rect 217797 199961 217825 199989
rect 217859 199961 217887 199989
rect 217921 199961 217949 199989
rect 217983 199961 218011 199989
rect 217797 191147 217825 191175
rect 217859 191147 217887 191175
rect 217921 191147 217949 191175
rect 217983 191147 218011 191175
rect 217797 191085 217825 191113
rect 217859 191085 217887 191113
rect 217921 191085 217949 191113
rect 217983 191085 218011 191113
rect 217797 191023 217825 191051
rect 217859 191023 217887 191051
rect 217921 191023 217949 191051
rect 217983 191023 218011 191051
rect 217797 190961 217825 190989
rect 217859 190961 217887 190989
rect 217921 190961 217949 190989
rect 217983 190961 218011 190989
rect 217797 182147 217825 182175
rect 217859 182147 217887 182175
rect 217921 182147 217949 182175
rect 217983 182147 218011 182175
rect 217797 182085 217825 182113
rect 217859 182085 217887 182113
rect 217921 182085 217949 182113
rect 217983 182085 218011 182113
rect 217797 182023 217825 182051
rect 217859 182023 217887 182051
rect 217921 182023 217949 182051
rect 217983 182023 218011 182051
rect 217797 181961 217825 181989
rect 217859 181961 217887 181989
rect 217921 181961 217949 181989
rect 217983 181961 218011 181989
rect 207939 173147 207967 173175
rect 208001 173147 208029 173175
rect 207939 173085 207967 173113
rect 208001 173085 208029 173113
rect 207939 173023 207967 173051
rect 208001 173023 208029 173051
rect 207939 172961 207967 172989
rect 208001 172961 208029 172989
rect 217797 173147 217825 173175
rect 217859 173147 217887 173175
rect 217921 173147 217949 173175
rect 217983 173147 218011 173175
rect 217797 173085 217825 173113
rect 217859 173085 217887 173113
rect 217921 173085 217949 173113
rect 217983 173085 218011 173113
rect 217797 173023 217825 173051
rect 217859 173023 217887 173051
rect 217921 173023 217949 173051
rect 217983 173023 218011 173051
rect 217797 172961 217825 172989
rect 217859 172961 217887 172989
rect 217921 172961 217949 172989
rect 217983 172961 218011 172989
rect 204297 167147 204325 167175
rect 204359 167147 204387 167175
rect 204421 167147 204449 167175
rect 204483 167147 204511 167175
rect 204297 167085 204325 167113
rect 204359 167085 204387 167113
rect 204421 167085 204449 167113
rect 204483 167085 204511 167113
rect 204297 167023 204325 167051
rect 204359 167023 204387 167051
rect 204421 167023 204449 167051
rect 204483 167023 204511 167051
rect 204297 166961 204325 166989
rect 204359 166961 204387 166989
rect 204421 166961 204449 166989
rect 204483 166961 204511 166989
rect 215619 167147 215647 167175
rect 215681 167147 215709 167175
rect 215619 167085 215647 167113
rect 215681 167085 215709 167113
rect 215619 167023 215647 167051
rect 215681 167023 215709 167051
rect 215619 166961 215647 166989
rect 215681 166961 215709 166989
rect 207939 164147 207967 164175
rect 208001 164147 208029 164175
rect 207939 164085 207967 164113
rect 208001 164085 208029 164113
rect 207939 164023 207967 164051
rect 208001 164023 208029 164051
rect 207939 163961 207967 163989
rect 208001 163961 208029 163989
rect 217797 164147 217825 164175
rect 217859 164147 217887 164175
rect 217921 164147 217949 164175
rect 217983 164147 218011 164175
rect 217797 164085 217825 164113
rect 217859 164085 217887 164113
rect 217921 164085 217949 164113
rect 217983 164085 218011 164113
rect 217797 164023 217825 164051
rect 217859 164023 217887 164051
rect 217921 164023 217949 164051
rect 217983 164023 218011 164051
rect 217797 163961 217825 163989
rect 217859 163961 217887 163989
rect 217921 163961 217949 163989
rect 217983 163961 218011 163989
rect 204297 158147 204325 158175
rect 204359 158147 204387 158175
rect 204421 158147 204449 158175
rect 204483 158147 204511 158175
rect 204297 158085 204325 158113
rect 204359 158085 204387 158113
rect 204421 158085 204449 158113
rect 204483 158085 204511 158113
rect 204297 158023 204325 158051
rect 204359 158023 204387 158051
rect 204421 158023 204449 158051
rect 204483 158023 204511 158051
rect 204297 157961 204325 157989
rect 204359 157961 204387 157989
rect 204421 157961 204449 157989
rect 204483 157961 204511 157989
rect 215619 158147 215647 158175
rect 215681 158147 215709 158175
rect 215619 158085 215647 158113
rect 215681 158085 215709 158113
rect 215619 158023 215647 158051
rect 215681 158023 215709 158051
rect 215619 157961 215647 157989
rect 215681 157961 215709 157989
rect 207939 155147 207967 155175
rect 208001 155147 208029 155175
rect 207939 155085 207967 155113
rect 208001 155085 208029 155113
rect 207939 155023 207967 155051
rect 208001 155023 208029 155051
rect 207939 154961 207967 154989
rect 208001 154961 208029 154989
rect 217797 155147 217825 155175
rect 217859 155147 217887 155175
rect 217921 155147 217949 155175
rect 217983 155147 218011 155175
rect 217797 155085 217825 155113
rect 217859 155085 217887 155113
rect 217921 155085 217949 155113
rect 217983 155085 218011 155113
rect 217797 155023 217825 155051
rect 217859 155023 217887 155051
rect 217921 155023 217949 155051
rect 217983 155023 218011 155051
rect 217797 154961 217825 154989
rect 217859 154961 217887 154989
rect 217921 154961 217949 154989
rect 217983 154961 218011 154989
rect 204297 149147 204325 149175
rect 204359 149147 204387 149175
rect 204421 149147 204449 149175
rect 204483 149147 204511 149175
rect 204297 149085 204325 149113
rect 204359 149085 204387 149113
rect 204421 149085 204449 149113
rect 204483 149085 204511 149113
rect 204297 149023 204325 149051
rect 204359 149023 204387 149051
rect 204421 149023 204449 149051
rect 204483 149023 204511 149051
rect 204297 148961 204325 148989
rect 204359 148961 204387 148989
rect 204421 148961 204449 148989
rect 204483 148961 204511 148989
rect 215619 149147 215647 149175
rect 215681 149147 215709 149175
rect 215619 149085 215647 149113
rect 215681 149085 215709 149113
rect 215619 149023 215647 149051
rect 215681 149023 215709 149051
rect 215619 148961 215647 148989
rect 215681 148961 215709 148989
rect 207939 146147 207967 146175
rect 208001 146147 208029 146175
rect 207939 146085 207967 146113
rect 208001 146085 208029 146113
rect 207939 146023 207967 146051
rect 208001 146023 208029 146051
rect 207939 145961 207967 145989
rect 208001 145961 208029 145989
rect 217797 146147 217825 146175
rect 217859 146147 217887 146175
rect 217921 146147 217949 146175
rect 217983 146147 218011 146175
rect 217797 146085 217825 146113
rect 217859 146085 217887 146113
rect 217921 146085 217949 146113
rect 217983 146085 218011 146113
rect 217797 146023 217825 146051
rect 217859 146023 217887 146051
rect 217921 146023 217949 146051
rect 217983 146023 218011 146051
rect 217797 145961 217825 145989
rect 217859 145961 217887 145989
rect 217921 145961 217949 145989
rect 217983 145961 218011 145989
rect 204297 140147 204325 140175
rect 204359 140147 204387 140175
rect 204421 140147 204449 140175
rect 204483 140147 204511 140175
rect 204297 140085 204325 140113
rect 204359 140085 204387 140113
rect 204421 140085 204449 140113
rect 204483 140085 204511 140113
rect 204297 140023 204325 140051
rect 204359 140023 204387 140051
rect 204421 140023 204449 140051
rect 204483 140023 204511 140051
rect 204297 139961 204325 139989
rect 204359 139961 204387 139989
rect 204421 139961 204449 139989
rect 204483 139961 204511 139989
rect 215619 140147 215647 140175
rect 215681 140147 215709 140175
rect 215619 140085 215647 140113
rect 215681 140085 215709 140113
rect 215619 140023 215647 140051
rect 215681 140023 215709 140051
rect 215619 139961 215647 139989
rect 215681 139961 215709 139989
rect 207939 137147 207967 137175
rect 208001 137147 208029 137175
rect 207939 137085 207967 137113
rect 208001 137085 208029 137113
rect 207939 137023 207967 137051
rect 208001 137023 208029 137051
rect 207939 136961 207967 136989
rect 208001 136961 208029 136989
rect 217797 137147 217825 137175
rect 217859 137147 217887 137175
rect 217921 137147 217949 137175
rect 217983 137147 218011 137175
rect 217797 137085 217825 137113
rect 217859 137085 217887 137113
rect 217921 137085 217949 137113
rect 217983 137085 218011 137113
rect 217797 137023 217825 137051
rect 217859 137023 217887 137051
rect 217921 137023 217949 137051
rect 217983 137023 218011 137051
rect 217797 136961 217825 136989
rect 217859 136961 217887 136989
rect 217921 136961 217949 136989
rect 217983 136961 218011 136989
rect 204297 131147 204325 131175
rect 204359 131147 204387 131175
rect 204421 131147 204449 131175
rect 204483 131147 204511 131175
rect 204297 131085 204325 131113
rect 204359 131085 204387 131113
rect 204421 131085 204449 131113
rect 204483 131085 204511 131113
rect 204297 131023 204325 131051
rect 204359 131023 204387 131051
rect 204421 131023 204449 131051
rect 204483 131023 204511 131051
rect 204297 130961 204325 130989
rect 204359 130961 204387 130989
rect 204421 130961 204449 130989
rect 204483 130961 204511 130989
rect 215619 131147 215647 131175
rect 215681 131147 215709 131175
rect 215619 131085 215647 131113
rect 215681 131085 215709 131113
rect 215619 131023 215647 131051
rect 215681 131023 215709 131051
rect 215619 130961 215647 130989
rect 215681 130961 215709 130989
rect 207939 128147 207967 128175
rect 208001 128147 208029 128175
rect 207939 128085 207967 128113
rect 208001 128085 208029 128113
rect 207939 128023 207967 128051
rect 208001 128023 208029 128051
rect 207939 127961 207967 127989
rect 208001 127961 208029 127989
rect 217797 128147 217825 128175
rect 217859 128147 217887 128175
rect 217921 128147 217949 128175
rect 217983 128147 218011 128175
rect 217797 128085 217825 128113
rect 217859 128085 217887 128113
rect 217921 128085 217949 128113
rect 217983 128085 218011 128113
rect 217797 128023 217825 128051
rect 217859 128023 217887 128051
rect 217921 128023 217949 128051
rect 217983 128023 218011 128051
rect 217797 127961 217825 127989
rect 217859 127961 217887 127989
rect 217921 127961 217949 127989
rect 217983 127961 218011 127989
rect 204297 122147 204325 122175
rect 204359 122147 204387 122175
rect 204421 122147 204449 122175
rect 204483 122147 204511 122175
rect 204297 122085 204325 122113
rect 204359 122085 204387 122113
rect 204421 122085 204449 122113
rect 204483 122085 204511 122113
rect 204297 122023 204325 122051
rect 204359 122023 204387 122051
rect 204421 122023 204449 122051
rect 204483 122023 204511 122051
rect 204297 121961 204325 121989
rect 204359 121961 204387 121989
rect 204421 121961 204449 121989
rect 204483 121961 204511 121989
rect 215619 122147 215647 122175
rect 215681 122147 215709 122175
rect 215619 122085 215647 122113
rect 215681 122085 215709 122113
rect 215619 122023 215647 122051
rect 215681 122023 215709 122051
rect 215619 121961 215647 121989
rect 215681 121961 215709 121989
rect 207939 119147 207967 119175
rect 208001 119147 208029 119175
rect 207939 119085 207967 119113
rect 208001 119085 208029 119113
rect 207939 119023 207967 119051
rect 208001 119023 208029 119051
rect 207939 118961 207967 118989
rect 208001 118961 208029 118989
rect 217797 119147 217825 119175
rect 217859 119147 217887 119175
rect 217921 119147 217949 119175
rect 217983 119147 218011 119175
rect 217797 119085 217825 119113
rect 217859 119085 217887 119113
rect 217921 119085 217949 119113
rect 217983 119085 218011 119113
rect 217797 119023 217825 119051
rect 217859 119023 217887 119051
rect 217921 119023 217949 119051
rect 217983 119023 218011 119051
rect 217797 118961 217825 118989
rect 217859 118961 217887 118989
rect 217921 118961 217949 118989
rect 217983 118961 218011 118989
rect 204297 113147 204325 113175
rect 204359 113147 204387 113175
rect 204421 113147 204449 113175
rect 204483 113147 204511 113175
rect 204297 113085 204325 113113
rect 204359 113085 204387 113113
rect 204421 113085 204449 113113
rect 204483 113085 204511 113113
rect 204297 113023 204325 113051
rect 204359 113023 204387 113051
rect 204421 113023 204449 113051
rect 204483 113023 204511 113051
rect 204297 112961 204325 112989
rect 204359 112961 204387 112989
rect 204421 112961 204449 112989
rect 204483 112961 204511 112989
rect 215619 113147 215647 113175
rect 215681 113147 215709 113175
rect 215619 113085 215647 113113
rect 215681 113085 215709 113113
rect 215619 113023 215647 113051
rect 215681 113023 215709 113051
rect 215619 112961 215647 112989
rect 215681 112961 215709 112989
rect 207939 110147 207967 110175
rect 208001 110147 208029 110175
rect 207939 110085 207967 110113
rect 208001 110085 208029 110113
rect 207939 110023 207967 110051
rect 208001 110023 208029 110051
rect 207939 109961 207967 109989
rect 208001 109961 208029 109989
rect 217797 110147 217825 110175
rect 217859 110147 217887 110175
rect 217921 110147 217949 110175
rect 217983 110147 218011 110175
rect 217797 110085 217825 110113
rect 217859 110085 217887 110113
rect 217921 110085 217949 110113
rect 217983 110085 218011 110113
rect 217797 110023 217825 110051
rect 217859 110023 217887 110051
rect 217921 110023 217949 110051
rect 217983 110023 218011 110051
rect 217797 109961 217825 109989
rect 217859 109961 217887 109989
rect 217921 109961 217949 109989
rect 217983 109961 218011 109989
rect 204297 104147 204325 104175
rect 204359 104147 204387 104175
rect 204421 104147 204449 104175
rect 204483 104147 204511 104175
rect 204297 104085 204325 104113
rect 204359 104085 204387 104113
rect 204421 104085 204449 104113
rect 204483 104085 204511 104113
rect 204297 104023 204325 104051
rect 204359 104023 204387 104051
rect 204421 104023 204449 104051
rect 204483 104023 204511 104051
rect 204297 103961 204325 103989
rect 204359 103961 204387 103989
rect 204421 103961 204449 103989
rect 204483 103961 204511 103989
rect 215619 104147 215647 104175
rect 215681 104147 215709 104175
rect 215619 104085 215647 104113
rect 215681 104085 215709 104113
rect 215619 104023 215647 104051
rect 215681 104023 215709 104051
rect 215619 103961 215647 103989
rect 215681 103961 215709 103989
rect 207939 101147 207967 101175
rect 208001 101147 208029 101175
rect 207939 101085 207967 101113
rect 208001 101085 208029 101113
rect 207939 101023 207967 101051
rect 208001 101023 208029 101051
rect 207939 100961 207967 100989
rect 208001 100961 208029 100989
rect 217797 101147 217825 101175
rect 217859 101147 217887 101175
rect 217921 101147 217949 101175
rect 217983 101147 218011 101175
rect 217797 101085 217825 101113
rect 217859 101085 217887 101113
rect 217921 101085 217949 101113
rect 217983 101085 218011 101113
rect 217797 101023 217825 101051
rect 217859 101023 217887 101051
rect 217921 101023 217949 101051
rect 217983 101023 218011 101051
rect 217797 100961 217825 100989
rect 217859 100961 217887 100989
rect 217921 100961 217949 100989
rect 217983 100961 218011 100989
rect 204297 95147 204325 95175
rect 204359 95147 204387 95175
rect 204421 95147 204449 95175
rect 204483 95147 204511 95175
rect 204297 95085 204325 95113
rect 204359 95085 204387 95113
rect 204421 95085 204449 95113
rect 204483 95085 204511 95113
rect 204297 95023 204325 95051
rect 204359 95023 204387 95051
rect 204421 95023 204449 95051
rect 204483 95023 204511 95051
rect 204297 94961 204325 94989
rect 204359 94961 204387 94989
rect 204421 94961 204449 94989
rect 204483 94961 204511 94989
rect 215619 95147 215647 95175
rect 215681 95147 215709 95175
rect 215619 95085 215647 95113
rect 215681 95085 215709 95113
rect 215619 95023 215647 95051
rect 215681 95023 215709 95051
rect 215619 94961 215647 94989
rect 215681 94961 215709 94989
rect 207939 92147 207967 92175
rect 208001 92147 208029 92175
rect 207939 92085 207967 92113
rect 208001 92085 208029 92113
rect 207939 92023 207967 92051
rect 208001 92023 208029 92051
rect 207939 91961 207967 91989
rect 208001 91961 208029 91989
rect 217797 92147 217825 92175
rect 217859 92147 217887 92175
rect 217921 92147 217949 92175
rect 217983 92147 218011 92175
rect 217797 92085 217825 92113
rect 217859 92085 217887 92113
rect 217921 92085 217949 92113
rect 217983 92085 218011 92113
rect 217797 92023 217825 92051
rect 217859 92023 217887 92051
rect 217921 92023 217949 92051
rect 217983 92023 218011 92051
rect 217797 91961 217825 91989
rect 217859 91961 217887 91989
rect 217921 91961 217949 91989
rect 217983 91961 218011 91989
rect 204297 86147 204325 86175
rect 204359 86147 204387 86175
rect 204421 86147 204449 86175
rect 204483 86147 204511 86175
rect 204297 86085 204325 86113
rect 204359 86085 204387 86113
rect 204421 86085 204449 86113
rect 204483 86085 204511 86113
rect 204297 86023 204325 86051
rect 204359 86023 204387 86051
rect 204421 86023 204449 86051
rect 204483 86023 204511 86051
rect 204297 85961 204325 85989
rect 204359 85961 204387 85989
rect 204421 85961 204449 85989
rect 204483 85961 204511 85989
rect 215619 86147 215647 86175
rect 215681 86147 215709 86175
rect 215619 86085 215647 86113
rect 215681 86085 215709 86113
rect 215619 86023 215647 86051
rect 215681 86023 215709 86051
rect 215619 85961 215647 85989
rect 215681 85961 215709 85989
rect 207939 83147 207967 83175
rect 208001 83147 208029 83175
rect 207939 83085 207967 83113
rect 208001 83085 208029 83113
rect 207939 83023 207967 83051
rect 208001 83023 208029 83051
rect 207939 82961 207967 82989
rect 208001 82961 208029 82989
rect 217797 83147 217825 83175
rect 217859 83147 217887 83175
rect 217921 83147 217949 83175
rect 217983 83147 218011 83175
rect 217797 83085 217825 83113
rect 217859 83085 217887 83113
rect 217921 83085 217949 83113
rect 217983 83085 218011 83113
rect 217797 83023 217825 83051
rect 217859 83023 217887 83051
rect 217921 83023 217949 83051
rect 217983 83023 218011 83051
rect 217797 82961 217825 82989
rect 217859 82961 217887 82989
rect 217921 82961 217949 82989
rect 217983 82961 218011 82989
rect 204297 77147 204325 77175
rect 204359 77147 204387 77175
rect 204421 77147 204449 77175
rect 204483 77147 204511 77175
rect 204297 77085 204325 77113
rect 204359 77085 204387 77113
rect 204421 77085 204449 77113
rect 204483 77085 204511 77113
rect 204297 77023 204325 77051
rect 204359 77023 204387 77051
rect 204421 77023 204449 77051
rect 204483 77023 204511 77051
rect 204297 76961 204325 76989
rect 204359 76961 204387 76989
rect 204421 76961 204449 76989
rect 204483 76961 204511 76989
rect 215619 77147 215647 77175
rect 215681 77147 215709 77175
rect 215619 77085 215647 77113
rect 215681 77085 215709 77113
rect 215619 77023 215647 77051
rect 215681 77023 215709 77051
rect 215619 76961 215647 76989
rect 215681 76961 215709 76989
rect 207939 74147 207967 74175
rect 208001 74147 208029 74175
rect 207939 74085 207967 74113
rect 208001 74085 208029 74113
rect 207939 74023 207967 74051
rect 208001 74023 208029 74051
rect 207939 73961 207967 73989
rect 208001 73961 208029 73989
rect 217797 74147 217825 74175
rect 217859 74147 217887 74175
rect 217921 74147 217949 74175
rect 217983 74147 218011 74175
rect 217797 74085 217825 74113
rect 217859 74085 217887 74113
rect 217921 74085 217949 74113
rect 217983 74085 218011 74113
rect 217797 74023 217825 74051
rect 217859 74023 217887 74051
rect 217921 74023 217949 74051
rect 217983 74023 218011 74051
rect 217797 73961 217825 73989
rect 217859 73961 217887 73989
rect 217921 73961 217949 73989
rect 217983 73961 218011 73989
rect 204297 68147 204325 68175
rect 204359 68147 204387 68175
rect 204421 68147 204449 68175
rect 204483 68147 204511 68175
rect 204297 68085 204325 68113
rect 204359 68085 204387 68113
rect 204421 68085 204449 68113
rect 204483 68085 204511 68113
rect 204297 68023 204325 68051
rect 204359 68023 204387 68051
rect 204421 68023 204449 68051
rect 204483 68023 204511 68051
rect 204297 67961 204325 67989
rect 204359 67961 204387 67989
rect 204421 67961 204449 67989
rect 204483 67961 204511 67989
rect 215619 68147 215647 68175
rect 215681 68147 215709 68175
rect 215619 68085 215647 68113
rect 215681 68085 215709 68113
rect 215619 68023 215647 68051
rect 215681 68023 215709 68051
rect 215619 67961 215647 67989
rect 215681 67961 215709 67989
rect 207939 65147 207967 65175
rect 208001 65147 208029 65175
rect 207939 65085 207967 65113
rect 208001 65085 208029 65113
rect 207939 65023 207967 65051
rect 208001 65023 208029 65051
rect 207939 64961 207967 64989
rect 208001 64961 208029 64989
rect 217797 65147 217825 65175
rect 217859 65147 217887 65175
rect 217921 65147 217949 65175
rect 217983 65147 218011 65175
rect 217797 65085 217825 65113
rect 217859 65085 217887 65113
rect 217921 65085 217949 65113
rect 217983 65085 218011 65113
rect 217797 65023 217825 65051
rect 217859 65023 217887 65051
rect 217921 65023 217949 65051
rect 217983 65023 218011 65051
rect 217797 64961 217825 64989
rect 217859 64961 217887 64989
rect 217921 64961 217949 64989
rect 217983 64961 218011 64989
rect 204297 59147 204325 59175
rect 204359 59147 204387 59175
rect 204421 59147 204449 59175
rect 204483 59147 204511 59175
rect 204297 59085 204325 59113
rect 204359 59085 204387 59113
rect 204421 59085 204449 59113
rect 204483 59085 204511 59113
rect 204297 59023 204325 59051
rect 204359 59023 204387 59051
rect 204421 59023 204449 59051
rect 204483 59023 204511 59051
rect 204297 58961 204325 58989
rect 204359 58961 204387 58989
rect 204421 58961 204449 58989
rect 204483 58961 204511 58989
rect 215619 59147 215647 59175
rect 215681 59147 215709 59175
rect 215619 59085 215647 59113
rect 215681 59085 215709 59113
rect 215619 59023 215647 59051
rect 215681 59023 215709 59051
rect 215619 58961 215647 58989
rect 215681 58961 215709 58989
rect 207939 56147 207967 56175
rect 208001 56147 208029 56175
rect 207939 56085 207967 56113
rect 208001 56085 208029 56113
rect 207939 56023 207967 56051
rect 208001 56023 208029 56051
rect 207939 55961 207967 55989
rect 208001 55961 208029 55989
rect 217797 56147 217825 56175
rect 217859 56147 217887 56175
rect 217921 56147 217949 56175
rect 217983 56147 218011 56175
rect 217797 56085 217825 56113
rect 217859 56085 217887 56113
rect 217921 56085 217949 56113
rect 217983 56085 218011 56113
rect 217797 56023 217825 56051
rect 217859 56023 217887 56051
rect 217921 56023 217949 56051
rect 217983 56023 218011 56051
rect 217797 55961 217825 55989
rect 217859 55961 217887 55989
rect 217921 55961 217949 55989
rect 217983 55961 218011 55989
rect 204297 50147 204325 50175
rect 204359 50147 204387 50175
rect 204421 50147 204449 50175
rect 204483 50147 204511 50175
rect 204297 50085 204325 50113
rect 204359 50085 204387 50113
rect 204421 50085 204449 50113
rect 204483 50085 204511 50113
rect 204297 50023 204325 50051
rect 204359 50023 204387 50051
rect 204421 50023 204449 50051
rect 204483 50023 204511 50051
rect 204297 49961 204325 49989
rect 204359 49961 204387 49989
rect 204421 49961 204449 49989
rect 204483 49961 204511 49989
rect 215619 50147 215647 50175
rect 215681 50147 215709 50175
rect 215619 50085 215647 50113
rect 215681 50085 215709 50113
rect 215619 50023 215647 50051
rect 215681 50023 215709 50051
rect 215619 49961 215647 49989
rect 215681 49961 215709 49989
rect 207939 47147 207967 47175
rect 208001 47147 208029 47175
rect 207939 47085 207967 47113
rect 208001 47085 208029 47113
rect 207939 47023 207967 47051
rect 208001 47023 208029 47051
rect 207939 46961 207967 46989
rect 208001 46961 208029 46989
rect 217797 47147 217825 47175
rect 217859 47147 217887 47175
rect 217921 47147 217949 47175
rect 217983 47147 218011 47175
rect 217797 47085 217825 47113
rect 217859 47085 217887 47113
rect 217921 47085 217949 47113
rect 217983 47085 218011 47113
rect 217797 47023 217825 47051
rect 217859 47023 217887 47051
rect 217921 47023 217949 47051
rect 217983 47023 218011 47051
rect 217797 46961 217825 46989
rect 217859 46961 217887 46989
rect 217921 46961 217949 46989
rect 217983 46961 218011 46989
rect 204297 41147 204325 41175
rect 204359 41147 204387 41175
rect 204421 41147 204449 41175
rect 204483 41147 204511 41175
rect 204297 41085 204325 41113
rect 204359 41085 204387 41113
rect 204421 41085 204449 41113
rect 204483 41085 204511 41113
rect 204297 41023 204325 41051
rect 204359 41023 204387 41051
rect 204421 41023 204449 41051
rect 204483 41023 204511 41051
rect 204297 40961 204325 40989
rect 204359 40961 204387 40989
rect 204421 40961 204449 40989
rect 204483 40961 204511 40989
rect 215619 41147 215647 41175
rect 215681 41147 215709 41175
rect 215619 41085 215647 41113
rect 215681 41085 215709 41113
rect 215619 41023 215647 41051
rect 215681 41023 215709 41051
rect 215619 40961 215647 40989
rect 215681 40961 215709 40989
rect 207939 38147 207967 38175
rect 208001 38147 208029 38175
rect 207939 38085 207967 38113
rect 208001 38085 208029 38113
rect 207939 38023 207967 38051
rect 208001 38023 208029 38051
rect 207939 37961 207967 37989
rect 208001 37961 208029 37989
rect 217797 38147 217825 38175
rect 217859 38147 217887 38175
rect 217921 38147 217949 38175
rect 217983 38147 218011 38175
rect 217797 38085 217825 38113
rect 217859 38085 217887 38113
rect 217921 38085 217949 38113
rect 217983 38085 218011 38113
rect 217797 38023 217825 38051
rect 217859 38023 217887 38051
rect 217921 38023 217949 38051
rect 217983 38023 218011 38051
rect 217797 37961 217825 37989
rect 217859 37961 217887 37989
rect 217921 37961 217949 37989
rect 217983 37961 218011 37989
rect 204297 32147 204325 32175
rect 204359 32147 204387 32175
rect 204421 32147 204449 32175
rect 204483 32147 204511 32175
rect 204297 32085 204325 32113
rect 204359 32085 204387 32113
rect 204421 32085 204449 32113
rect 204483 32085 204511 32113
rect 204297 32023 204325 32051
rect 204359 32023 204387 32051
rect 204421 32023 204449 32051
rect 204483 32023 204511 32051
rect 204297 31961 204325 31989
rect 204359 31961 204387 31989
rect 204421 31961 204449 31989
rect 204483 31961 204511 31989
rect 215619 32147 215647 32175
rect 215681 32147 215709 32175
rect 215619 32085 215647 32113
rect 215681 32085 215709 32113
rect 215619 32023 215647 32051
rect 215681 32023 215709 32051
rect 215619 31961 215647 31989
rect 215681 31961 215709 31989
rect 207939 29147 207967 29175
rect 208001 29147 208029 29175
rect 207939 29085 207967 29113
rect 208001 29085 208029 29113
rect 207939 29023 207967 29051
rect 208001 29023 208029 29051
rect 207939 28961 207967 28989
rect 208001 28961 208029 28989
rect 217797 29147 217825 29175
rect 217859 29147 217887 29175
rect 217921 29147 217949 29175
rect 217983 29147 218011 29175
rect 217797 29085 217825 29113
rect 217859 29085 217887 29113
rect 217921 29085 217949 29113
rect 217983 29085 218011 29113
rect 217797 29023 217825 29051
rect 217859 29023 217887 29051
rect 217921 29023 217949 29051
rect 217983 29023 218011 29051
rect 217797 28961 217825 28989
rect 217859 28961 217887 28989
rect 217921 28961 217949 28989
rect 217983 28961 218011 28989
rect 204297 23147 204325 23175
rect 204359 23147 204387 23175
rect 204421 23147 204449 23175
rect 204483 23147 204511 23175
rect 204297 23085 204325 23113
rect 204359 23085 204387 23113
rect 204421 23085 204449 23113
rect 204483 23085 204511 23113
rect 204297 23023 204325 23051
rect 204359 23023 204387 23051
rect 204421 23023 204449 23051
rect 204483 23023 204511 23051
rect 204297 22961 204325 22989
rect 204359 22961 204387 22989
rect 204421 22961 204449 22989
rect 204483 22961 204511 22989
rect 215619 23147 215647 23175
rect 215681 23147 215709 23175
rect 215619 23085 215647 23113
rect 215681 23085 215709 23113
rect 215619 23023 215647 23051
rect 215681 23023 215709 23051
rect 215619 22961 215647 22989
rect 215681 22961 215709 22989
rect 207939 20147 207967 20175
rect 208001 20147 208029 20175
rect 207939 20085 207967 20113
rect 208001 20085 208029 20113
rect 207939 20023 207967 20051
rect 208001 20023 208029 20051
rect 207939 19961 207967 19989
rect 208001 19961 208029 19989
rect 217797 20147 217825 20175
rect 217859 20147 217887 20175
rect 217921 20147 217949 20175
rect 217983 20147 218011 20175
rect 217797 20085 217825 20113
rect 217859 20085 217887 20113
rect 217921 20085 217949 20113
rect 217983 20085 218011 20113
rect 217797 20023 217825 20051
rect 217859 20023 217887 20051
rect 217921 20023 217949 20051
rect 217983 20023 218011 20051
rect 217797 19961 217825 19989
rect 217859 19961 217887 19989
rect 217921 19961 217949 19989
rect 217983 19961 218011 19989
rect 204297 14147 204325 14175
rect 204359 14147 204387 14175
rect 204421 14147 204449 14175
rect 204483 14147 204511 14175
rect 204297 14085 204325 14113
rect 204359 14085 204387 14113
rect 204421 14085 204449 14113
rect 204483 14085 204511 14113
rect 204297 14023 204325 14051
rect 204359 14023 204387 14051
rect 204421 14023 204449 14051
rect 204483 14023 204511 14051
rect 204297 13961 204325 13989
rect 204359 13961 204387 13989
rect 204421 13961 204449 13989
rect 204483 13961 204511 13989
rect 215619 14147 215647 14175
rect 215681 14147 215709 14175
rect 215619 14085 215647 14113
rect 215681 14085 215709 14113
rect 215619 14023 215647 14051
rect 215681 14023 215709 14051
rect 215619 13961 215647 13989
rect 215681 13961 215709 13989
rect 207939 11147 207967 11175
rect 208001 11147 208029 11175
rect 207939 11085 207967 11113
rect 208001 11085 208029 11113
rect 207939 11023 207967 11051
rect 208001 11023 208029 11051
rect 207939 10961 207967 10989
rect 208001 10961 208029 10989
rect 217797 11147 217825 11175
rect 217859 11147 217887 11175
rect 217921 11147 217949 11175
rect 217983 11147 218011 11175
rect 217797 11085 217825 11113
rect 217859 11085 217887 11113
rect 217921 11085 217949 11113
rect 217983 11085 218011 11113
rect 217797 11023 217825 11051
rect 217859 11023 217887 11051
rect 217921 11023 217949 11051
rect 217983 11023 218011 11051
rect 217797 10961 217825 10989
rect 217859 10961 217887 10989
rect 217921 10961 217949 10989
rect 217983 10961 218011 10989
rect 204297 5147 204325 5175
rect 204359 5147 204387 5175
rect 204421 5147 204449 5175
rect 204483 5147 204511 5175
rect 204297 5085 204325 5113
rect 204359 5085 204387 5113
rect 204421 5085 204449 5113
rect 204483 5085 204511 5113
rect 204297 5023 204325 5051
rect 204359 5023 204387 5051
rect 204421 5023 204449 5051
rect 204483 5023 204511 5051
rect 204297 4961 204325 4989
rect 204359 4961 204387 4989
rect 204421 4961 204449 4989
rect 204483 4961 204511 4989
rect 215619 5147 215647 5175
rect 215681 5147 215709 5175
rect 215619 5085 215647 5113
rect 215681 5085 215709 5113
rect 215619 5023 215647 5051
rect 215681 5023 215709 5051
rect 215619 4961 215647 4989
rect 215681 4961 215709 4989
rect 204297 -588 204325 -560
rect 204359 -588 204387 -560
rect 204421 -588 204449 -560
rect 204483 -588 204511 -560
rect 204297 -650 204325 -622
rect 204359 -650 204387 -622
rect 204421 -650 204449 -622
rect 204483 -650 204511 -622
rect 204297 -712 204325 -684
rect 204359 -712 204387 -684
rect 204421 -712 204449 -684
rect 204483 -712 204511 -684
rect 204297 -774 204325 -746
rect 204359 -774 204387 -746
rect 204421 -774 204449 -746
rect 204483 -774 204511 -746
rect 217797 2147 217825 2175
rect 217859 2147 217887 2175
rect 217921 2147 217949 2175
rect 217983 2147 218011 2175
rect 217797 2085 217825 2113
rect 217859 2085 217887 2113
rect 217921 2085 217949 2113
rect 217983 2085 218011 2113
rect 217797 2023 217825 2051
rect 217859 2023 217887 2051
rect 217921 2023 217949 2051
rect 217983 2023 218011 2051
rect 217797 1961 217825 1989
rect 217859 1961 217887 1989
rect 217921 1961 217949 1989
rect 217983 1961 218011 1989
rect 217797 -108 217825 -80
rect 217859 -108 217887 -80
rect 217921 -108 217949 -80
rect 217983 -108 218011 -80
rect 217797 -170 217825 -142
rect 217859 -170 217887 -142
rect 217921 -170 217949 -142
rect 217983 -170 218011 -142
rect 217797 -232 217825 -204
rect 217859 -232 217887 -204
rect 217921 -232 217949 -204
rect 217983 -232 218011 -204
rect 217797 -294 217825 -266
rect 217859 -294 217887 -266
rect 217921 -294 217949 -266
rect 217983 -294 218011 -266
rect 219657 299058 219685 299086
rect 219719 299058 219747 299086
rect 219781 299058 219809 299086
rect 219843 299058 219871 299086
rect 219657 298996 219685 299024
rect 219719 298996 219747 299024
rect 219781 298996 219809 299024
rect 219843 298996 219871 299024
rect 219657 298934 219685 298962
rect 219719 298934 219747 298962
rect 219781 298934 219809 298962
rect 219843 298934 219871 298962
rect 219657 298872 219685 298900
rect 219719 298872 219747 298900
rect 219781 298872 219809 298900
rect 219843 298872 219871 298900
rect 219657 293147 219685 293175
rect 219719 293147 219747 293175
rect 219781 293147 219809 293175
rect 219843 293147 219871 293175
rect 219657 293085 219685 293113
rect 219719 293085 219747 293113
rect 219781 293085 219809 293113
rect 219843 293085 219871 293113
rect 219657 293023 219685 293051
rect 219719 293023 219747 293051
rect 219781 293023 219809 293051
rect 219843 293023 219871 293051
rect 219657 292961 219685 292989
rect 219719 292961 219747 292989
rect 219781 292961 219809 292989
rect 219843 292961 219871 292989
rect 219657 284147 219685 284175
rect 219719 284147 219747 284175
rect 219781 284147 219809 284175
rect 219843 284147 219871 284175
rect 219657 284085 219685 284113
rect 219719 284085 219747 284113
rect 219781 284085 219809 284113
rect 219843 284085 219871 284113
rect 219657 284023 219685 284051
rect 219719 284023 219747 284051
rect 219781 284023 219809 284051
rect 219843 284023 219871 284051
rect 219657 283961 219685 283989
rect 219719 283961 219747 283989
rect 219781 283961 219809 283989
rect 219843 283961 219871 283989
rect 219657 275147 219685 275175
rect 219719 275147 219747 275175
rect 219781 275147 219809 275175
rect 219843 275147 219871 275175
rect 219657 275085 219685 275113
rect 219719 275085 219747 275113
rect 219781 275085 219809 275113
rect 219843 275085 219871 275113
rect 219657 275023 219685 275051
rect 219719 275023 219747 275051
rect 219781 275023 219809 275051
rect 219843 275023 219871 275051
rect 219657 274961 219685 274989
rect 219719 274961 219747 274989
rect 219781 274961 219809 274989
rect 219843 274961 219871 274989
rect 219657 266147 219685 266175
rect 219719 266147 219747 266175
rect 219781 266147 219809 266175
rect 219843 266147 219871 266175
rect 219657 266085 219685 266113
rect 219719 266085 219747 266113
rect 219781 266085 219809 266113
rect 219843 266085 219871 266113
rect 219657 266023 219685 266051
rect 219719 266023 219747 266051
rect 219781 266023 219809 266051
rect 219843 266023 219871 266051
rect 219657 265961 219685 265989
rect 219719 265961 219747 265989
rect 219781 265961 219809 265989
rect 219843 265961 219871 265989
rect 219657 257147 219685 257175
rect 219719 257147 219747 257175
rect 219781 257147 219809 257175
rect 219843 257147 219871 257175
rect 219657 257085 219685 257113
rect 219719 257085 219747 257113
rect 219781 257085 219809 257113
rect 219843 257085 219871 257113
rect 219657 257023 219685 257051
rect 219719 257023 219747 257051
rect 219781 257023 219809 257051
rect 219843 257023 219871 257051
rect 219657 256961 219685 256989
rect 219719 256961 219747 256989
rect 219781 256961 219809 256989
rect 219843 256961 219871 256989
rect 219657 248147 219685 248175
rect 219719 248147 219747 248175
rect 219781 248147 219809 248175
rect 219843 248147 219871 248175
rect 219657 248085 219685 248113
rect 219719 248085 219747 248113
rect 219781 248085 219809 248113
rect 219843 248085 219871 248113
rect 219657 248023 219685 248051
rect 219719 248023 219747 248051
rect 219781 248023 219809 248051
rect 219843 248023 219871 248051
rect 219657 247961 219685 247989
rect 219719 247961 219747 247989
rect 219781 247961 219809 247989
rect 219843 247961 219871 247989
rect 219657 239147 219685 239175
rect 219719 239147 219747 239175
rect 219781 239147 219809 239175
rect 219843 239147 219871 239175
rect 219657 239085 219685 239113
rect 219719 239085 219747 239113
rect 219781 239085 219809 239113
rect 219843 239085 219871 239113
rect 219657 239023 219685 239051
rect 219719 239023 219747 239051
rect 219781 239023 219809 239051
rect 219843 239023 219871 239051
rect 219657 238961 219685 238989
rect 219719 238961 219747 238989
rect 219781 238961 219809 238989
rect 219843 238961 219871 238989
rect 219657 230147 219685 230175
rect 219719 230147 219747 230175
rect 219781 230147 219809 230175
rect 219843 230147 219871 230175
rect 219657 230085 219685 230113
rect 219719 230085 219747 230113
rect 219781 230085 219809 230113
rect 219843 230085 219871 230113
rect 219657 230023 219685 230051
rect 219719 230023 219747 230051
rect 219781 230023 219809 230051
rect 219843 230023 219871 230051
rect 219657 229961 219685 229989
rect 219719 229961 219747 229989
rect 219781 229961 219809 229989
rect 219843 229961 219871 229989
rect 219657 221147 219685 221175
rect 219719 221147 219747 221175
rect 219781 221147 219809 221175
rect 219843 221147 219871 221175
rect 219657 221085 219685 221113
rect 219719 221085 219747 221113
rect 219781 221085 219809 221113
rect 219843 221085 219871 221113
rect 219657 221023 219685 221051
rect 219719 221023 219747 221051
rect 219781 221023 219809 221051
rect 219843 221023 219871 221051
rect 219657 220961 219685 220989
rect 219719 220961 219747 220989
rect 219781 220961 219809 220989
rect 219843 220961 219871 220989
rect 219657 212147 219685 212175
rect 219719 212147 219747 212175
rect 219781 212147 219809 212175
rect 219843 212147 219871 212175
rect 219657 212085 219685 212113
rect 219719 212085 219747 212113
rect 219781 212085 219809 212113
rect 219843 212085 219871 212113
rect 219657 212023 219685 212051
rect 219719 212023 219747 212051
rect 219781 212023 219809 212051
rect 219843 212023 219871 212051
rect 219657 211961 219685 211989
rect 219719 211961 219747 211989
rect 219781 211961 219809 211989
rect 219843 211961 219871 211989
rect 219657 203147 219685 203175
rect 219719 203147 219747 203175
rect 219781 203147 219809 203175
rect 219843 203147 219871 203175
rect 219657 203085 219685 203113
rect 219719 203085 219747 203113
rect 219781 203085 219809 203113
rect 219843 203085 219871 203113
rect 219657 203023 219685 203051
rect 219719 203023 219747 203051
rect 219781 203023 219809 203051
rect 219843 203023 219871 203051
rect 219657 202961 219685 202989
rect 219719 202961 219747 202989
rect 219781 202961 219809 202989
rect 219843 202961 219871 202989
rect 219657 194147 219685 194175
rect 219719 194147 219747 194175
rect 219781 194147 219809 194175
rect 219843 194147 219871 194175
rect 219657 194085 219685 194113
rect 219719 194085 219747 194113
rect 219781 194085 219809 194113
rect 219843 194085 219871 194113
rect 219657 194023 219685 194051
rect 219719 194023 219747 194051
rect 219781 194023 219809 194051
rect 219843 194023 219871 194051
rect 219657 193961 219685 193989
rect 219719 193961 219747 193989
rect 219781 193961 219809 193989
rect 219843 193961 219871 193989
rect 219657 185147 219685 185175
rect 219719 185147 219747 185175
rect 219781 185147 219809 185175
rect 219843 185147 219871 185175
rect 219657 185085 219685 185113
rect 219719 185085 219747 185113
rect 219781 185085 219809 185113
rect 219843 185085 219871 185113
rect 219657 185023 219685 185051
rect 219719 185023 219747 185051
rect 219781 185023 219809 185051
rect 219843 185023 219871 185051
rect 219657 184961 219685 184989
rect 219719 184961 219747 184989
rect 219781 184961 219809 184989
rect 219843 184961 219871 184989
rect 219657 176147 219685 176175
rect 219719 176147 219747 176175
rect 219781 176147 219809 176175
rect 219843 176147 219871 176175
rect 219657 176085 219685 176113
rect 219719 176085 219747 176113
rect 219781 176085 219809 176113
rect 219843 176085 219871 176113
rect 219657 176023 219685 176051
rect 219719 176023 219747 176051
rect 219781 176023 219809 176051
rect 219843 176023 219871 176051
rect 219657 175961 219685 175989
rect 219719 175961 219747 175989
rect 219781 175961 219809 175989
rect 219843 175961 219871 175989
rect 233157 298578 233185 298606
rect 233219 298578 233247 298606
rect 233281 298578 233309 298606
rect 233343 298578 233371 298606
rect 233157 298516 233185 298544
rect 233219 298516 233247 298544
rect 233281 298516 233309 298544
rect 233343 298516 233371 298544
rect 233157 298454 233185 298482
rect 233219 298454 233247 298482
rect 233281 298454 233309 298482
rect 233343 298454 233371 298482
rect 233157 298392 233185 298420
rect 233219 298392 233247 298420
rect 233281 298392 233309 298420
rect 233343 298392 233371 298420
rect 233157 290147 233185 290175
rect 233219 290147 233247 290175
rect 233281 290147 233309 290175
rect 233343 290147 233371 290175
rect 233157 290085 233185 290113
rect 233219 290085 233247 290113
rect 233281 290085 233309 290113
rect 233343 290085 233371 290113
rect 233157 290023 233185 290051
rect 233219 290023 233247 290051
rect 233281 290023 233309 290051
rect 233343 290023 233371 290051
rect 233157 289961 233185 289989
rect 233219 289961 233247 289989
rect 233281 289961 233309 289989
rect 233343 289961 233371 289989
rect 233157 281147 233185 281175
rect 233219 281147 233247 281175
rect 233281 281147 233309 281175
rect 233343 281147 233371 281175
rect 233157 281085 233185 281113
rect 233219 281085 233247 281113
rect 233281 281085 233309 281113
rect 233343 281085 233371 281113
rect 233157 281023 233185 281051
rect 233219 281023 233247 281051
rect 233281 281023 233309 281051
rect 233343 281023 233371 281051
rect 233157 280961 233185 280989
rect 233219 280961 233247 280989
rect 233281 280961 233309 280989
rect 233343 280961 233371 280989
rect 233157 272147 233185 272175
rect 233219 272147 233247 272175
rect 233281 272147 233309 272175
rect 233343 272147 233371 272175
rect 233157 272085 233185 272113
rect 233219 272085 233247 272113
rect 233281 272085 233309 272113
rect 233343 272085 233371 272113
rect 233157 272023 233185 272051
rect 233219 272023 233247 272051
rect 233281 272023 233309 272051
rect 233343 272023 233371 272051
rect 233157 271961 233185 271989
rect 233219 271961 233247 271989
rect 233281 271961 233309 271989
rect 233343 271961 233371 271989
rect 233157 263147 233185 263175
rect 233219 263147 233247 263175
rect 233281 263147 233309 263175
rect 233343 263147 233371 263175
rect 233157 263085 233185 263113
rect 233219 263085 233247 263113
rect 233281 263085 233309 263113
rect 233343 263085 233371 263113
rect 233157 263023 233185 263051
rect 233219 263023 233247 263051
rect 233281 263023 233309 263051
rect 233343 263023 233371 263051
rect 233157 262961 233185 262989
rect 233219 262961 233247 262989
rect 233281 262961 233309 262989
rect 233343 262961 233371 262989
rect 233157 254147 233185 254175
rect 233219 254147 233247 254175
rect 233281 254147 233309 254175
rect 233343 254147 233371 254175
rect 233157 254085 233185 254113
rect 233219 254085 233247 254113
rect 233281 254085 233309 254113
rect 233343 254085 233371 254113
rect 233157 254023 233185 254051
rect 233219 254023 233247 254051
rect 233281 254023 233309 254051
rect 233343 254023 233371 254051
rect 233157 253961 233185 253989
rect 233219 253961 233247 253989
rect 233281 253961 233309 253989
rect 233343 253961 233371 253989
rect 233157 245147 233185 245175
rect 233219 245147 233247 245175
rect 233281 245147 233309 245175
rect 233343 245147 233371 245175
rect 233157 245085 233185 245113
rect 233219 245085 233247 245113
rect 233281 245085 233309 245113
rect 233343 245085 233371 245113
rect 233157 245023 233185 245051
rect 233219 245023 233247 245051
rect 233281 245023 233309 245051
rect 233343 245023 233371 245051
rect 233157 244961 233185 244989
rect 233219 244961 233247 244989
rect 233281 244961 233309 244989
rect 233343 244961 233371 244989
rect 233157 236147 233185 236175
rect 233219 236147 233247 236175
rect 233281 236147 233309 236175
rect 233343 236147 233371 236175
rect 233157 236085 233185 236113
rect 233219 236085 233247 236113
rect 233281 236085 233309 236113
rect 233343 236085 233371 236113
rect 233157 236023 233185 236051
rect 233219 236023 233247 236051
rect 233281 236023 233309 236051
rect 233343 236023 233371 236051
rect 233157 235961 233185 235989
rect 233219 235961 233247 235989
rect 233281 235961 233309 235989
rect 233343 235961 233371 235989
rect 233157 227147 233185 227175
rect 233219 227147 233247 227175
rect 233281 227147 233309 227175
rect 233343 227147 233371 227175
rect 233157 227085 233185 227113
rect 233219 227085 233247 227113
rect 233281 227085 233309 227113
rect 233343 227085 233371 227113
rect 233157 227023 233185 227051
rect 233219 227023 233247 227051
rect 233281 227023 233309 227051
rect 233343 227023 233371 227051
rect 233157 226961 233185 226989
rect 233219 226961 233247 226989
rect 233281 226961 233309 226989
rect 233343 226961 233371 226989
rect 233157 218147 233185 218175
rect 233219 218147 233247 218175
rect 233281 218147 233309 218175
rect 233343 218147 233371 218175
rect 233157 218085 233185 218113
rect 233219 218085 233247 218113
rect 233281 218085 233309 218113
rect 233343 218085 233371 218113
rect 233157 218023 233185 218051
rect 233219 218023 233247 218051
rect 233281 218023 233309 218051
rect 233343 218023 233371 218051
rect 233157 217961 233185 217989
rect 233219 217961 233247 217989
rect 233281 217961 233309 217989
rect 233343 217961 233371 217989
rect 233157 209147 233185 209175
rect 233219 209147 233247 209175
rect 233281 209147 233309 209175
rect 233343 209147 233371 209175
rect 233157 209085 233185 209113
rect 233219 209085 233247 209113
rect 233281 209085 233309 209113
rect 233343 209085 233371 209113
rect 233157 209023 233185 209051
rect 233219 209023 233247 209051
rect 233281 209023 233309 209051
rect 233343 209023 233371 209051
rect 233157 208961 233185 208989
rect 233219 208961 233247 208989
rect 233281 208961 233309 208989
rect 233343 208961 233371 208989
rect 233157 200147 233185 200175
rect 233219 200147 233247 200175
rect 233281 200147 233309 200175
rect 233343 200147 233371 200175
rect 233157 200085 233185 200113
rect 233219 200085 233247 200113
rect 233281 200085 233309 200113
rect 233343 200085 233371 200113
rect 233157 200023 233185 200051
rect 233219 200023 233247 200051
rect 233281 200023 233309 200051
rect 233343 200023 233371 200051
rect 233157 199961 233185 199989
rect 233219 199961 233247 199989
rect 233281 199961 233309 199989
rect 233343 199961 233371 199989
rect 233157 191147 233185 191175
rect 233219 191147 233247 191175
rect 233281 191147 233309 191175
rect 233343 191147 233371 191175
rect 233157 191085 233185 191113
rect 233219 191085 233247 191113
rect 233281 191085 233309 191113
rect 233343 191085 233371 191113
rect 233157 191023 233185 191051
rect 233219 191023 233247 191051
rect 233281 191023 233309 191051
rect 233343 191023 233371 191051
rect 233157 190961 233185 190989
rect 233219 190961 233247 190989
rect 233281 190961 233309 190989
rect 233343 190961 233371 190989
rect 233157 182147 233185 182175
rect 233219 182147 233247 182175
rect 233281 182147 233309 182175
rect 233343 182147 233371 182175
rect 233157 182085 233185 182113
rect 233219 182085 233247 182113
rect 233281 182085 233309 182113
rect 233343 182085 233371 182113
rect 233157 182023 233185 182051
rect 233219 182023 233247 182051
rect 233281 182023 233309 182051
rect 233343 182023 233371 182051
rect 233157 181961 233185 181989
rect 233219 181961 233247 181989
rect 233281 181961 233309 181989
rect 233343 181961 233371 181989
rect 223299 173147 223327 173175
rect 223361 173147 223389 173175
rect 223299 173085 223327 173113
rect 223361 173085 223389 173113
rect 223299 173023 223327 173051
rect 223361 173023 223389 173051
rect 223299 172961 223327 172989
rect 223361 172961 223389 172989
rect 233157 173147 233185 173175
rect 233219 173147 233247 173175
rect 233281 173147 233309 173175
rect 233343 173147 233371 173175
rect 233157 173085 233185 173113
rect 233219 173085 233247 173113
rect 233281 173085 233309 173113
rect 233343 173085 233371 173113
rect 233157 173023 233185 173051
rect 233219 173023 233247 173051
rect 233281 173023 233309 173051
rect 233343 173023 233371 173051
rect 233157 172961 233185 172989
rect 233219 172961 233247 172989
rect 233281 172961 233309 172989
rect 233343 172961 233371 172989
rect 219657 167147 219685 167175
rect 219719 167147 219747 167175
rect 219781 167147 219809 167175
rect 219843 167147 219871 167175
rect 219657 167085 219685 167113
rect 219719 167085 219747 167113
rect 219781 167085 219809 167113
rect 219843 167085 219871 167113
rect 219657 167023 219685 167051
rect 219719 167023 219747 167051
rect 219781 167023 219809 167051
rect 219843 167023 219871 167051
rect 219657 166961 219685 166989
rect 219719 166961 219747 166989
rect 219781 166961 219809 166989
rect 219843 166961 219871 166989
rect 230979 167147 231007 167175
rect 231041 167147 231069 167175
rect 230979 167085 231007 167113
rect 231041 167085 231069 167113
rect 230979 167023 231007 167051
rect 231041 167023 231069 167051
rect 230979 166961 231007 166989
rect 231041 166961 231069 166989
rect 223299 164147 223327 164175
rect 223361 164147 223389 164175
rect 223299 164085 223327 164113
rect 223361 164085 223389 164113
rect 223299 164023 223327 164051
rect 223361 164023 223389 164051
rect 223299 163961 223327 163989
rect 223361 163961 223389 163989
rect 233157 164147 233185 164175
rect 233219 164147 233247 164175
rect 233281 164147 233309 164175
rect 233343 164147 233371 164175
rect 233157 164085 233185 164113
rect 233219 164085 233247 164113
rect 233281 164085 233309 164113
rect 233343 164085 233371 164113
rect 233157 164023 233185 164051
rect 233219 164023 233247 164051
rect 233281 164023 233309 164051
rect 233343 164023 233371 164051
rect 233157 163961 233185 163989
rect 233219 163961 233247 163989
rect 233281 163961 233309 163989
rect 233343 163961 233371 163989
rect 219657 158147 219685 158175
rect 219719 158147 219747 158175
rect 219781 158147 219809 158175
rect 219843 158147 219871 158175
rect 219657 158085 219685 158113
rect 219719 158085 219747 158113
rect 219781 158085 219809 158113
rect 219843 158085 219871 158113
rect 219657 158023 219685 158051
rect 219719 158023 219747 158051
rect 219781 158023 219809 158051
rect 219843 158023 219871 158051
rect 219657 157961 219685 157989
rect 219719 157961 219747 157989
rect 219781 157961 219809 157989
rect 219843 157961 219871 157989
rect 230979 158147 231007 158175
rect 231041 158147 231069 158175
rect 230979 158085 231007 158113
rect 231041 158085 231069 158113
rect 230979 158023 231007 158051
rect 231041 158023 231069 158051
rect 230979 157961 231007 157989
rect 231041 157961 231069 157989
rect 223299 155147 223327 155175
rect 223361 155147 223389 155175
rect 223299 155085 223327 155113
rect 223361 155085 223389 155113
rect 223299 155023 223327 155051
rect 223361 155023 223389 155051
rect 223299 154961 223327 154989
rect 223361 154961 223389 154989
rect 233157 155147 233185 155175
rect 233219 155147 233247 155175
rect 233281 155147 233309 155175
rect 233343 155147 233371 155175
rect 233157 155085 233185 155113
rect 233219 155085 233247 155113
rect 233281 155085 233309 155113
rect 233343 155085 233371 155113
rect 233157 155023 233185 155051
rect 233219 155023 233247 155051
rect 233281 155023 233309 155051
rect 233343 155023 233371 155051
rect 233157 154961 233185 154989
rect 233219 154961 233247 154989
rect 233281 154961 233309 154989
rect 233343 154961 233371 154989
rect 219657 149147 219685 149175
rect 219719 149147 219747 149175
rect 219781 149147 219809 149175
rect 219843 149147 219871 149175
rect 219657 149085 219685 149113
rect 219719 149085 219747 149113
rect 219781 149085 219809 149113
rect 219843 149085 219871 149113
rect 219657 149023 219685 149051
rect 219719 149023 219747 149051
rect 219781 149023 219809 149051
rect 219843 149023 219871 149051
rect 219657 148961 219685 148989
rect 219719 148961 219747 148989
rect 219781 148961 219809 148989
rect 219843 148961 219871 148989
rect 230979 149147 231007 149175
rect 231041 149147 231069 149175
rect 230979 149085 231007 149113
rect 231041 149085 231069 149113
rect 230979 149023 231007 149051
rect 231041 149023 231069 149051
rect 230979 148961 231007 148989
rect 231041 148961 231069 148989
rect 223299 146147 223327 146175
rect 223361 146147 223389 146175
rect 223299 146085 223327 146113
rect 223361 146085 223389 146113
rect 223299 146023 223327 146051
rect 223361 146023 223389 146051
rect 223299 145961 223327 145989
rect 223361 145961 223389 145989
rect 233157 146147 233185 146175
rect 233219 146147 233247 146175
rect 233281 146147 233309 146175
rect 233343 146147 233371 146175
rect 233157 146085 233185 146113
rect 233219 146085 233247 146113
rect 233281 146085 233309 146113
rect 233343 146085 233371 146113
rect 233157 146023 233185 146051
rect 233219 146023 233247 146051
rect 233281 146023 233309 146051
rect 233343 146023 233371 146051
rect 233157 145961 233185 145989
rect 233219 145961 233247 145989
rect 233281 145961 233309 145989
rect 233343 145961 233371 145989
rect 219657 140147 219685 140175
rect 219719 140147 219747 140175
rect 219781 140147 219809 140175
rect 219843 140147 219871 140175
rect 219657 140085 219685 140113
rect 219719 140085 219747 140113
rect 219781 140085 219809 140113
rect 219843 140085 219871 140113
rect 219657 140023 219685 140051
rect 219719 140023 219747 140051
rect 219781 140023 219809 140051
rect 219843 140023 219871 140051
rect 219657 139961 219685 139989
rect 219719 139961 219747 139989
rect 219781 139961 219809 139989
rect 219843 139961 219871 139989
rect 230979 140147 231007 140175
rect 231041 140147 231069 140175
rect 230979 140085 231007 140113
rect 231041 140085 231069 140113
rect 230979 140023 231007 140051
rect 231041 140023 231069 140051
rect 230979 139961 231007 139989
rect 231041 139961 231069 139989
rect 223299 137147 223327 137175
rect 223361 137147 223389 137175
rect 223299 137085 223327 137113
rect 223361 137085 223389 137113
rect 223299 137023 223327 137051
rect 223361 137023 223389 137051
rect 223299 136961 223327 136989
rect 223361 136961 223389 136989
rect 233157 137147 233185 137175
rect 233219 137147 233247 137175
rect 233281 137147 233309 137175
rect 233343 137147 233371 137175
rect 233157 137085 233185 137113
rect 233219 137085 233247 137113
rect 233281 137085 233309 137113
rect 233343 137085 233371 137113
rect 233157 137023 233185 137051
rect 233219 137023 233247 137051
rect 233281 137023 233309 137051
rect 233343 137023 233371 137051
rect 233157 136961 233185 136989
rect 233219 136961 233247 136989
rect 233281 136961 233309 136989
rect 233343 136961 233371 136989
rect 219657 131147 219685 131175
rect 219719 131147 219747 131175
rect 219781 131147 219809 131175
rect 219843 131147 219871 131175
rect 219657 131085 219685 131113
rect 219719 131085 219747 131113
rect 219781 131085 219809 131113
rect 219843 131085 219871 131113
rect 219657 131023 219685 131051
rect 219719 131023 219747 131051
rect 219781 131023 219809 131051
rect 219843 131023 219871 131051
rect 219657 130961 219685 130989
rect 219719 130961 219747 130989
rect 219781 130961 219809 130989
rect 219843 130961 219871 130989
rect 230979 131147 231007 131175
rect 231041 131147 231069 131175
rect 230979 131085 231007 131113
rect 231041 131085 231069 131113
rect 230979 131023 231007 131051
rect 231041 131023 231069 131051
rect 230979 130961 231007 130989
rect 231041 130961 231069 130989
rect 223299 128147 223327 128175
rect 223361 128147 223389 128175
rect 223299 128085 223327 128113
rect 223361 128085 223389 128113
rect 223299 128023 223327 128051
rect 223361 128023 223389 128051
rect 223299 127961 223327 127989
rect 223361 127961 223389 127989
rect 233157 128147 233185 128175
rect 233219 128147 233247 128175
rect 233281 128147 233309 128175
rect 233343 128147 233371 128175
rect 233157 128085 233185 128113
rect 233219 128085 233247 128113
rect 233281 128085 233309 128113
rect 233343 128085 233371 128113
rect 233157 128023 233185 128051
rect 233219 128023 233247 128051
rect 233281 128023 233309 128051
rect 233343 128023 233371 128051
rect 233157 127961 233185 127989
rect 233219 127961 233247 127989
rect 233281 127961 233309 127989
rect 233343 127961 233371 127989
rect 219657 122147 219685 122175
rect 219719 122147 219747 122175
rect 219781 122147 219809 122175
rect 219843 122147 219871 122175
rect 219657 122085 219685 122113
rect 219719 122085 219747 122113
rect 219781 122085 219809 122113
rect 219843 122085 219871 122113
rect 219657 122023 219685 122051
rect 219719 122023 219747 122051
rect 219781 122023 219809 122051
rect 219843 122023 219871 122051
rect 219657 121961 219685 121989
rect 219719 121961 219747 121989
rect 219781 121961 219809 121989
rect 219843 121961 219871 121989
rect 230979 122147 231007 122175
rect 231041 122147 231069 122175
rect 230979 122085 231007 122113
rect 231041 122085 231069 122113
rect 230979 122023 231007 122051
rect 231041 122023 231069 122051
rect 230979 121961 231007 121989
rect 231041 121961 231069 121989
rect 223299 119147 223327 119175
rect 223361 119147 223389 119175
rect 223299 119085 223327 119113
rect 223361 119085 223389 119113
rect 223299 119023 223327 119051
rect 223361 119023 223389 119051
rect 223299 118961 223327 118989
rect 223361 118961 223389 118989
rect 233157 119147 233185 119175
rect 233219 119147 233247 119175
rect 233281 119147 233309 119175
rect 233343 119147 233371 119175
rect 233157 119085 233185 119113
rect 233219 119085 233247 119113
rect 233281 119085 233309 119113
rect 233343 119085 233371 119113
rect 233157 119023 233185 119051
rect 233219 119023 233247 119051
rect 233281 119023 233309 119051
rect 233343 119023 233371 119051
rect 233157 118961 233185 118989
rect 233219 118961 233247 118989
rect 233281 118961 233309 118989
rect 233343 118961 233371 118989
rect 219657 113147 219685 113175
rect 219719 113147 219747 113175
rect 219781 113147 219809 113175
rect 219843 113147 219871 113175
rect 219657 113085 219685 113113
rect 219719 113085 219747 113113
rect 219781 113085 219809 113113
rect 219843 113085 219871 113113
rect 219657 113023 219685 113051
rect 219719 113023 219747 113051
rect 219781 113023 219809 113051
rect 219843 113023 219871 113051
rect 219657 112961 219685 112989
rect 219719 112961 219747 112989
rect 219781 112961 219809 112989
rect 219843 112961 219871 112989
rect 230979 113147 231007 113175
rect 231041 113147 231069 113175
rect 230979 113085 231007 113113
rect 231041 113085 231069 113113
rect 230979 113023 231007 113051
rect 231041 113023 231069 113051
rect 230979 112961 231007 112989
rect 231041 112961 231069 112989
rect 223299 110147 223327 110175
rect 223361 110147 223389 110175
rect 223299 110085 223327 110113
rect 223361 110085 223389 110113
rect 223299 110023 223327 110051
rect 223361 110023 223389 110051
rect 223299 109961 223327 109989
rect 223361 109961 223389 109989
rect 233157 110147 233185 110175
rect 233219 110147 233247 110175
rect 233281 110147 233309 110175
rect 233343 110147 233371 110175
rect 233157 110085 233185 110113
rect 233219 110085 233247 110113
rect 233281 110085 233309 110113
rect 233343 110085 233371 110113
rect 233157 110023 233185 110051
rect 233219 110023 233247 110051
rect 233281 110023 233309 110051
rect 233343 110023 233371 110051
rect 233157 109961 233185 109989
rect 233219 109961 233247 109989
rect 233281 109961 233309 109989
rect 233343 109961 233371 109989
rect 219657 104147 219685 104175
rect 219719 104147 219747 104175
rect 219781 104147 219809 104175
rect 219843 104147 219871 104175
rect 219657 104085 219685 104113
rect 219719 104085 219747 104113
rect 219781 104085 219809 104113
rect 219843 104085 219871 104113
rect 219657 104023 219685 104051
rect 219719 104023 219747 104051
rect 219781 104023 219809 104051
rect 219843 104023 219871 104051
rect 219657 103961 219685 103989
rect 219719 103961 219747 103989
rect 219781 103961 219809 103989
rect 219843 103961 219871 103989
rect 230979 104147 231007 104175
rect 231041 104147 231069 104175
rect 230979 104085 231007 104113
rect 231041 104085 231069 104113
rect 230979 104023 231007 104051
rect 231041 104023 231069 104051
rect 230979 103961 231007 103989
rect 231041 103961 231069 103989
rect 223299 101147 223327 101175
rect 223361 101147 223389 101175
rect 223299 101085 223327 101113
rect 223361 101085 223389 101113
rect 223299 101023 223327 101051
rect 223361 101023 223389 101051
rect 223299 100961 223327 100989
rect 223361 100961 223389 100989
rect 233157 101147 233185 101175
rect 233219 101147 233247 101175
rect 233281 101147 233309 101175
rect 233343 101147 233371 101175
rect 233157 101085 233185 101113
rect 233219 101085 233247 101113
rect 233281 101085 233309 101113
rect 233343 101085 233371 101113
rect 233157 101023 233185 101051
rect 233219 101023 233247 101051
rect 233281 101023 233309 101051
rect 233343 101023 233371 101051
rect 233157 100961 233185 100989
rect 233219 100961 233247 100989
rect 233281 100961 233309 100989
rect 233343 100961 233371 100989
rect 219657 95147 219685 95175
rect 219719 95147 219747 95175
rect 219781 95147 219809 95175
rect 219843 95147 219871 95175
rect 219657 95085 219685 95113
rect 219719 95085 219747 95113
rect 219781 95085 219809 95113
rect 219843 95085 219871 95113
rect 219657 95023 219685 95051
rect 219719 95023 219747 95051
rect 219781 95023 219809 95051
rect 219843 95023 219871 95051
rect 219657 94961 219685 94989
rect 219719 94961 219747 94989
rect 219781 94961 219809 94989
rect 219843 94961 219871 94989
rect 230979 95147 231007 95175
rect 231041 95147 231069 95175
rect 230979 95085 231007 95113
rect 231041 95085 231069 95113
rect 230979 95023 231007 95051
rect 231041 95023 231069 95051
rect 230979 94961 231007 94989
rect 231041 94961 231069 94989
rect 223299 92147 223327 92175
rect 223361 92147 223389 92175
rect 223299 92085 223327 92113
rect 223361 92085 223389 92113
rect 223299 92023 223327 92051
rect 223361 92023 223389 92051
rect 223299 91961 223327 91989
rect 223361 91961 223389 91989
rect 233157 92147 233185 92175
rect 233219 92147 233247 92175
rect 233281 92147 233309 92175
rect 233343 92147 233371 92175
rect 233157 92085 233185 92113
rect 233219 92085 233247 92113
rect 233281 92085 233309 92113
rect 233343 92085 233371 92113
rect 233157 92023 233185 92051
rect 233219 92023 233247 92051
rect 233281 92023 233309 92051
rect 233343 92023 233371 92051
rect 233157 91961 233185 91989
rect 233219 91961 233247 91989
rect 233281 91961 233309 91989
rect 233343 91961 233371 91989
rect 219657 86147 219685 86175
rect 219719 86147 219747 86175
rect 219781 86147 219809 86175
rect 219843 86147 219871 86175
rect 219657 86085 219685 86113
rect 219719 86085 219747 86113
rect 219781 86085 219809 86113
rect 219843 86085 219871 86113
rect 219657 86023 219685 86051
rect 219719 86023 219747 86051
rect 219781 86023 219809 86051
rect 219843 86023 219871 86051
rect 219657 85961 219685 85989
rect 219719 85961 219747 85989
rect 219781 85961 219809 85989
rect 219843 85961 219871 85989
rect 230979 86147 231007 86175
rect 231041 86147 231069 86175
rect 230979 86085 231007 86113
rect 231041 86085 231069 86113
rect 230979 86023 231007 86051
rect 231041 86023 231069 86051
rect 230979 85961 231007 85989
rect 231041 85961 231069 85989
rect 223299 83147 223327 83175
rect 223361 83147 223389 83175
rect 223299 83085 223327 83113
rect 223361 83085 223389 83113
rect 223299 83023 223327 83051
rect 223361 83023 223389 83051
rect 223299 82961 223327 82989
rect 223361 82961 223389 82989
rect 233157 83147 233185 83175
rect 233219 83147 233247 83175
rect 233281 83147 233309 83175
rect 233343 83147 233371 83175
rect 233157 83085 233185 83113
rect 233219 83085 233247 83113
rect 233281 83085 233309 83113
rect 233343 83085 233371 83113
rect 233157 83023 233185 83051
rect 233219 83023 233247 83051
rect 233281 83023 233309 83051
rect 233343 83023 233371 83051
rect 233157 82961 233185 82989
rect 233219 82961 233247 82989
rect 233281 82961 233309 82989
rect 233343 82961 233371 82989
rect 219657 77147 219685 77175
rect 219719 77147 219747 77175
rect 219781 77147 219809 77175
rect 219843 77147 219871 77175
rect 219657 77085 219685 77113
rect 219719 77085 219747 77113
rect 219781 77085 219809 77113
rect 219843 77085 219871 77113
rect 219657 77023 219685 77051
rect 219719 77023 219747 77051
rect 219781 77023 219809 77051
rect 219843 77023 219871 77051
rect 219657 76961 219685 76989
rect 219719 76961 219747 76989
rect 219781 76961 219809 76989
rect 219843 76961 219871 76989
rect 230979 77147 231007 77175
rect 231041 77147 231069 77175
rect 230979 77085 231007 77113
rect 231041 77085 231069 77113
rect 230979 77023 231007 77051
rect 231041 77023 231069 77051
rect 230979 76961 231007 76989
rect 231041 76961 231069 76989
rect 223299 74147 223327 74175
rect 223361 74147 223389 74175
rect 223299 74085 223327 74113
rect 223361 74085 223389 74113
rect 223299 74023 223327 74051
rect 223361 74023 223389 74051
rect 223299 73961 223327 73989
rect 223361 73961 223389 73989
rect 233157 74147 233185 74175
rect 233219 74147 233247 74175
rect 233281 74147 233309 74175
rect 233343 74147 233371 74175
rect 233157 74085 233185 74113
rect 233219 74085 233247 74113
rect 233281 74085 233309 74113
rect 233343 74085 233371 74113
rect 233157 74023 233185 74051
rect 233219 74023 233247 74051
rect 233281 74023 233309 74051
rect 233343 74023 233371 74051
rect 233157 73961 233185 73989
rect 233219 73961 233247 73989
rect 233281 73961 233309 73989
rect 233343 73961 233371 73989
rect 219657 68147 219685 68175
rect 219719 68147 219747 68175
rect 219781 68147 219809 68175
rect 219843 68147 219871 68175
rect 219657 68085 219685 68113
rect 219719 68085 219747 68113
rect 219781 68085 219809 68113
rect 219843 68085 219871 68113
rect 219657 68023 219685 68051
rect 219719 68023 219747 68051
rect 219781 68023 219809 68051
rect 219843 68023 219871 68051
rect 219657 67961 219685 67989
rect 219719 67961 219747 67989
rect 219781 67961 219809 67989
rect 219843 67961 219871 67989
rect 230979 68147 231007 68175
rect 231041 68147 231069 68175
rect 230979 68085 231007 68113
rect 231041 68085 231069 68113
rect 230979 68023 231007 68051
rect 231041 68023 231069 68051
rect 230979 67961 231007 67989
rect 231041 67961 231069 67989
rect 223299 65147 223327 65175
rect 223361 65147 223389 65175
rect 223299 65085 223327 65113
rect 223361 65085 223389 65113
rect 223299 65023 223327 65051
rect 223361 65023 223389 65051
rect 223299 64961 223327 64989
rect 223361 64961 223389 64989
rect 233157 65147 233185 65175
rect 233219 65147 233247 65175
rect 233281 65147 233309 65175
rect 233343 65147 233371 65175
rect 233157 65085 233185 65113
rect 233219 65085 233247 65113
rect 233281 65085 233309 65113
rect 233343 65085 233371 65113
rect 233157 65023 233185 65051
rect 233219 65023 233247 65051
rect 233281 65023 233309 65051
rect 233343 65023 233371 65051
rect 233157 64961 233185 64989
rect 233219 64961 233247 64989
rect 233281 64961 233309 64989
rect 233343 64961 233371 64989
rect 219657 59147 219685 59175
rect 219719 59147 219747 59175
rect 219781 59147 219809 59175
rect 219843 59147 219871 59175
rect 219657 59085 219685 59113
rect 219719 59085 219747 59113
rect 219781 59085 219809 59113
rect 219843 59085 219871 59113
rect 219657 59023 219685 59051
rect 219719 59023 219747 59051
rect 219781 59023 219809 59051
rect 219843 59023 219871 59051
rect 219657 58961 219685 58989
rect 219719 58961 219747 58989
rect 219781 58961 219809 58989
rect 219843 58961 219871 58989
rect 230979 59147 231007 59175
rect 231041 59147 231069 59175
rect 230979 59085 231007 59113
rect 231041 59085 231069 59113
rect 230979 59023 231007 59051
rect 231041 59023 231069 59051
rect 230979 58961 231007 58989
rect 231041 58961 231069 58989
rect 223299 56147 223327 56175
rect 223361 56147 223389 56175
rect 223299 56085 223327 56113
rect 223361 56085 223389 56113
rect 223299 56023 223327 56051
rect 223361 56023 223389 56051
rect 223299 55961 223327 55989
rect 223361 55961 223389 55989
rect 233157 56147 233185 56175
rect 233219 56147 233247 56175
rect 233281 56147 233309 56175
rect 233343 56147 233371 56175
rect 233157 56085 233185 56113
rect 233219 56085 233247 56113
rect 233281 56085 233309 56113
rect 233343 56085 233371 56113
rect 233157 56023 233185 56051
rect 233219 56023 233247 56051
rect 233281 56023 233309 56051
rect 233343 56023 233371 56051
rect 233157 55961 233185 55989
rect 233219 55961 233247 55989
rect 233281 55961 233309 55989
rect 233343 55961 233371 55989
rect 219657 50147 219685 50175
rect 219719 50147 219747 50175
rect 219781 50147 219809 50175
rect 219843 50147 219871 50175
rect 219657 50085 219685 50113
rect 219719 50085 219747 50113
rect 219781 50085 219809 50113
rect 219843 50085 219871 50113
rect 219657 50023 219685 50051
rect 219719 50023 219747 50051
rect 219781 50023 219809 50051
rect 219843 50023 219871 50051
rect 219657 49961 219685 49989
rect 219719 49961 219747 49989
rect 219781 49961 219809 49989
rect 219843 49961 219871 49989
rect 230979 50147 231007 50175
rect 231041 50147 231069 50175
rect 230979 50085 231007 50113
rect 231041 50085 231069 50113
rect 230979 50023 231007 50051
rect 231041 50023 231069 50051
rect 230979 49961 231007 49989
rect 231041 49961 231069 49989
rect 223299 47147 223327 47175
rect 223361 47147 223389 47175
rect 223299 47085 223327 47113
rect 223361 47085 223389 47113
rect 223299 47023 223327 47051
rect 223361 47023 223389 47051
rect 223299 46961 223327 46989
rect 223361 46961 223389 46989
rect 233157 47147 233185 47175
rect 233219 47147 233247 47175
rect 233281 47147 233309 47175
rect 233343 47147 233371 47175
rect 233157 47085 233185 47113
rect 233219 47085 233247 47113
rect 233281 47085 233309 47113
rect 233343 47085 233371 47113
rect 233157 47023 233185 47051
rect 233219 47023 233247 47051
rect 233281 47023 233309 47051
rect 233343 47023 233371 47051
rect 233157 46961 233185 46989
rect 233219 46961 233247 46989
rect 233281 46961 233309 46989
rect 233343 46961 233371 46989
rect 219657 41147 219685 41175
rect 219719 41147 219747 41175
rect 219781 41147 219809 41175
rect 219843 41147 219871 41175
rect 219657 41085 219685 41113
rect 219719 41085 219747 41113
rect 219781 41085 219809 41113
rect 219843 41085 219871 41113
rect 219657 41023 219685 41051
rect 219719 41023 219747 41051
rect 219781 41023 219809 41051
rect 219843 41023 219871 41051
rect 219657 40961 219685 40989
rect 219719 40961 219747 40989
rect 219781 40961 219809 40989
rect 219843 40961 219871 40989
rect 230979 41147 231007 41175
rect 231041 41147 231069 41175
rect 230979 41085 231007 41113
rect 231041 41085 231069 41113
rect 230979 41023 231007 41051
rect 231041 41023 231069 41051
rect 230979 40961 231007 40989
rect 231041 40961 231069 40989
rect 223299 38147 223327 38175
rect 223361 38147 223389 38175
rect 223299 38085 223327 38113
rect 223361 38085 223389 38113
rect 223299 38023 223327 38051
rect 223361 38023 223389 38051
rect 223299 37961 223327 37989
rect 223361 37961 223389 37989
rect 233157 38147 233185 38175
rect 233219 38147 233247 38175
rect 233281 38147 233309 38175
rect 233343 38147 233371 38175
rect 233157 38085 233185 38113
rect 233219 38085 233247 38113
rect 233281 38085 233309 38113
rect 233343 38085 233371 38113
rect 233157 38023 233185 38051
rect 233219 38023 233247 38051
rect 233281 38023 233309 38051
rect 233343 38023 233371 38051
rect 233157 37961 233185 37989
rect 233219 37961 233247 37989
rect 233281 37961 233309 37989
rect 233343 37961 233371 37989
rect 219657 32147 219685 32175
rect 219719 32147 219747 32175
rect 219781 32147 219809 32175
rect 219843 32147 219871 32175
rect 219657 32085 219685 32113
rect 219719 32085 219747 32113
rect 219781 32085 219809 32113
rect 219843 32085 219871 32113
rect 219657 32023 219685 32051
rect 219719 32023 219747 32051
rect 219781 32023 219809 32051
rect 219843 32023 219871 32051
rect 219657 31961 219685 31989
rect 219719 31961 219747 31989
rect 219781 31961 219809 31989
rect 219843 31961 219871 31989
rect 230979 32147 231007 32175
rect 231041 32147 231069 32175
rect 230979 32085 231007 32113
rect 231041 32085 231069 32113
rect 230979 32023 231007 32051
rect 231041 32023 231069 32051
rect 230979 31961 231007 31989
rect 231041 31961 231069 31989
rect 223299 29147 223327 29175
rect 223361 29147 223389 29175
rect 223299 29085 223327 29113
rect 223361 29085 223389 29113
rect 223299 29023 223327 29051
rect 223361 29023 223389 29051
rect 223299 28961 223327 28989
rect 223361 28961 223389 28989
rect 233157 29147 233185 29175
rect 233219 29147 233247 29175
rect 233281 29147 233309 29175
rect 233343 29147 233371 29175
rect 233157 29085 233185 29113
rect 233219 29085 233247 29113
rect 233281 29085 233309 29113
rect 233343 29085 233371 29113
rect 233157 29023 233185 29051
rect 233219 29023 233247 29051
rect 233281 29023 233309 29051
rect 233343 29023 233371 29051
rect 233157 28961 233185 28989
rect 233219 28961 233247 28989
rect 233281 28961 233309 28989
rect 233343 28961 233371 28989
rect 219657 23147 219685 23175
rect 219719 23147 219747 23175
rect 219781 23147 219809 23175
rect 219843 23147 219871 23175
rect 219657 23085 219685 23113
rect 219719 23085 219747 23113
rect 219781 23085 219809 23113
rect 219843 23085 219871 23113
rect 219657 23023 219685 23051
rect 219719 23023 219747 23051
rect 219781 23023 219809 23051
rect 219843 23023 219871 23051
rect 219657 22961 219685 22989
rect 219719 22961 219747 22989
rect 219781 22961 219809 22989
rect 219843 22961 219871 22989
rect 230979 23147 231007 23175
rect 231041 23147 231069 23175
rect 230979 23085 231007 23113
rect 231041 23085 231069 23113
rect 230979 23023 231007 23051
rect 231041 23023 231069 23051
rect 230979 22961 231007 22989
rect 231041 22961 231069 22989
rect 223299 20147 223327 20175
rect 223361 20147 223389 20175
rect 223299 20085 223327 20113
rect 223361 20085 223389 20113
rect 223299 20023 223327 20051
rect 223361 20023 223389 20051
rect 223299 19961 223327 19989
rect 223361 19961 223389 19989
rect 233157 20147 233185 20175
rect 233219 20147 233247 20175
rect 233281 20147 233309 20175
rect 233343 20147 233371 20175
rect 233157 20085 233185 20113
rect 233219 20085 233247 20113
rect 233281 20085 233309 20113
rect 233343 20085 233371 20113
rect 233157 20023 233185 20051
rect 233219 20023 233247 20051
rect 233281 20023 233309 20051
rect 233343 20023 233371 20051
rect 233157 19961 233185 19989
rect 233219 19961 233247 19989
rect 233281 19961 233309 19989
rect 233343 19961 233371 19989
rect 219657 14147 219685 14175
rect 219719 14147 219747 14175
rect 219781 14147 219809 14175
rect 219843 14147 219871 14175
rect 219657 14085 219685 14113
rect 219719 14085 219747 14113
rect 219781 14085 219809 14113
rect 219843 14085 219871 14113
rect 219657 14023 219685 14051
rect 219719 14023 219747 14051
rect 219781 14023 219809 14051
rect 219843 14023 219871 14051
rect 219657 13961 219685 13989
rect 219719 13961 219747 13989
rect 219781 13961 219809 13989
rect 219843 13961 219871 13989
rect 230979 14147 231007 14175
rect 231041 14147 231069 14175
rect 230979 14085 231007 14113
rect 231041 14085 231069 14113
rect 230979 14023 231007 14051
rect 231041 14023 231069 14051
rect 230979 13961 231007 13989
rect 231041 13961 231069 13989
rect 223299 11147 223327 11175
rect 223361 11147 223389 11175
rect 223299 11085 223327 11113
rect 223361 11085 223389 11113
rect 223299 11023 223327 11051
rect 223361 11023 223389 11051
rect 223299 10961 223327 10989
rect 223361 10961 223389 10989
rect 233157 11147 233185 11175
rect 233219 11147 233247 11175
rect 233281 11147 233309 11175
rect 233343 11147 233371 11175
rect 233157 11085 233185 11113
rect 233219 11085 233247 11113
rect 233281 11085 233309 11113
rect 233343 11085 233371 11113
rect 233157 11023 233185 11051
rect 233219 11023 233247 11051
rect 233281 11023 233309 11051
rect 233343 11023 233371 11051
rect 233157 10961 233185 10989
rect 233219 10961 233247 10989
rect 233281 10961 233309 10989
rect 233343 10961 233371 10989
rect 219657 5147 219685 5175
rect 219719 5147 219747 5175
rect 219781 5147 219809 5175
rect 219843 5147 219871 5175
rect 219657 5085 219685 5113
rect 219719 5085 219747 5113
rect 219781 5085 219809 5113
rect 219843 5085 219871 5113
rect 219657 5023 219685 5051
rect 219719 5023 219747 5051
rect 219781 5023 219809 5051
rect 219843 5023 219871 5051
rect 219657 4961 219685 4989
rect 219719 4961 219747 4989
rect 219781 4961 219809 4989
rect 219843 4961 219871 4989
rect 230979 5147 231007 5175
rect 231041 5147 231069 5175
rect 230979 5085 231007 5113
rect 231041 5085 231069 5113
rect 230979 5023 231007 5051
rect 231041 5023 231069 5051
rect 230979 4961 231007 4989
rect 231041 4961 231069 4989
rect 219657 -588 219685 -560
rect 219719 -588 219747 -560
rect 219781 -588 219809 -560
rect 219843 -588 219871 -560
rect 219657 -650 219685 -622
rect 219719 -650 219747 -622
rect 219781 -650 219809 -622
rect 219843 -650 219871 -622
rect 219657 -712 219685 -684
rect 219719 -712 219747 -684
rect 219781 -712 219809 -684
rect 219843 -712 219871 -684
rect 219657 -774 219685 -746
rect 219719 -774 219747 -746
rect 219781 -774 219809 -746
rect 219843 -774 219871 -746
rect 233157 2147 233185 2175
rect 233219 2147 233247 2175
rect 233281 2147 233309 2175
rect 233343 2147 233371 2175
rect 233157 2085 233185 2113
rect 233219 2085 233247 2113
rect 233281 2085 233309 2113
rect 233343 2085 233371 2113
rect 233157 2023 233185 2051
rect 233219 2023 233247 2051
rect 233281 2023 233309 2051
rect 233343 2023 233371 2051
rect 233157 1961 233185 1989
rect 233219 1961 233247 1989
rect 233281 1961 233309 1989
rect 233343 1961 233371 1989
rect 233157 -108 233185 -80
rect 233219 -108 233247 -80
rect 233281 -108 233309 -80
rect 233343 -108 233371 -80
rect 233157 -170 233185 -142
rect 233219 -170 233247 -142
rect 233281 -170 233309 -142
rect 233343 -170 233371 -142
rect 233157 -232 233185 -204
rect 233219 -232 233247 -204
rect 233281 -232 233309 -204
rect 233343 -232 233371 -204
rect 233157 -294 233185 -266
rect 233219 -294 233247 -266
rect 233281 -294 233309 -266
rect 233343 -294 233371 -266
rect 235017 299058 235045 299086
rect 235079 299058 235107 299086
rect 235141 299058 235169 299086
rect 235203 299058 235231 299086
rect 235017 298996 235045 299024
rect 235079 298996 235107 299024
rect 235141 298996 235169 299024
rect 235203 298996 235231 299024
rect 235017 298934 235045 298962
rect 235079 298934 235107 298962
rect 235141 298934 235169 298962
rect 235203 298934 235231 298962
rect 235017 298872 235045 298900
rect 235079 298872 235107 298900
rect 235141 298872 235169 298900
rect 235203 298872 235231 298900
rect 235017 293147 235045 293175
rect 235079 293147 235107 293175
rect 235141 293147 235169 293175
rect 235203 293147 235231 293175
rect 235017 293085 235045 293113
rect 235079 293085 235107 293113
rect 235141 293085 235169 293113
rect 235203 293085 235231 293113
rect 235017 293023 235045 293051
rect 235079 293023 235107 293051
rect 235141 293023 235169 293051
rect 235203 293023 235231 293051
rect 235017 292961 235045 292989
rect 235079 292961 235107 292989
rect 235141 292961 235169 292989
rect 235203 292961 235231 292989
rect 235017 284147 235045 284175
rect 235079 284147 235107 284175
rect 235141 284147 235169 284175
rect 235203 284147 235231 284175
rect 235017 284085 235045 284113
rect 235079 284085 235107 284113
rect 235141 284085 235169 284113
rect 235203 284085 235231 284113
rect 235017 284023 235045 284051
rect 235079 284023 235107 284051
rect 235141 284023 235169 284051
rect 235203 284023 235231 284051
rect 235017 283961 235045 283989
rect 235079 283961 235107 283989
rect 235141 283961 235169 283989
rect 235203 283961 235231 283989
rect 235017 275147 235045 275175
rect 235079 275147 235107 275175
rect 235141 275147 235169 275175
rect 235203 275147 235231 275175
rect 235017 275085 235045 275113
rect 235079 275085 235107 275113
rect 235141 275085 235169 275113
rect 235203 275085 235231 275113
rect 235017 275023 235045 275051
rect 235079 275023 235107 275051
rect 235141 275023 235169 275051
rect 235203 275023 235231 275051
rect 235017 274961 235045 274989
rect 235079 274961 235107 274989
rect 235141 274961 235169 274989
rect 235203 274961 235231 274989
rect 235017 266147 235045 266175
rect 235079 266147 235107 266175
rect 235141 266147 235169 266175
rect 235203 266147 235231 266175
rect 235017 266085 235045 266113
rect 235079 266085 235107 266113
rect 235141 266085 235169 266113
rect 235203 266085 235231 266113
rect 235017 266023 235045 266051
rect 235079 266023 235107 266051
rect 235141 266023 235169 266051
rect 235203 266023 235231 266051
rect 235017 265961 235045 265989
rect 235079 265961 235107 265989
rect 235141 265961 235169 265989
rect 235203 265961 235231 265989
rect 235017 257147 235045 257175
rect 235079 257147 235107 257175
rect 235141 257147 235169 257175
rect 235203 257147 235231 257175
rect 235017 257085 235045 257113
rect 235079 257085 235107 257113
rect 235141 257085 235169 257113
rect 235203 257085 235231 257113
rect 235017 257023 235045 257051
rect 235079 257023 235107 257051
rect 235141 257023 235169 257051
rect 235203 257023 235231 257051
rect 235017 256961 235045 256989
rect 235079 256961 235107 256989
rect 235141 256961 235169 256989
rect 235203 256961 235231 256989
rect 235017 248147 235045 248175
rect 235079 248147 235107 248175
rect 235141 248147 235169 248175
rect 235203 248147 235231 248175
rect 235017 248085 235045 248113
rect 235079 248085 235107 248113
rect 235141 248085 235169 248113
rect 235203 248085 235231 248113
rect 235017 248023 235045 248051
rect 235079 248023 235107 248051
rect 235141 248023 235169 248051
rect 235203 248023 235231 248051
rect 235017 247961 235045 247989
rect 235079 247961 235107 247989
rect 235141 247961 235169 247989
rect 235203 247961 235231 247989
rect 235017 239147 235045 239175
rect 235079 239147 235107 239175
rect 235141 239147 235169 239175
rect 235203 239147 235231 239175
rect 235017 239085 235045 239113
rect 235079 239085 235107 239113
rect 235141 239085 235169 239113
rect 235203 239085 235231 239113
rect 235017 239023 235045 239051
rect 235079 239023 235107 239051
rect 235141 239023 235169 239051
rect 235203 239023 235231 239051
rect 235017 238961 235045 238989
rect 235079 238961 235107 238989
rect 235141 238961 235169 238989
rect 235203 238961 235231 238989
rect 235017 230147 235045 230175
rect 235079 230147 235107 230175
rect 235141 230147 235169 230175
rect 235203 230147 235231 230175
rect 235017 230085 235045 230113
rect 235079 230085 235107 230113
rect 235141 230085 235169 230113
rect 235203 230085 235231 230113
rect 235017 230023 235045 230051
rect 235079 230023 235107 230051
rect 235141 230023 235169 230051
rect 235203 230023 235231 230051
rect 235017 229961 235045 229989
rect 235079 229961 235107 229989
rect 235141 229961 235169 229989
rect 235203 229961 235231 229989
rect 235017 221147 235045 221175
rect 235079 221147 235107 221175
rect 235141 221147 235169 221175
rect 235203 221147 235231 221175
rect 235017 221085 235045 221113
rect 235079 221085 235107 221113
rect 235141 221085 235169 221113
rect 235203 221085 235231 221113
rect 235017 221023 235045 221051
rect 235079 221023 235107 221051
rect 235141 221023 235169 221051
rect 235203 221023 235231 221051
rect 235017 220961 235045 220989
rect 235079 220961 235107 220989
rect 235141 220961 235169 220989
rect 235203 220961 235231 220989
rect 235017 212147 235045 212175
rect 235079 212147 235107 212175
rect 235141 212147 235169 212175
rect 235203 212147 235231 212175
rect 235017 212085 235045 212113
rect 235079 212085 235107 212113
rect 235141 212085 235169 212113
rect 235203 212085 235231 212113
rect 235017 212023 235045 212051
rect 235079 212023 235107 212051
rect 235141 212023 235169 212051
rect 235203 212023 235231 212051
rect 235017 211961 235045 211989
rect 235079 211961 235107 211989
rect 235141 211961 235169 211989
rect 235203 211961 235231 211989
rect 235017 203147 235045 203175
rect 235079 203147 235107 203175
rect 235141 203147 235169 203175
rect 235203 203147 235231 203175
rect 235017 203085 235045 203113
rect 235079 203085 235107 203113
rect 235141 203085 235169 203113
rect 235203 203085 235231 203113
rect 235017 203023 235045 203051
rect 235079 203023 235107 203051
rect 235141 203023 235169 203051
rect 235203 203023 235231 203051
rect 235017 202961 235045 202989
rect 235079 202961 235107 202989
rect 235141 202961 235169 202989
rect 235203 202961 235231 202989
rect 235017 194147 235045 194175
rect 235079 194147 235107 194175
rect 235141 194147 235169 194175
rect 235203 194147 235231 194175
rect 235017 194085 235045 194113
rect 235079 194085 235107 194113
rect 235141 194085 235169 194113
rect 235203 194085 235231 194113
rect 235017 194023 235045 194051
rect 235079 194023 235107 194051
rect 235141 194023 235169 194051
rect 235203 194023 235231 194051
rect 235017 193961 235045 193989
rect 235079 193961 235107 193989
rect 235141 193961 235169 193989
rect 235203 193961 235231 193989
rect 235017 185147 235045 185175
rect 235079 185147 235107 185175
rect 235141 185147 235169 185175
rect 235203 185147 235231 185175
rect 235017 185085 235045 185113
rect 235079 185085 235107 185113
rect 235141 185085 235169 185113
rect 235203 185085 235231 185113
rect 235017 185023 235045 185051
rect 235079 185023 235107 185051
rect 235141 185023 235169 185051
rect 235203 185023 235231 185051
rect 235017 184961 235045 184989
rect 235079 184961 235107 184989
rect 235141 184961 235169 184989
rect 235203 184961 235231 184989
rect 235017 176147 235045 176175
rect 235079 176147 235107 176175
rect 235141 176147 235169 176175
rect 235203 176147 235231 176175
rect 235017 176085 235045 176113
rect 235079 176085 235107 176113
rect 235141 176085 235169 176113
rect 235203 176085 235231 176113
rect 235017 176023 235045 176051
rect 235079 176023 235107 176051
rect 235141 176023 235169 176051
rect 235203 176023 235231 176051
rect 235017 175961 235045 175989
rect 235079 175961 235107 175989
rect 235141 175961 235169 175989
rect 235203 175961 235231 175989
rect 248517 298578 248545 298606
rect 248579 298578 248607 298606
rect 248641 298578 248669 298606
rect 248703 298578 248731 298606
rect 248517 298516 248545 298544
rect 248579 298516 248607 298544
rect 248641 298516 248669 298544
rect 248703 298516 248731 298544
rect 248517 298454 248545 298482
rect 248579 298454 248607 298482
rect 248641 298454 248669 298482
rect 248703 298454 248731 298482
rect 248517 298392 248545 298420
rect 248579 298392 248607 298420
rect 248641 298392 248669 298420
rect 248703 298392 248731 298420
rect 248517 290147 248545 290175
rect 248579 290147 248607 290175
rect 248641 290147 248669 290175
rect 248703 290147 248731 290175
rect 248517 290085 248545 290113
rect 248579 290085 248607 290113
rect 248641 290085 248669 290113
rect 248703 290085 248731 290113
rect 248517 290023 248545 290051
rect 248579 290023 248607 290051
rect 248641 290023 248669 290051
rect 248703 290023 248731 290051
rect 248517 289961 248545 289989
rect 248579 289961 248607 289989
rect 248641 289961 248669 289989
rect 248703 289961 248731 289989
rect 248517 281147 248545 281175
rect 248579 281147 248607 281175
rect 248641 281147 248669 281175
rect 248703 281147 248731 281175
rect 248517 281085 248545 281113
rect 248579 281085 248607 281113
rect 248641 281085 248669 281113
rect 248703 281085 248731 281113
rect 248517 281023 248545 281051
rect 248579 281023 248607 281051
rect 248641 281023 248669 281051
rect 248703 281023 248731 281051
rect 248517 280961 248545 280989
rect 248579 280961 248607 280989
rect 248641 280961 248669 280989
rect 248703 280961 248731 280989
rect 248517 272147 248545 272175
rect 248579 272147 248607 272175
rect 248641 272147 248669 272175
rect 248703 272147 248731 272175
rect 248517 272085 248545 272113
rect 248579 272085 248607 272113
rect 248641 272085 248669 272113
rect 248703 272085 248731 272113
rect 248517 272023 248545 272051
rect 248579 272023 248607 272051
rect 248641 272023 248669 272051
rect 248703 272023 248731 272051
rect 248517 271961 248545 271989
rect 248579 271961 248607 271989
rect 248641 271961 248669 271989
rect 248703 271961 248731 271989
rect 248517 263147 248545 263175
rect 248579 263147 248607 263175
rect 248641 263147 248669 263175
rect 248703 263147 248731 263175
rect 248517 263085 248545 263113
rect 248579 263085 248607 263113
rect 248641 263085 248669 263113
rect 248703 263085 248731 263113
rect 248517 263023 248545 263051
rect 248579 263023 248607 263051
rect 248641 263023 248669 263051
rect 248703 263023 248731 263051
rect 248517 262961 248545 262989
rect 248579 262961 248607 262989
rect 248641 262961 248669 262989
rect 248703 262961 248731 262989
rect 248517 254147 248545 254175
rect 248579 254147 248607 254175
rect 248641 254147 248669 254175
rect 248703 254147 248731 254175
rect 248517 254085 248545 254113
rect 248579 254085 248607 254113
rect 248641 254085 248669 254113
rect 248703 254085 248731 254113
rect 248517 254023 248545 254051
rect 248579 254023 248607 254051
rect 248641 254023 248669 254051
rect 248703 254023 248731 254051
rect 248517 253961 248545 253989
rect 248579 253961 248607 253989
rect 248641 253961 248669 253989
rect 248703 253961 248731 253989
rect 248517 245147 248545 245175
rect 248579 245147 248607 245175
rect 248641 245147 248669 245175
rect 248703 245147 248731 245175
rect 248517 245085 248545 245113
rect 248579 245085 248607 245113
rect 248641 245085 248669 245113
rect 248703 245085 248731 245113
rect 248517 245023 248545 245051
rect 248579 245023 248607 245051
rect 248641 245023 248669 245051
rect 248703 245023 248731 245051
rect 248517 244961 248545 244989
rect 248579 244961 248607 244989
rect 248641 244961 248669 244989
rect 248703 244961 248731 244989
rect 248517 236147 248545 236175
rect 248579 236147 248607 236175
rect 248641 236147 248669 236175
rect 248703 236147 248731 236175
rect 248517 236085 248545 236113
rect 248579 236085 248607 236113
rect 248641 236085 248669 236113
rect 248703 236085 248731 236113
rect 248517 236023 248545 236051
rect 248579 236023 248607 236051
rect 248641 236023 248669 236051
rect 248703 236023 248731 236051
rect 248517 235961 248545 235989
rect 248579 235961 248607 235989
rect 248641 235961 248669 235989
rect 248703 235961 248731 235989
rect 248517 227147 248545 227175
rect 248579 227147 248607 227175
rect 248641 227147 248669 227175
rect 248703 227147 248731 227175
rect 248517 227085 248545 227113
rect 248579 227085 248607 227113
rect 248641 227085 248669 227113
rect 248703 227085 248731 227113
rect 248517 227023 248545 227051
rect 248579 227023 248607 227051
rect 248641 227023 248669 227051
rect 248703 227023 248731 227051
rect 248517 226961 248545 226989
rect 248579 226961 248607 226989
rect 248641 226961 248669 226989
rect 248703 226961 248731 226989
rect 248517 218147 248545 218175
rect 248579 218147 248607 218175
rect 248641 218147 248669 218175
rect 248703 218147 248731 218175
rect 248517 218085 248545 218113
rect 248579 218085 248607 218113
rect 248641 218085 248669 218113
rect 248703 218085 248731 218113
rect 248517 218023 248545 218051
rect 248579 218023 248607 218051
rect 248641 218023 248669 218051
rect 248703 218023 248731 218051
rect 248517 217961 248545 217989
rect 248579 217961 248607 217989
rect 248641 217961 248669 217989
rect 248703 217961 248731 217989
rect 248517 209147 248545 209175
rect 248579 209147 248607 209175
rect 248641 209147 248669 209175
rect 248703 209147 248731 209175
rect 248517 209085 248545 209113
rect 248579 209085 248607 209113
rect 248641 209085 248669 209113
rect 248703 209085 248731 209113
rect 248517 209023 248545 209051
rect 248579 209023 248607 209051
rect 248641 209023 248669 209051
rect 248703 209023 248731 209051
rect 248517 208961 248545 208989
rect 248579 208961 248607 208989
rect 248641 208961 248669 208989
rect 248703 208961 248731 208989
rect 248517 200147 248545 200175
rect 248579 200147 248607 200175
rect 248641 200147 248669 200175
rect 248703 200147 248731 200175
rect 248517 200085 248545 200113
rect 248579 200085 248607 200113
rect 248641 200085 248669 200113
rect 248703 200085 248731 200113
rect 248517 200023 248545 200051
rect 248579 200023 248607 200051
rect 248641 200023 248669 200051
rect 248703 200023 248731 200051
rect 248517 199961 248545 199989
rect 248579 199961 248607 199989
rect 248641 199961 248669 199989
rect 248703 199961 248731 199989
rect 248517 191147 248545 191175
rect 248579 191147 248607 191175
rect 248641 191147 248669 191175
rect 248703 191147 248731 191175
rect 248517 191085 248545 191113
rect 248579 191085 248607 191113
rect 248641 191085 248669 191113
rect 248703 191085 248731 191113
rect 248517 191023 248545 191051
rect 248579 191023 248607 191051
rect 248641 191023 248669 191051
rect 248703 191023 248731 191051
rect 248517 190961 248545 190989
rect 248579 190961 248607 190989
rect 248641 190961 248669 190989
rect 248703 190961 248731 190989
rect 248517 182147 248545 182175
rect 248579 182147 248607 182175
rect 248641 182147 248669 182175
rect 248703 182147 248731 182175
rect 248517 182085 248545 182113
rect 248579 182085 248607 182113
rect 248641 182085 248669 182113
rect 248703 182085 248731 182113
rect 248517 182023 248545 182051
rect 248579 182023 248607 182051
rect 248641 182023 248669 182051
rect 248703 182023 248731 182051
rect 248517 181961 248545 181989
rect 248579 181961 248607 181989
rect 248641 181961 248669 181989
rect 248703 181961 248731 181989
rect 238659 173147 238687 173175
rect 238721 173147 238749 173175
rect 238659 173085 238687 173113
rect 238721 173085 238749 173113
rect 238659 173023 238687 173051
rect 238721 173023 238749 173051
rect 238659 172961 238687 172989
rect 238721 172961 238749 172989
rect 248517 173147 248545 173175
rect 248579 173147 248607 173175
rect 248641 173147 248669 173175
rect 248703 173147 248731 173175
rect 248517 173085 248545 173113
rect 248579 173085 248607 173113
rect 248641 173085 248669 173113
rect 248703 173085 248731 173113
rect 248517 173023 248545 173051
rect 248579 173023 248607 173051
rect 248641 173023 248669 173051
rect 248703 173023 248731 173051
rect 248517 172961 248545 172989
rect 248579 172961 248607 172989
rect 248641 172961 248669 172989
rect 248703 172961 248731 172989
rect 235017 167147 235045 167175
rect 235079 167147 235107 167175
rect 235141 167147 235169 167175
rect 235203 167147 235231 167175
rect 235017 167085 235045 167113
rect 235079 167085 235107 167113
rect 235141 167085 235169 167113
rect 235203 167085 235231 167113
rect 235017 167023 235045 167051
rect 235079 167023 235107 167051
rect 235141 167023 235169 167051
rect 235203 167023 235231 167051
rect 235017 166961 235045 166989
rect 235079 166961 235107 166989
rect 235141 166961 235169 166989
rect 235203 166961 235231 166989
rect 246339 167147 246367 167175
rect 246401 167147 246429 167175
rect 246339 167085 246367 167113
rect 246401 167085 246429 167113
rect 246339 167023 246367 167051
rect 246401 167023 246429 167051
rect 246339 166961 246367 166989
rect 246401 166961 246429 166989
rect 238659 164147 238687 164175
rect 238721 164147 238749 164175
rect 238659 164085 238687 164113
rect 238721 164085 238749 164113
rect 238659 164023 238687 164051
rect 238721 164023 238749 164051
rect 238659 163961 238687 163989
rect 238721 163961 238749 163989
rect 248517 164147 248545 164175
rect 248579 164147 248607 164175
rect 248641 164147 248669 164175
rect 248703 164147 248731 164175
rect 248517 164085 248545 164113
rect 248579 164085 248607 164113
rect 248641 164085 248669 164113
rect 248703 164085 248731 164113
rect 248517 164023 248545 164051
rect 248579 164023 248607 164051
rect 248641 164023 248669 164051
rect 248703 164023 248731 164051
rect 248517 163961 248545 163989
rect 248579 163961 248607 163989
rect 248641 163961 248669 163989
rect 248703 163961 248731 163989
rect 235017 158147 235045 158175
rect 235079 158147 235107 158175
rect 235141 158147 235169 158175
rect 235203 158147 235231 158175
rect 235017 158085 235045 158113
rect 235079 158085 235107 158113
rect 235141 158085 235169 158113
rect 235203 158085 235231 158113
rect 235017 158023 235045 158051
rect 235079 158023 235107 158051
rect 235141 158023 235169 158051
rect 235203 158023 235231 158051
rect 235017 157961 235045 157989
rect 235079 157961 235107 157989
rect 235141 157961 235169 157989
rect 235203 157961 235231 157989
rect 246339 158147 246367 158175
rect 246401 158147 246429 158175
rect 246339 158085 246367 158113
rect 246401 158085 246429 158113
rect 246339 158023 246367 158051
rect 246401 158023 246429 158051
rect 246339 157961 246367 157989
rect 246401 157961 246429 157989
rect 238659 155147 238687 155175
rect 238721 155147 238749 155175
rect 238659 155085 238687 155113
rect 238721 155085 238749 155113
rect 238659 155023 238687 155051
rect 238721 155023 238749 155051
rect 238659 154961 238687 154989
rect 238721 154961 238749 154989
rect 248517 155147 248545 155175
rect 248579 155147 248607 155175
rect 248641 155147 248669 155175
rect 248703 155147 248731 155175
rect 248517 155085 248545 155113
rect 248579 155085 248607 155113
rect 248641 155085 248669 155113
rect 248703 155085 248731 155113
rect 248517 155023 248545 155051
rect 248579 155023 248607 155051
rect 248641 155023 248669 155051
rect 248703 155023 248731 155051
rect 248517 154961 248545 154989
rect 248579 154961 248607 154989
rect 248641 154961 248669 154989
rect 248703 154961 248731 154989
rect 235017 149147 235045 149175
rect 235079 149147 235107 149175
rect 235141 149147 235169 149175
rect 235203 149147 235231 149175
rect 235017 149085 235045 149113
rect 235079 149085 235107 149113
rect 235141 149085 235169 149113
rect 235203 149085 235231 149113
rect 235017 149023 235045 149051
rect 235079 149023 235107 149051
rect 235141 149023 235169 149051
rect 235203 149023 235231 149051
rect 235017 148961 235045 148989
rect 235079 148961 235107 148989
rect 235141 148961 235169 148989
rect 235203 148961 235231 148989
rect 246339 149147 246367 149175
rect 246401 149147 246429 149175
rect 246339 149085 246367 149113
rect 246401 149085 246429 149113
rect 246339 149023 246367 149051
rect 246401 149023 246429 149051
rect 246339 148961 246367 148989
rect 246401 148961 246429 148989
rect 238659 146147 238687 146175
rect 238721 146147 238749 146175
rect 238659 146085 238687 146113
rect 238721 146085 238749 146113
rect 238659 146023 238687 146051
rect 238721 146023 238749 146051
rect 238659 145961 238687 145989
rect 238721 145961 238749 145989
rect 248517 146147 248545 146175
rect 248579 146147 248607 146175
rect 248641 146147 248669 146175
rect 248703 146147 248731 146175
rect 248517 146085 248545 146113
rect 248579 146085 248607 146113
rect 248641 146085 248669 146113
rect 248703 146085 248731 146113
rect 248517 146023 248545 146051
rect 248579 146023 248607 146051
rect 248641 146023 248669 146051
rect 248703 146023 248731 146051
rect 248517 145961 248545 145989
rect 248579 145961 248607 145989
rect 248641 145961 248669 145989
rect 248703 145961 248731 145989
rect 235017 140147 235045 140175
rect 235079 140147 235107 140175
rect 235141 140147 235169 140175
rect 235203 140147 235231 140175
rect 235017 140085 235045 140113
rect 235079 140085 235107 140113
rect 235141 140085 235169 140113
rect 235203 140085 235231 140113
rect 235017 140023 235045 140051
rect 235079 140023 235107 140051
rect 235141 140023 235169 140051
rect 235203 140023 235231 140051
rect 235017 139961 235045 139989
rect 235079 139961 235107 139989
rect 235141 139961 235169 139989
rect 235203 139961 235231 139989
rect 246339 140147 246367 140175
rect 246401 140147 246429 140175
rect 246339 140085 246367 140113
rect 246401 140085 246429 140113
rect 246339 140023 246367 140051
rect 246401 140023 246429 140051
rect 246339 139961 246367 139989
rect 246401 139961 246429 139989
rect 238659 137147 238687 137175
rect 238721 137147 238749 137175
rect 238659 137085 238687 137113
rect 238721 137085 238749 137113
rect 238659 137023 238687 137051
rect 238721 137023 238749 137051
rect 238659 136961 238687 136989
rect 238721 136961 238749 136989
rect 248517 137147 248545 137175
rect 248579 137147 248607 137175
rect 248641 137147 248669 137175
rect 248703 137147 248731 137175
rect 248517 137085 248545 137113
rect 248579 137085 248607 137113
rect 248641 137085 248669 137113
rect 248703 137085 248731 137113
rect 248517 137023 248545 137051
rect 248579 137023 248607 137051
rect 248641 137023 248669 137051
rect 248703 137023 248731 137051
rect 248517 136961 248545 136989
rect 248579 136961 248607 136989
rect 248641 136961 248669 136989
rect 248703 136961 248731 136989
rect 235017 131147 235045 131175
rect 235079 131147 235107 131175
rect 235141 131147 235169 131175
rect 235203 131147 235231 131175
rect 235017 131085 235045 131113
rect 235079 131085 235107 131113
rect 235141 131085 235169 131113
rect 235203 131085 235231 131113
rect 235017 131023 235045 131051
rect 235079 131023 235107 131051
rect 235141 131023 235169 131051
rect 235203 131023 235231 131051
rect 235017 130961 235045 130989
rect 235079 130961 235107 130989
rect 235141 130961 235169 130989
rect 235203 130961 235231 130989
rect 246339 131147 246367 131175
rect 246401 131147 246429 131175
rect 246339 131085 246367 131113
rect 246401 131085 246429 131113
rect 246339 131023 246367 131051
rect 246401 131023 246429 131051
rect 246339 130961 246367 130989
rect 246401 130961 246429 130989
rect 238659 128147 238687 128175
rect 238721 128147 238749 128175
rect 238659 128085 238687 128113
rect 238721 128085 238749 128113
rect 238659 128023 238687 128051
rect 238721 128023 238749 128051
rect 238659 127961 238687 127989
rect 238721 127961 238749 127989
rect 248517 128147 248545 128175
rect 248579 128147 248607 128175
rect 248641 128147 248669 128175
rect 248703 128147 248731 128175
rect 248517 128085 248545 128113
rect 248579 128085 248607 128113
rect 248641 128085 248669 128113
rect 248703 128085 248731 128113
rect 248517 128023 248545 128051
rect 248579 128023 248607 128051
rect 248641 128023 248669 128051
rect 248703 128023 248731 128051
rect 248517 127961 248545 127989
rect 248579 127961 248607 127989
rect 248641 127961 248669 127989
rect 248703 127961 248731 127989
rect 235017 122147 235045 122175
rect 235079 122147 235107 122175
rect 235141 122147 235169 122175
rect 235203 122147 235231 122175
rect 235017 122085 235045 122113
rect 235079 122085 235107 122113
rect 235141 122085 235169 122113
rect 235203 122085 235231 122113
rect 235017 122023 235045 122051
rect 235079 122023 235107 122051
rect 235141 122023 235169 122051
rect 235203 122023 235231 122051
rect 235017 121961 235045 121989
rect 235079 121961 235107 121989
rect 235141 121961 235169 121989
rect 235203 121961 235231 121989
rect 246339 122147 246367 122175
rect 246401 122147 246429 122175
rect 246339 122085 246367 122113
rect 246401 122085 246429 122113
rect 246339 122023 246367 122051
rect 246401 122023 246429 122051
rect 246339 121961 246367 121989
rect 246401 121961 246429 121989
rect 238659 119147 238687 119175
rect 238721 119147 238749 119175
rect 238659 119085 238687 119113
rect 238721 119085 238749 119113
rect 238659 119023 238687 119051
rect 238721 119023 238749 119051
rect 238659 118961 238687 118989
rect 238721 118961 238749 118989
rect 248517 119147 248545 119175
rect 248579 119147 248607 119175
rect 248641 119147 248669 119175
rect 248703 119147 248731 119175
rect 248517 119085 248545 119113
rect 248579 119085 248607 119113
rect 248641 119085 248669 119113
rect 248703 119085 248731 119113
rect 248517 119023 248545 119051
rect 248579 119023 248607 119051
rect 248641 119023 248669 119051
rect 248703 119023 248731 119051
rect 248517 118961 248545 118989
rect 248579 118961 248607 118989
rect 248641 118961 248669 118989
rect 248703 118961 248731 118989
rect 235017 113147 235045 113175
rect 235079 113147 235107 113175
rect 235141 113147 235169 113175
rect 235203 113147 235231 113175
rect 235017 113085 235045 113113
rect 235079 113085 235107 113113
rect 235141 113085 235169 113113
rect 235203 113085 235231 113113
rect 235017 113023 235045 113051
rect 235079 113023 235107 113051
rect 235141 113023 235169 113051
rect 235203 113023 235231 113051
rect 235017 112961 235045 112989
rect 235079 112961 235107 112989
rect 235141 112961 235169 112989
rect 235203 112961 235231 112989
rect 246339 113147 246367 113175
rect 246401 113147 246429 113175
rect 246339 113085 246367 113113
rect 246401 113085 246429 113113
rect 246339 113023 246367 113051
rect 246401 113023 246429 113051
rect 246339 112961 246367 112989
rect 246401 112961 246429 112989
rect 238659 110147 238687 110175
rect 238721 110147 238749 110175
rect 238659 110085 238687 110113
rect 238721 110085 238749 110113
rect 238659 110023 238687 110051
rect 238721 110023 238749 110051
rect 238659 109961 238687 109989
rect 238721 109961 238749 109989
rect 248517 110147 248545 110175
rect 248579 110147 248607 110175
rect 248641 110147 248669 110175
rect 248703 110147 248731 110175
rect 248517 110085 248545 110113
rect 248579 110085 248607 110113
rect 248641 110085 248669 110113
rect 248703 110085 248731 110113
rect 248517 110023 248545 110051
rect 248579 110023 248607 110051
rect 248641 110023 248669 110051
rect 248703 110023 248731 110051
rect 248517 109961 248545 109989
rect 248579 109961 248607 109989
rect 248641 109961 248669 109989
rect 248703 109961 248731 109989
rect 235017 104147 235045 104175
rect 235079 104147 235107 104175
rect 235141 104147 235169 104175
rect 235203 104147 235231 104175
rect 235017 104085 235045 104113
rect 235079 104085 235107 104113
rect 235141 104085 235169 104113
rect 235203 104085 235231 104113
rect 235017 104023 235045 104051
rect 235079 104023 235107 104051
rect 235141 104023 235169 104051
rect 235203 104023 235231 104051
rect 235017 103961 235045 103989
rect 235079 103961 235107 103989
rect 235141 103961 235169 103989
rect 235203 103961 235231 103989
rect 246339 104147 246367 104175
rect 246401 104147 246429 104175
rect 246339 104085 246367 104113
rect 246401 104085 246429 104113
rect 246339 104023 246367 104051
rect 246401 104023 246429 104051
rect 246339 103961 246367 103989
rect 246401 103961 246429 103989
rect 238659 101147 238687 101175
rect 238721 101147 238749 101175
rect 238659 101085 238687 101113
rect 238721 101085 238749 101113
rect 238659 101023 238687 101051
rect 238721 101023 238749 101051
rect 238659 100961 238687 100989
rect 238721 100961 238749 100989
rect 248517 101147 248545 101175
rect 248579 101147 248607 101175
rect 248641 101147 248669 101175
rect 248703 101147 248731 101175
rect 248517 101085 248545 101113
rect 248579 101085 248607 101113
rect 248641 101085 248669 101113
rect 248703 101085 248731 101113
rect 248517 101023 248545 101051
rect 248579 101023 248607 101051
rect 248641 101023 248669 101051
rect 248703 101023 248731 101051
rect 248517 100961 248545 100989
rect 248579 100961 248607 100989
rect 248641 100961 248669 100989
rect 248703 100961 248731 100989
rect 235017 95147 235045 95175
rect 235079 95147 235107 95175
rect 235141 95147 235169 95175
rect 235203 95147 235231 95175
rect 235017 95085 235045 95113
rect 235079 95085 235107 95113
rect 235141 95085 235169 95113
rect 235203 95085 235231 95113
rect 235017 95023 235045 95051
rect 235079 95023 235107 95051
rect 235141 95023 235169 95051
rect 235203 95023 235231 95051
rect 235017 94961 235045 94989
rect 235079 94961 235107 94989
rect 235141 94961 235169 94989
rect 235203 94961 235231 94989
rect 246339 95147 246367 95175
rect 246401 95147 246429 95175
rect 246339 95085 246367 95113
rect 246401 95085 246429 95113
rect 246339 95023 246367 95051
rect 246401 95023 246429 95051
rect 246339 94961 246367 94989
rect 246401 94961 246429 94989
rect 238659 92147 238687 92175
rect 238721 92147 238749 92175
rect 238659 92085 238687 92113
rect 238721 92085 238749 92113
rect 238659 92023 238687 92051
rect 238721 92023 238749 92051
rect 238659 91961 238687 91989
rect 238721 91961 238749 91989
rect 248517 92147 248545 92175
rect 248579 92147 248607 92175
rect 248641 92147 248669 92175
rect 248703 92147 248731 92175
rect 248517 92085 248545 92113
rect 248579 92085 248607 92113
rect 248641 92085 248669 92113
rect 248703 92085 248731 92113
rect 248517 92023 248545 92051
rect 248579 92023 248607 92051
rect 248641 92023 248669 92051
rect 248703 92023 248731 92051
rect 248517 91961 248545 91989
rect 248579 91961 248607 91989
rect 248641 91961 248669 91989
rect 248703 91961 248731 91989
rect 235017 86147 235045 86175
rect 235079 86147 235107 86175
rect 235141 86147 235169 86175
rect 235203 86147 235231 86175
rect 235017 86085 235045 86113
rect 235079 86085 235107 86113
rect 235141 86085 235169 86113
rect 235203 86085 235231 86113
rect 235017 86023 235045 86051
rect 235079 86023 235107 86051
rect 235141 86023 235169 86051
rect 235203 86023 235231 86051
rect 235017 85961 235045 85989
rect 235079 85961 235107 85989
rect 235141 85961 235169 85989
rect 235203 85961 235231 85989
rect 246339 86147 246367 86175
rect 246401 86147 246429 86175
rect 246339 86085 246367 86113
rect 246401 86085 246429 86113
rect 246339 86023 246367 86051
rect 246401 86023 246429 86051
rect 246339 85961 246367 85989
rect 246401 85961 246429 85989
rect 238659 83147 238687 83175
rect 238721 83147 238749 83175
rect 238659 83085 238687 83113
rect 238721 83085 238749 83113
rect 238659 83023 238687 83051
rect 238721 83023 238749 83051
rect 238659 82961 238687 82989
rect 238721 82961 238749 82989
rect 248517 83147 248545 83175
rect 248579 83147 248607 83175
rect 248641 83147 248669 83175
rect 248703 83147 248731 83175
rect 248517 83085 248545 83113
rect 248579 83085 248607 83113
rect 248641 83085 248669 83113
rect 248703 83085 248731 83113
rect 248517 83023 248545 83051
rect 248579 83023 248607 83051
rect 248641 83023 248669 83051
rect 248703 83023 248731 83051
rect 248517 82961 248545 82989
rect 248579 82961 248607 82989
rect 248641 82961 248669 82989
rect 248703 82961 248731 82989
rect 235017 77147 235045 77175
rect 235079 77147 235107 77175
rect 235141 77147 235169 77175
rect 235203 77147 235231 77175
rect 235017 77085 235045 77113
rect 235079 77085 235107 77113
rect 235141 77085 235169 77113
rect 235203 77085 235231 77113
rect 235017 77023 235045 77051
rect 235079 77023 235107 77051
rect 235141 77023 235169 77051
rect 235203 77023 235231 77051
rect 235017 76961 235045 76989
rect 235079 76961 235107 76989
rect 235141 76961 235169 76989
rect 235203 76961 235231 76989
rect 246339 77147 246367 77175
rect 246401 77147 246429 77175
rect 246339 77085 246367 77113
rect 246401 77085 246429 77113
rect 246339 77023 246367 77051
rect 246401 77023 246429 77051
rect 246339 76961 246367 76989
rect 246401 76961 246429 76989
rect 238659 74147 238687 74175
rect 238721 74147 238749 74175
rect 238659 74085 238687 74113
rect 238721 74085 238749 74113
rect 238659 74023 238687 74051
rect 238721 74023 238749 74051
rect 238659 73961 238687 73989
rect 238721 73961 238749 73989
rect 248517 74147 248545 74175
rect 248579 74147 248607 74175
rect 248641 74147 248669 74175
rect 248703 74147 248731 74175
rect 248517 74085 248545 74113
rect 248579 74085 248607 74113
rect 248641 74085 248669 74113
rect 248703 74085 248731 74113
rect 248517 74023 248545 74051
rect 248579 74023 248607 74051
rect 248641 74023 248669 74051
rect 248703 74023 248731 74051
rect 248517 73961 248545 73989
rect 248579 73961 248607 73989
rect 248641 73961 248669 73989
rect 248703 73961 248731 73989
rect 235017 68147 235045 68175
rect 235079 68147 235107 68175
rect 235141 68147 235169 68175
rect 235203 68147 235231 68175
rect 235017 68085 235045 68113
rect 235079 68085 235107 68113
rect 235141 68085 235169 68113
rect 235203 68085 235231 68113
rect 235017 68023 235045 68051
rect 235079 68023 235107 68051
rect 235141 68023 235169 68051
rect 235203 68023 235231 68051
rect 235017 67961 235045 67989
rect 235079 67961 235107 67989
rect 235141 67961 235169 67989
rect 235203 67961 235231 67989
rect 246339 68147 246367 68175
rect 246401 68147 246429 68175
rect 246339 68085 246367 68113
rect 246401 68085 246429 68113
rect 246339 68023 246367 68051
rect 246401 68023 246429 68051
rect 246339 67961 246367 67989
rect 246401 67961 246429 67989
rect 238659 65147 238687 65175
rect 238721 65147 238749 65175
rect 238659 65085 238687 65113
rect 238721 65085 238749 65113
rect 238659 65023 238687 65051
rect 238721 65023 238749 65051
rect 238659 64961 238687 64989
rect 238721 64961 238749 64989
rect 248517 65147 248545 65175
rect 248579 65147 248607 65175
rect 248641 65147 248669 65175
rect 248703 65147 248731 65175
rect 248517 65085 248545 65113
rect 248579 65085 248607 65113
rect 248641 65085 248669 65113
rect 248703 65085 248731 65113
rect 248517 65023 248545 65051
rect 248579 65023 248607 65051
rect 248641 65023 248669 65051
rect 248703 65023 248731 65051
rect 248517 64961 248545 64989
rect 248579 64961 248607 64989
rect 248641 64961 248669 64989
rect 248703 64961 248731 64989
rect 235017 59147 235045 59175
rect 235079 59147 235107 59175
rect 235141 59147 235169 59175
rect 235203 59147 235231 59175
rect 235017 59085 235045 59113
rect 235079 59085 235107 59113
rect 235141 59085 235169 59113
rect 235203 59085 235231 59113
rect 235017 59023 235045 59051
rect 235079 59023 235107 59051
rect 235141 59023 235169 59051
rect 235203 59023 235231 59051
rect 235017 58961 235045 58989
rect 235079 58961 235107 58989
rect 235141 58961 235169 58989
rect 235203 58961 235231 58989
rect 246339 59147 246367 59175
rect 246401 59147 246429 59175
rect 246339 59085 246367 59113
rect 246401 59085 246429 59113
rect 246339 59023 246367 59051
rect 246401 59023 246429 59051
rect 246339 58961 246367 58989
rect 246401 58961 246429 58989
rect 238659 56147 238687 56175
rect 238721 56147 238749 56175
rect 238659 56085 238687 56113
rect 238721 56085 238749 56113
rect 238659 56023 238687 56051
rect 238721 56023 238749 56051
rect 238659 55961 238687 55989
rect 238721 55961 238749 55989
rect 248517 56147 248545 56175
rect 248579 56147 248607 56175
rect 248641 56147 248669 56175
rect 248703 56147 248731 56175
rect 248517 56085 248545 56113
rect 248579 56085 248607 56113
rect 248641 56085 248669 56113
rect 248703 56085 248731 56113
rect 248517 56023 248545 56051
rect 248579 56023 248607 56051
rect 248641 56023 248669 56051
rect 248703 56023 248731 56051
rect 248517 55961 248545 55989
rect 248579 55961 248607 55989
rect 248641 55961 248669 55989
rect 248703 55961 248731 55989
rect 235017 50147 235045 50175
rect 235079 50147 235107 50175
rect 235141 50147 235169 50175
rect 235203 50147 235231 50175
rect 235017 50085 235045 50113
rect 235079 50085 235107 50113
rect 235141 50085 235169 50113
rect 235203 50085 235231 50113
rect 235017 50023 235045 50051
rect 235079 50023 235107 50051
rect 235141 50023 235169 50051
rect 235203 50023 235231 50051
rect 235017 49961 235045 49989
rect 235079 49961 235107 49989
rect 235141 49961 235169 49989
rect 235203 49961 235231 49989
rect 246339 50147 246367 50175
rect 246401 50147 246429 50175
rect 246339 50085 246367 50113
rect 246401 50085 246429 50113
rect 246339 50023 246367 50051
rect 246401 50023 246429 50051
rect 246339 49961 246367 49989
rect 246401 49961 246429 49989
rect 238659 47147 238687 47175
rect 238721 47147 238749 47175
rect 238659 47085 238687 47113
rect 238721 47085 238749 47113
rect 238659 47023 238687 47051
rect 238721 47023 238749 47051
rect 238659 46961 238687 46989
rect 238721 46961 238749 46989
rect 248517 47147 248545 47175
rect 248579 47147 248607 47175
rect 248641 47147 248669 47175
rect 248703 47147 248731 47175
rect 248517 47085 248545 47113
rect 248579 47085 248607 47113
rect 248641 47085 248669 47113
rect 248703 47085 248731 47113
rect 248517 47023 248545 47051
rect 248579 47023 248607 47051
rect 248641 47023 248669 47051
rect 248703 47023 248731 47051
rect 248517 46961 248545 46989
rect 248579 46961 248607 46989
rect 248641 46961 248669 46989
rect 248703 46961 248731 46989
rect 235017 41147 235045 41175
rect 235079 41147 235107 41175
rect 235141 41147 235169 41175
rect 235203 41147 235231 41175
rect 235017 41085 235045 41113
rect 235079 41085 235107 41113
rect 235141 41085 235169 41113
rect 235203 41085 235231 41113
rect 235017 41023 235045 41051
rect 235079 41023 235107 41051
rect 235141 41023 235169 41051
rect 235203 41023 235231 41051
rect 235017 40961 235045 40989
rect 235079 40961 235107 40989
rect 235141 40961 235169 40989
rect 235203 40961 235231 40989
rect 246339 41147 246367 41175
rect 246401 41147 246429 41175
rect 246339 41085 246367 41113
rect 246401 41085 246429 41113
rect 246339 41023 246367 41051
rect 246401 41023 246429 41051
rect 246339 40961 246367 40989
rect 246401 40961 246429 40989
rect 238659 38147 238687 38175
rect 238721 38147 238749 38175
rect 238659 38085 238687 38113
rect 238721 38085 238749 38113
rect 238659 38023 238687 38051
rect 238721 38023 238749 38051
rect 238659 37961 238687 37989
rect 238721 37961 238749 37989
rect 248517 38147 248545 38175
rect 248579 38147 248607 38175
rect 248641 38147 248669 38175
rect 248703 38147 248731 38175
rect 248517 38085 248545 38113
rect 248579 38085 248607 38113
rect 248641 38085 248669 38113
rect 248703 38085 248731 38113
rect 248517 38023 248545 38051
rect 248579 38023 248607 38051
rect 248641 38023 248669 38051
rect 248703 38023 248731 38051
rect 248517 37961 248545 37989
rect 248579 37961 248607 37989
rect 248641 37961 248669 37989
rect 248703 37961 248731 37989
rect 235017 32147 235045 32175
rect 235079 32147 235107 32175
rect 235141 32147 235169 32175
rect 235203 32147 235231 32175
rect 235017 32085 235045 32113
rect 235079 32085 235107 32113
rect 235141 32085 235169 32113
rect 235203 32085 235231 32113
rect 235017 32023 235045 32051
rect 235079 32023 235107 32051
rect 235141 32023 235169 32051
rect 235203 32023 235231 32051
rect 235017 31961 235045 31989
rect 235079 31961 235107 31989
rect 235141 31961 235169 31989
rect 235203 31961 235231 31989
rect 246339 32147 246367 32175
rect 246401 32147 246429 32175
rect 246339 32085 246367 32113
rect 246401 32085 246429 32113
rect 246339 32023 246367 32051
rect 246401 32023 246429 32051
rect 246339 31961 246367 31989
rect 246401 31961 246429 31989
rect 238659 29147 238687 29175
rect 238721 29147 238749 29175
rect 238659 29085 238687 29113
rect 238721 29085 238749 29113
rect 238659 29023 238687 29051
rect 238721 29023 238749 29051
rect 238659 28961 238687 28989
rect 238721 28961 238749 28989
rect 248517 29147 248545 29175
rect 248579 29147 248607 29175
rect 248641 29147 248669 29175
rect 248703 29147 248731 29175
rect 248517 29085 248545 29113
rect 248579 29085 248607 29113
rect 248641 29085 248669 29113
rect 248703 29085 248731 29113
rect 248517 29023 248545 29051
rect 248579 29023 248607 29051
rect 248641 29023 248669 29051
rect 248703 29023 248731 29051
rect 248517 28961 248545 28989
rect 248579 28961 248607 28989
rect 248641 28961 248669 28989
rect 248703 28961 248731 28989
rect 235017 23147 235045 23175
rect 235079 23147 235107 23175
rect 235141 23147 235169 23175
rect 235203 23147 235231 23175
rect 235017 23085 235045 23113
rect 235079 23085 235107 23113
rect 235141 23085 235169 23113
rect 235203 23085 235231 23113
rect 235017 23023 235045 23051
rect 235079 23023 235107 23051
rect 235141 23023 235169 23051
rect 235203 23023 235231 23051
rect 235017 22961 235045 22989
rect 235079 22961 235107 22989
rect 235141 22961 235169 22989
rect 235203 22961 235231 22989
rect 246339 23147 246367 23175
rect 246401 23147 246429 23175
rect 246339 23085 246367 23113
rect 246401 23085 246429 23113
rect 246339 23023 246367 23051
rect 246401 23023 246429 23051
rect 246339 22961 246367 22989
rect 246401 22961 246429 22989
rect 238659 20147 238687 20175
rect 238721 20147 238749 20175
rect 238659 20085 238687 20113
rect 238721 20085 238749 20113
rect 238659 20023 238687 20051
rect 238721 20023 238749 20051
rect 238659 19961 238687 19989
rect 238721 19961 238749 19989
rect 248517 20147 248545 20175
rect 248579 20147 248607 20175
rect 248641 20147 248669 20175
rect 248703 20147 248731 20175
rect 248517 20085 248545 20113
rect 248579 20085 248607 20113
rect 248641 20085 248669 20113
rect 248703 20085 248731 20113
rect 248517 20023 248545 20051
rect 248579 20023 248607 20051
rect 248641 20023 248669 20051
rect 248703 20023 248731 20051
rect 248517 19961 248545 19989
rect 248579 19961 248607 19989
rect 248641 19961 248669 19989
rect 248703 19961 248731 19989
rect 235017 14147 235045 14175
rect 235079 14147 235107 14175
rect 235141 14147 235169 14175
rect 235203 14147 235231 14175
rect 235017 14085 235045 14113
rect 235079 14085 235107 14113
rect 235141 14085 235169 14113
rect 235203 14085 235231 14113
rect 235017 14023 235045 14051
rect 235079 14023 235107 14051
rect 235141 14023 235169 14051
rect 235203 14023 235231 14051
rect 235017 13961 235045 13989
rect 235079 13961 235107 13989
rect 235141 13961 235169 13989
rect 235203 13961 235231 13989
rect 246339 14147 246367 14175
rect 246401 14147 246429 14175
rect 246339 14085 246367 14113
rect 246401 14085 246429 14113
rect 246339 14023 246367 14051
rect 246401 14023 246429 14051
rect 246339 13961 246367 13989
rect 246401 13961 246429 13989
rect 238659 11147 238687 11175
rect 238721 11147 238749 11175
rect 238659 11085 238687 11113
rect 238721 11085 238749 11113
rect 238659 11023 238687 11051
rect 238721 11023 238749 11051
rect 238659 10961 238687 10989
rect 238721 10961 238749 10989
rect 248517 11147 248545 11175
rect 248579 11147 248607 11175
rect 248641 11147 248669 11175
rect 248703 11147 248731 11175
rect 248517 11085 248545 11113
rect 248579 11085 248607 11113
rect 248641 11085 248669 11113
rect 248703 11085 248731 11113
rect 248517 11023 248545 11051
rect 248579 11023 248607 11051
rect 248641 11023 248669 11051
rect 248703 11023 248731 11051
rect 248517 10961 248545 10989
rect 248579 10961 248607 10989
rect 248641 10961 248669 10989
rect 248703 10961 248731 10989
rect 235017 5147 235045 5175
rect 235079 5147 235107 5175
rect 235141 5147 235169 5175
rect 235203 5147 235231 5175
rect 235017 5085 235045 5113
rect 235079 5085 235107 5113
rect 235141 5085 235169 5113
rect 235203 5085 235231 5113
rect 235017 5023 235045 5051
rect 235079 5023 235107 5051
rect 235141 5023 235169 5051
rect 235203 5023 235231 5051
rect 235017 4961 235045 4989
rect 235079 4961 235107 4989
rect 235141 4961 235169 4989
rect 235203 4961 235231 4989
rect 246339 5147 246367 5175
rect 246401 5147 246429 5175
rect 246339 5085 246367 5113
rect 246401 5085 246429 5113
rect 246339 5023 246367 5051
rect 246401 5023 246429 5051
rect 246339 4961 246367 4989
rect 246401 4961 246429 4989
rect 235017 -588 235045 -560
rect 235079 -588 235107 -560
rect 235141 -588 235169 -560
rect 235203 -588 235231 -560
rect 235017 -650 235045 -622
rect 235079 -650 235107 -622
rect 235141 -650 235169 -622
rect 235203 -650 235231 -622
rect 235017 -712 235045 -684
rect 235079 -712 235107 -684
rect 235141 -712 235169 -684
rect 235203 -712 235231 -684
rect 235017 -774 235045 -746
rect 235079 -774 235107 -746
rect 235141 -774 235169 -746
rect 235203 -774 235231 -746
rect 248517 2147 248545 2175
rect 248579 2147 248607 2175
rect 248641 2147 248669 2175
rect 248703 2147 248731 2175
rect 248517 2085 248545 2113
rect 248579 2085 248607 2113
rect 248641 2085 248669 2113
rect 248703 2085 248731 2113
rect 248517 2023 248545 2051
rect 248579 2023 248607 2051
rect 248641 2023 248669 2051
rect 248703 2023 248731 2051
rect 248517 1961 248545 1989
rect 248579 1961 248607 1989
rect 248641 1961 248669 1989
rect 248703 1961 248731 1989
rect 248517 -108 248545 -80
rect 248579 -108 248607 -80
rect 248641 -108 248669 -80
rect 248703 -108 248731 -80
rect 248517 -170 248545 -142
rect 248579 -170 248607 -142
rect 248641 -170 248669 -142
rect 248703 -170 248731 -142
rect 248517 -232 248545 -204
rect 248579 -232 248607 -204
rect 248641 -232 248669 -204
rect 248703 -232 248731 -204
rect 248517 -294 248545 -266
rect 248579 -294 248607 -266
rect 248641 -294 248669 -266
rect 248703 -294 248731 -266
rect 250377 299058 250405 299086
rect 250439 299058 250467 299086
rect 250501 299058 250529 299086
rect 250563 299058 250591 299086
rect 250377 298996 250405 299024
rect 250439 298996 250467 299024
rect 250501 298996 250529 299024
rect 250563 298996 250591 299024
rect 250377 298934 250405 298962
rect 250439 298934 250467 298962
rect 250501 298934 250529 298962
rect 250563 298934 250591 298962
rect 250377 298872 250405 298900
rect 250439 298872 250467 298900
rect 250501 298872 250529 298900
rect 250563 298872 250591 298900
rect 250377 293147 250405 293175
rect 250439 293147 250467 293175
rect 250501 293147 250529 293175
rect 250563 293147 250591 293175
rect 250377 293085 250405 293113
rect 250439 293085 250467 293113
rect 250501 293085 250529 293113
rect 250563 293085 250591 293113
rect 250377 293023 250405 293051
rect 250439 293023 250467 293051
rect 250501 293023 250529 293051
rect 250563 293023 250591 293051
rect 250377 292961 250405 292989
rect 250439 292961 250467 292989
rect 250501 292961 250529 292989
rect 250563 292961 250591 292989
rect 250377 284147 250405 284175
rect 250439 284147 250467 284175
rect 250501 284147 250529 284175
rect 250563 284147 250591 284175
rect 250377 284085 250405 284113
rect 250439 284085 250467 284113
rect 250501 284085 250529 284113
rect 250563 284085 250591 284113
rect 250377 284023 250405 284051
rect 250439 284023 250467 284051
rect 250501 284023 250529 284051
rect 250563 284023 250591 284051
rect 250377 283961 250405 283989
rect 250439 283961 250467 283989
rect 250501 283961 250529 283989
rect 250563 283961 250591 283989
rect 250377 275147 250405 275175
rect 250439 275147 250467 275175
rect 250501 275147 250529 275175
rect 250563 275147 250591 275175
rect 250377 275085 250405 275113
rect 250439 275085 250467 275113
rect 250501 275085 250529 275113
rect 250563 275085 250591 275113
rect 250377 275023 250405 275051
rect 250439 275023 250467 275051
rect 250501 275023 250529 275051
rect 250563 275023 250591 275051
rect 250377 274961 250405 274989
rect 250439 274961 250467 274989
rect 250501 274961 250529 274989
rect 250563 274961 250591 274989
rect 250377 266147 250405 266175
rect 250439 266147 250467 266175
rect 250501 266147 250529 266175
rect 250563 266147 250591 266175
rect 250377 266085 250405 266113
rect 250439 266085 250467 266113
rect 250501 266085 250529 266113
rect 250563 266085 250591 266113
rect 250377 266023 250405 266051
rect 250439 266023 250467 266051
rect 250501 266023 250529 266051
rect 250563 266023 250591 266051
rect 250377 265961 250405 265989
rect 250439 265961 250467 265989
rect 250501 265961 250529 265989
rect 250563 265961 250591 265989
rect 250377 257147 250405 257175
rect 250439 257147 250467 257175
rect 250501 257147 250529 257175
rect 250563 257147 250591 257175
rect 250377 257085 250405 257113
rect 250439 257085 250467 257113
rect 250501 257085 250529 257113
rect 250563 257085 250591 257113
rect 250377 257023 250405 257051
rect 250439 257023 250467 257051
rect 250501 257023 250529 257051
rect 250563 257023 250591 257051
rect 250377 256961 250405 256989
rect 250439 256961 250467 256989
rect 250501 256961 250529 256989
rect 250563 256961 250591 256989
rect 250377 248147 250405 248175
rect 250439 248147 250467 248175
rect 250501 248147 250529 248175
rect 250563 248147 250591 248175
rect 250377 248085 250405 248113
rect 250439 248085 250467 248113
rect 250501 248085 250529 248113
rect 250563 248085 250591 248113
rect 250377 248023 250405 248051
rect 250439 248023 250467 248051
rect 250501 248023 250529 248051
rect 250563 248023 250591 248051
rect 250377 247961 250405 247989
rect 250439 247961 250467 247989
rect 250501 247961 250529 247989
rect 250563 247961 250591 247989
rect 250377 239147 250405 239175
rect 250439 239147 250467 239175
rect 250501 239147 250529 239175
rect 250563 239147 250591 239175
rect 250377 239085 250405 239113
rect 250439 239085 250467 239113
rect 250501 239085 250529 239113
rect 250563 239085 250591 239113
rect 250377 239023 250405 239051
rect 250439 239023 250467 239051
rect 250501 239023 250529 239051
rect 250563 239023 250591 239051
rect 250377 238961 250405 238989
rect 250439 238961 250467 238989
rect 250501 238961 250529 238989
rect 250563 238961 250591 238989
rect 250377 230147 250405 230175
rect 250439 230147 250467 230175
rect 250501 230147 250529 230175
rect 250563 230147 250591 230175
rect 250377 230085 250405 230113
rect 250439 230085 250467 230113
rect 250501 230085 250529 230113
rect 250563 230085 250591 230113
rect 250377 230023 250405 230051
rect 250439 230023 250467 230051
rect 250501 230023 250529 230051
rect 250563 230023 250591 230051
rect 250377 229961 250405 229989
rect 250439 229961 250467 229989
rect 250501 229961 250529 229989
rect 250563 229961 250591 229989
rect 250377 221147 250405 221175
rect 250439 221147 250467 221175
rect 250501 221147 250529 221175
rect 250563 221147 250591 221175
rect 250377 221085 250405 221113
rect 250439 221085 250467 221113
rect 250501 221085 250529 221113
rect 250563 221085 250591 221113
rect 250377 221023 250405 221051
rect 250439 221023 250467 221051
rect 250501 221023 250529 221051
rect 250563 221023 250591 221051
rect 250377 220961 250405 220989
rect 250439 220961 250467 220989
rect 250501 220961 250529 220989
rect 250563 220961 250591 220989
rect 250377 212147 250405 212175
rect 250439 212147 250467 212175
rect 250501 212147 250529 212175
rect 250563 212147 250591 212175
rect 250377 212085 250405 212113
rect 250439 212085 250467 212113
rect 250501 212085 250529 212113
rect 250563 212085 250591 212113
rect 250377 212023 250405 212051
rect 250439 212023 250467 212051
rect 250501 212023 250529 212051
rect 250563 212023 250591 212051
rect 250377 211961 250405 211989
rect 250439 211961 250467 211989
rect 250501 211961 250529 211989
rect 250563 211961 250591 211989
rect 250377 203147 250405 203175
rect 250439 203147 250467 203175
rect 250501 203147 250529 203175
rect 250563 203147 250591 203175
rect 250377 203085 250405 203113
rect 250439 203085 250467 203113
rect 250501 203085 250529 203113
rect 250563 203085 250591 203113
rect 250377 203023 250405 203051
rect 250439 203023 250467 203051
rect 250501 203023 250529 203051
rect 250563 203023 250591 203051
rect 250377 202961 250405 202989
rect 250439 202961 250467 202989
rect 250501 202961 250529 202989
rect 250563 202961 250591 202989
rect 250377 194147 250405 194175
rect 250439 194147 250467 194175
rect 250501 194147 250529 194175
rect 250563 194147 250591 194175
rect 250377 194085 250405 194113
rect 250439 194085 250467 194113
rect 250501 194085 250529 194113
rect 250563 194085 250591 194113
rect 250377 194023 250405 194051
rect 250439 194023 250467 194051
rect 250501 194023 250529 194051
rect 250563 194023 250591 194051
rect 250377 193961 250405 193989
rect 250439 193961 250467 193989
rect 250501 193961 250529 193989
rect 250563 193961 250591 193989
rect 250377 185147 250405 185175
rect 250439 185147 250467 185175
rect 250501 185147 250529 185175
rect 250563 185147 250591 185175
rect 250377 185085 250405 185113
rect 250439 185085 250467 185113
rect 250501 185085 250529 185113
rect 250563 185085 250591 185113
rect 250377 185023 250405 185051
rect 250439 185023 250467 185051
rect 250501 185023 250529 185051
rect 250563 185023 250591 185051
rect 250377 184961 250405 184989
rect 250439 184961 250467 184989
rect 250501 184961 250529 184989
rect 250563 184961 250591 184989
rect 250377 176147 250405 176175
rect 250439 176147 250467 176175
rect 250501 176147 250529 176175
rect 250563 176147 250591 176175
rect 250377 176085 250405 176113
rect 250439 176085 250467 176113
rect 250501 176085 250529 176113
rect 250563 176085 250591 176113
rect 250377 176023 250405 176051
rect 250439 176023 250467 176051
rect 250501 176023 250529 176051
rect 250563 176023 250591 176051
rect 250377 175961 250405 175989
rect 250439 175961 250467 175989
rect 250501 175961 250529 175989
rect 250563 175961 250591 175989
rect 263877 298578 263905 298606
rect 263939 298578 263967 298606
rect 264001 298578 264029 298606
rect 264063 298578 264091 298606
rect 263877 298516 263905 298544
rect 263939 298516 263967 298544
rect 264001 298516 264029 298544
rect 264063 298516 264091 298544
rect 263877 298454 263905 298482
rect 263939 298454 263967 298482
rect 264001 298454 264029 298482
rect 264063 298454 264091 298482
rect 263877 298392 263905 298420
rect 263939 298392 263967 298420
rect 264001 298392 264029 298420
rect 264063 298392 264091 298420
rect 263877 290147 263905 290175
rect 263939 290147 263967 290175
rect 264001 290147 264029 290175
rect 264063 290147 264091 290175
rect 263877 290085 263905 290113
rect 263939 290085 263967 290113
rect 264001 290085 264029 290113
rect 264063 290085 264091 290113
rect 263877 290023 263905 290051
rect 263939 290023 263967 290051
rect 264001 290023 264029 290051
rect 264063 290023 264091 290051
rect 263877 289961 263905 289989
rect 263939 289961 263967 289989
rect 264001 289961 264029 289989
rect 264063 289961 264091 289989
rect 263877 281147 263905 281175
rect 263939 281147 263967 281175
rect 264001 281147 264029 281175
rect 264063 281147 264091 281175
rect 263877 281085 263905 281113
rect 263939 281085 263967 281113
rect 264001 281085 264029 281113
rect 264063 281085 264091 281113
rect 263877 281023 263905 281051
rect 263939 281023 263967 281051
rect 264001 281023 264029 281051
rect 264063 281023 264091 281051
rect 263877 280961 263905 280989
rect 263939 280961 263967 280989
rect 264001 280961 264029 280989
rect 264063 280961 264091 280989
rect 263877 272147 263905 272175
rect 263939 272147 263967 272175
rect 264001 272147 264029 272175
rect 264063 272147 264091 272175
rect 263877 272085 263905 272113
rect 263939 272085 263967 272113
rect 264001 272085 264029 272113
rect 264063 272085 264091 272113
rect 263877 272023 263905 272051
rect 263939 272023 263967 272051
rect 264001 272023 264029 272051
rect 264063 272023 264091 272051
rect 263877 271961 263905 271989
rect 263939 271961 263967 271989
rect 264001 271961 264029 271989
rect 264063 271961 264091 271989
rect 263877 263147 263905 263175
rect 263939 263147 263967 263175
rect 264001 263147 264029 263175
rect 264063 263147 264091 263175
rect 263877 263085 263905 263113
rect 263939 263085 263967 263113
rect 264001 263085 264029 263113
rect 264063 263085 264091 263113
rect 263877 263023 263905 263051
rect 263939 263023 263967 263051
rect 264001 263023 264029 263051
rect 264063 263023 264091 263051
rect 263877 262961 263905 262989
rect 263939 262961 263967 262989
rect 264001 262961 264029 262989
rect 264063 262961 264091 262989
rect 263877 254147 263905 254175
rect 263939 254147 263967 254175
rect 264001 254147 264029 254175
rect 264063 254147 264091 254175
rect 263877 254085 263905 254113
rect 263939 254085 263967 254113
rect 264001 254085 264029 254113
rect 264063 254085 264091 254113
rect 263877 254023 263905 254051
rect 263939 254023 263967 254051
rect 264001 254023 264029 254051
rect 264063 254023 264091 254051
rect 263877 253961 263905 253989
rect 263939 253961 263967 253989
rect 264001 253961 264029 253989
rect 264063 253961 264091 253989
rect 263877 245147 263905 245175
rect 263939 245147 263967 245175
rect 264001 245147 264029 245175
rect 264063 245147 264091 245175
rect 263877 245085 263905 245113
rect 263939 245085 263967 245113
rect 264001 245085 264029 245113
rect 264063 245085 264091 245113
rect 263877 245023 263905 245051
rect 263939 245023 263967 245051
rect 264001 245023 264029 245051
rect 264063 245023 264091 245051
rect 263877 244961 263905 244989
rect 263939 244961 263967 244989
rect 264001 244961 264029 244989
rect 264063 244961 264091 244989
rect 263877 236147 263905 236175
rect 263939 236147 263967 236175
rect 264001 236147 264029 236175
rect 264063 236147 264091 236175
rect 263877 236085 263905 236113
rect 263939 236085 263967 236113
rect 264001 236085 264029 236113
rect 264063 236085 264091 236113
rect 263877 236023 263905 236051
rect 263939 236023 263967 236051
rect 264001 236023 264029 236051
rect 264063 236023 264091 236051
rect 263877 235961 263905 235989
rect 263939 235961 263967 235989
rect 264001 235961 264029 235989
rect 264063 235961 264091 235989
rect 263877 227147 263905 227175
rect 263939 227147 263967 227175
rect 264001 227147 264029 227175
rect 264063 227147 264091 227175
rect 263877 227085 263905 227113
rect 263939 227085 263967 227113
rect 264001 227085 264029 227113
rect 264063 227085 264091 227113
rect 263877 227023 263905 227051
rect 263939 227023 263967 227051
rect 264001 227023 264029 227051
rect 264063 227023 264091 227051
rect 263877 226961 263905 226989
rect 263939 226961 263967 226989
rect 264001 226961 264029 226989
rect 264063 226961 264091 226989
rect 263877 218147 263905 218175
rect 263939 218147 263967 218175
rect 264001 218147 264029 218175
rect 264063 218147 264091 218175
rect 263877 218085 263905 218113
rect 263939 218085 263967 218113
rect 264001 218085 264029 218113
rect 264063 218085 264091 218113
rect 263877 218023 263905 218051
rect 263939 218023 263967 218051
rect 264001 218023 264029 218051
rect 264063 218023 264091 218051
rect 263877 217961 263905 217989
rect 263939 217961 263967 217989
rect 264001 217961 264029 217989
rect 264063 217961 264091 217989
rect 263877 209147 263905 209175
rect 263939 209147 263967 209175
rect 264001 209147 264029 209175
rect 264063 209147 264091 209175
rect 263877 209085 263905 209113
rect 263939 209085 263967 209113
rect 264001 209085 264029 209113
rect 264063 209085 264091 209113
rect 263877 209023 263905 209051
rect 263939 209023 263967 209051
rect 264001 209023 264029 209051
rect 264063 209023 264091 209051
rect 263877 208961 263905 208989
rect 263939 208961 263967 208989
rect 264001 208961 264029 208989
rect 264063 208961 264091 208989
rect 263877 200147 263905 200175
rect 263939 200147 263967 200175
rect 264001 200147 264029 200175
rect 264063 200147 264091 200175
rect 263877 200085 263905 200113
rect 263939 200085 263967 200113
rect 264001 200085 264029 200113
rect 264063 200085 264091 200113
rect 263877 200023 263905 200051
rect 263939 200023 263967 200051
rect 264001 200023 264029 200051
rect 264063 200023 264091 200051
rect 263877 199961 263905 199989
rect 263939 199961 263967 199989
rect 264001 199961 264029 199989
rect 264063 199961 264091 199989
rect 263877 191147 263905 191175
rect 263939 191147 263967 191175
rect 264001 191147 264029 191175
rect 264063 191147 264091 191175
rect 263877 191085 263905 191113
rect 263939 191085 263967 191113
rect 264001 191085 264029 191113
rect 264063 191085 264091 191113
rect 263877 191023 263905 191051
rect 263939 191023 263967 191051
rect 264001 191023 264029 191051
rect 264063 191023 264091 191051
rect 263877 190961 263905 190989
rect 263939 190961 263967 190989
rect 264001 190961 264029 190989
rect 264063 190961 264091 190989
rect 263877 182147 263905 182175
rect 263939 182147 263967 182175
rect 264001 182147 264029 182175
rect 264063 182147 264091 182175
rect 263877 182085 263905 182113
rect 263939 182085 263967 182113
rect 264001 182085 264029 182113
rect 264063 182085 264091 182113
rect 263877 182023 263905 182051
rect 263939 182023 263967 182051
rect 264001 182023 264029 182051
rect 264063 182023 264091 182051
rect 263877 181961 263905 181989
rect 263939 181961 263967 181989
rect 264001 181961 264029 181989
rect 264063 181961 264091 181989
rect 254019 173147 254047 173175
rect 254081 173147 254109 173175
rect 254019 173085 254047 173113
rect 254081 173085 254109 173113
rect 254019 173023 254047 173051
rect 254081 173023 254109 173051
rect 254019 172961 254047 172989
rect 254081 172961 254109 172989
rect 263877 173147 263905 173175
rect 263939 173147 263967 173175
rect 264001 173147 264029 173175
rect 264063 173147 264091 173175
rect 263877 173085 263905 173113
rect 263939 173085 263967 173113
rect 264001 173085 264029 173113
rect 264063 173085 264091 173113
rect 263877 173023 263905 173051
rect 263939 173023 263967 173051
rect 264001 173023 264029 173051
rect 264063 173023 264091 173051
rect 263877 172961 263905 172989
rect 263939 172961 263967 172989
rect 264001 172961 264029 172989
rect 264063 172961 264091 172989
rect 250377 167147 250405 167175
rect 250439 167147 250467 167175
rect 250501 167147 250529 167175
rect 250563 167147 250591 167175
rect 250377 167085 250405 167113
rect 250439 167085 250467 167113
rect 250501 167085 250529 167113
rect 250563 167085 250591 167113
rect 250377 167023 250405 167051
rect 250439 167023 250467 167051
rect 250501 167023 250529 167051
rect 250563 167023 250591 167051
rect 250377 166961 250405 166989
rect 250439 166961 250467 166989
rect 250501 166961 250529 166989
rect 250563 166961 250591 166989
rect 261699 167147 261727 167175
rect 261761 167147 261789 167175
rect 261699 167085 261727 167113
rect 261761 167085 261789 167113
rect 261699 167023 261727 167051
rect 261761 167023 261789 167051
rect 261699 166961 261727 166989
rect 261761 166961 261789 166989
rect 254019 164147 254047 164175
rect 254081 164147 254109 164175
rect 254019 164085 254047 164113
rect 254081 164085 254109 164113
rect 254019 164023 254047 164051
rect 254081 164023 254109 164051
rect 254019 163961 254047 163989
rect 254081 163961 254109 163989
rect 263877 164147 263905 164175
rect 263939 164147 263967 164175
rect 264001 164147 264029 164175
rect 264063 164147 264091 164175
rect 263877 164085 263905 164113
rect 263939 164085 263967 164113
rect 264001 164085 264029 164113
rect 264063 164085 264091 164113
rect 263877 164023 263905 164051
rect 263939 164023 263967 164051
rect 264001 164023 264029 164051
rect 264063 164023 264091 164051
rect 263877 163961 263905 163989
rect 263939 163961 263967 163989
rect 264001 163961 264029 163989
rect 264063 163961 264091 163989
rect 250377 158147 250405 158175
rect 250439 158147 250467 158175
rect 250501 158147 250529 158175
rect 250563 158147 250591 158175
rect 250377 158085 250405 158113
rect 250439 158085 250467 158113
rect 250501 158085 250529 158113
rect 250563 158085 250591 158113
rect 250377 158023 250405 158051
rect 250439 158023 250467 158051
rect 250501 158023 250529 158051
rect 250563 158023 250591 158051
rect 250377 157961 250405 157989
rect 250439 157961 250467 157989
rect 250501 157961 250529 157989
rect 250563 157961 250591 157989
rect 261699 158147 261727 158175
rect 261761 158147 261789 158175
rect 261699 158085 261727 158113
rect 261761 158085 261789 158113
rect 261699 158023 261727 158051
rect 261761 158023 261789 158051
rect 261699 157961 261727 157989
rect 261761 157961 261789 157989
rect 254019 155147 254047 155175
rect 254081 155147 254109 155175
rect 254019 155085 254047 155113
rect 254081 155085 254109 155113
rect 254019 155023 254047 155051
rect 254081 155023 254109 155051
rect 254019 154961 254047 154989
rect 254081 154961 254109 154989
rect 263877 155147 263905 155175
rect 263939 155147 263967 155175
rect 264001 155147 264029 155175
rect 264063 155147 264091 155175
rect 263877 155085 263905 155113
rect 263939 155085 263967 155113
rect 264001 155085 264029 155113
rect 264063 155085 264091 155113
rect 263877 155023 263905 155051
rect 263939 155023 263967 155051
rect 264001 155023 264029 155051
rect 264063 155023 264091 155051
rect 263877 154961 263905 154989
rect 263939 154961 263967 154989
rect 264001 154961 264029 154989
rect 264063 154961 264091 154989
rect 250377 149147 250405 149175
rect 250439 149147 250467 149175
rect 250501 149147 250529 149175
rect 250563 149147 250591 149175
rect 250377 149085 250405 149113
rect 250439 149085 250467 149113
rect 250501 149085 250529 149113
rect 250563 149085 250591 149113
rect 250377 149023 250405 149051
rect 250439 149023 250467 149051
rect 250501 149023 250529 149051
rect 250563 149023 250591 149051
rect 250377 148961 250405 148989
rect 250439 148961 250467 148989
rect 250501 148961 250529 148989
rect 250563 148961 250591 148989
rect 261699 149147 261727 149175
rect 261761 149147 261789 149175
rect 261699 149085 261727 149113
rect 261761 149085 261789 149113
rect 261699 149023 261727 149051
rect 261761 149023 261789 149051
rect 261699 148961 261727 148989
rect 261761 148961 261789 148989
rect 254019 146147 254047 146175
rect 254081 146147 254109 146175
rect 254019 146085 254047 146113
rect 254081 146085 254109 146113
rect 254019 146023 254047 146051
rect 254081 146023 254109 146051
rect 254019 145961 254047 145989
rect 254081 145961 254109 145989
rect 263877 146147 263905 146175
rect 263939 146147 263967 146175
rect 264001 146147 264029 146175
rect 264063 146147 264091 146175
rect 263877 146085 263905 146113
rect 263939 146085 263967 146113
rect 264001 146085 264029 146113
rect 264063 146085 264091 146113
rect 263877 146023 263905 146051
rect 263939 146023 263967 146051
rect 264001 146023 264029 146051
rect 264063 146023 264091 146051
rect 263877 145961 263905 145989
rect 263939 145961 263967 145989
rect 264001 145961 264029 145989
rect 264063 145961 264091 145989
rect 250377 140147 250405 140175
rect 250439 140147 250467 140175
rect 250501 140147 250529 140175
rect 250563 140147 250591 140175
rect 250377 140085 250405 140113
rect 250439 140085 250467 140113
rect 250501 140085 250529 140113
rect 250563 140085 250591 140113
rect 250377 140023 250405 140051
rect 250439 140023 250467 140051
rect 250501 140023 250529 140051
rect 250563 140023 250591 140051
rect 250377 139961 250405 139989
rect 250439 139961 250467 139989
rect 250501 139961 250529 139989
rect 250563 139961 250591 139989
rect 261699 140147 261727 140175
rect 261761 140147 261789 140175
rect 261699 140085 261727 140113
rect 261761 140085 261789 140113
rect 261699 140023 261727 140051
rect 261761 140023 261789 140051
rect 261699 139961 261727 139989
rect 261761 139961 261789 139989
rect 254019 137147 254047 137175
rect 254081 137147 254109 137175
rect 254019 137085 254047 137113
rect 254081 137085 254109 137113
rect 254019 137023 254047 137051
rect 254081 137023 254109 137051
rect 254019 136961 254047 136989
rect 254081 136961 254109 136989
rect 263877 137147 263905 137175
rect 263939 137147 263967 137175
rect 264001 137147 264029 137175
rect 264063 137147 264091 137175
rect 263877 137085 263905 137113
rect 263939 137085 263967 137113
rect 264001 137085 264029 137113
rect 264063 137085 264091 137113
rect 263877 137023 263905 137051
rect 263939 137023 263967 137051
rect 264001 137023 264029 137051
rect 264063 137023 264091 137051
rect 263877 136961 263905 136989
rect 263939 136961 263967 136989
rect 264001 136961 264029 136989
rect 264063 136961 264091 136989
rect 250377 131147 250405 131175
rect 250439 131147 250467 131175
rect 250501 131147 250529 131175
rect 250563 131147 250591 131175
rect 250377 131085 250405 131113
rect 250439 131085 250467 131113
rect 250501 131085 250529 131113
rect 250563 131085 250591 131113
rect 250377 131023 250405 131051
rect 250439 131023 250467 131051
rect 250501 131023 250529 131051
rect 250563 131023 250591 131051
rect 250377 130961 250405 130989
rect 250439 130961 250467 130989
rect 250501 130961 250529 130989
rect 250563 130961 250591 130989
rect 261699 131147 261727 131175
rect 261761 131147 261789 131175
rect 261699 131085 261727 131113
rect 261761 131085 261789 131113
rect 261699 131023 261727 131051
rect 261761 131023 261789 131051
rect 261699 130961 261727 130989
rect 261761 130961 261789 130989
rect 254019 128147 254047 128175
rect 254081 128147 254109 128175
rect 254019 128085 254047 128113
rect 254081 128085 254109 128113
rect 254019 128023 254047 128051
rect 254081 128023 254109 128051
rect 254019 127961 254047 127989
rect 254081 127961 254109 127989
rect 263877 128147 263905 128175
rect 263939 128147 263967 128175
rect 264001 128147 264029 128175
rect 264063 128147 264091 128175
rect 263877 128085 263905 128113
rect 263939 128085 263967 128113
rect 264001 128085 264029 128113
rect 264063 128085 264091 128113
rect 263877 128023 263905 128051
rect 263939 128023 263967 128051
rect 264001 128023 264029 128051
rect 264063 128023 264091 128051
rect 263877 127961 263905 127989
rect 263939 127961 263967 127989
rect 264001 127961 264029 127989
rect 264063 127961 264091 127989
rect 250377 122147 250405 122175
rect 250439 122147 250467 122175
rect 250501 122147 250529 122175
rect 250563 122147 250591 122175
rect 250377 122085 250405 122113
rect 250439 122085 250467 122113
rect 250501 122085 250529 122113
rect 250563 122085 250591 122113
rect 250377 122023 250405 122051
rect 250439 122023 250467 122051
rect 250501 122023 250529 122051
rect 250563 122023 250591 122051
rect 250377 121961 250405 121989
rect 250439 121961 250467 121989
rect 250501 121961 250529 121989
rect 250563 121961 250591 121989
rect 261699 122147 261727 122175
rect 261761 122147 261789 122175
rect 261699 122085 261727 122113
rect 261761 122085 261789 122113
rect 261699 122023 261727 122051
rect 261761 122023 261789 122051
rect 261699 121961 261727 121989
rect 261761 121961 261789 121989
rect 254019 119147 254047 119175
rect 254081 119147 254109 119175
rect 254019 119085 254047 119113
rect 254081 119085 254109 119113
rect 254019 119023 254047 119051
rect 254081 119023 254109 119051
rect 254019 118961 254047 118989
rect 254081 118961 254109 118989
rect 263877 119147 263905 119175
rect 263939 119147 263967 119175
rect 264001 119147 264029 119175
rect 264063 119147 264091 119175
rect 263877 119085 263905 119113
rect 263939 119085 263967 119113
rect 264001 119085 264029 119113
rect 264063 119085 264091 119113
rect 263877 119023 263905 119051
rect 263939 119023 263967 119051
rect 264001 119023 264029 119051
rect 264063 119023 264091 119051
rect 263877 118961 263905 118989
rect 263939 118961 263967 118989
rect 264001 118961 264029 118989
rect 264063 118961 264091 118989
rect 250377 113147 250405 113175
rect 250439 113147 250467 113175
rect 250501 113147 250529 113175
rect 250563 113147 250591 113175
rect 250377 113085 250405 113113
rect 250439 113085 250467 113113
rect 250501 113085 250529 113113
rect 250563 113085 250591 113113
rect 250377 113023 250405 113051
rect 250439 113023 250467 113051
rect 250501 113023 250529 113051
rect 250563 113023 250591 113051
rect 250377 112961 250405 112989
rect 250439 112961 250467 112989
rect 250501 112961 250529 112989
rect 250563 112961 250591 112989
rect 261699 113147 261727 113175
rect 261761 113147 261789 113175
rect 261699 113085 261727 113113
rect 261761 113085 261789 113113
rect 261699 113023 261727 113051
rect 261761 113023 261789 113051
rect 261699 112961 261727 112989
rect 261761 112961 261789 112989
rect 254019 110147 254047 110175
rect 254081 110147 254109 110175
rect 254019 110085 254047 110113
rect 254081 110085 254109 110113
rect 254019 110023 254047 110051
rect 254081 110023 254109 110051
rect 254019 109961 254047 109989
rect 254081 109961 254109 109989
rect 263877 110147 263905 110175
rect 263939 110147 263967 110175
rect 264001 110147 264029 110175
rect 264063 110147 264091 110175
rect 263877 110085 263905 110113
rect 263939 110085 263967 110113
rect 264001 110085 264029 110113
rect 264063 110085 264091 110113
rect 263877 110023 263905 110051
rect 263939 110023 263967 110051
rect 264001 110023 264029 110051
rect 264063 110023 264091 110051
rect 263877 109961 263905 109989
rect 263939 109961 263967 109989
rect 264001 109961 264029 109989
rect 264063 109961 264091 109989
rect 250377 104147 250405 104175
rect 250439 104147 250467 104175
rect 250501 104147 250529 104175
rect 250563 104147 250591 104175
rect 250377 104085 250405 104113
rect 250439 104085 250467 104113
rect 250501 104085 250529 104113
rect 250563 104085 250591 104113
rect 250377 104023 250405 104051
rect 250439 104023 250467 104051
rect 250501 104023 250529 104051
rect 250563 104023 250591 104051
rect 250377 103961 250405 103989
rect 250439 103961 250467 103989
rect 250501 103961 250529 103989
rect 250563 103961 250591 103989
rect 261699 104147 261727 104175
rect 261761 104147 261789 104175
rect 261699 104085 261727 104113
rect 261761 104085 261789 104113
rect 261699 104023 261727 104051
rect 261761 104023 261789 104051
rect 261699 103961 261727 103989
rect 261761 103961 261789 103989
rect 254019 101147 254047 101175
rect 254081 101147 254109 101175
rect 254019 101085 254047 101113
rect 254081 101085 254109 101113
rect 254019 101023 254047 101051
rect 254081 101023 254109 101051
rect 254019 100961 254047 100989
rect 254081 100961 254109 100989
rect 263877 101147 263905 101175
rect 263939 101147 263967 101175
rect 264001 101147 264029 101175
rect 264063 101147 264091 101175
rect 263877 101085 263905 101113
rect 263939 101085 263967 101113
rect 264001 101085 264029 101113
rect 264063 101085 264091 101113
rect 263877 101023 263905 101051
rect 263939 101023 263967 101051
rect 264001 101023 264029 101051
rect 264063 101023 264091 101051
rect 263877 100961 263905 100989
rect 263939 100961 263967 100989
rect 264001 100961 264029 100989
rect 264063 100961 264091 100989
rect 250377 95147 250405 95175
rect 250439 95147 250467 95175
rect 250501 95147 250529 95175
rect 250563 95147 250591 95175
rect 250377 95085 250405 95113
rect 250439 95085 250467 95113
rect 250501 95085 250529 95113
rect 250563 95085 250591 95113
rect 250377 95023 250405 95051
rect 250439 95023 250467 95051
rect 250501 95023 250529 95051
rect 250563 95023 250591 95051
rect 250377 94961 250405 94989
rect 250439 94961 250467 94989
rect 250501 94961 250529 94989
rect 250563 94961 250591 94989
rect 261699 95147 261727 95175
rect 261761 95147 261789 95175
rect 261699 95085 261727 95113
rect 261761 95085 261789 95113
rect 261699 95023 261727 95051
rect 261761 95023 261789 95051
rect 261699 94961 261727 94989
rect 261761 94961 261789 94989
rect 254019 92147 254047 92175
rect 254081 92147 254109 92175
rect 254019 92085 254047 92113
rect 254081 92085 254109 92113
rect 254019 92023 254047 92051
rect 254081 92023 254109 92051
rect 254019 91961 254047 91989
rect 254081 91961 254109 91989
rect 263877 92147 263905 92175
rect 263939 92147 263967 92175
rect 264001 92147 264029 92175
rect 264063 92147 264091 92175
rect 263877 92085 263905 92113
rect 263939 92085 263967 92113
rect 264001 92085 264029 92113
rect 264063 92085 264091 92113
rect 263877 92023 263905 92051
rect 263939 92023 263967 92051
rect 264001 92023 264029 92051
rect 264063 92023 264091 92051
rect 263877 91961 263905 91989
rect 263939 91961 263967 91989
rect 264001 91961 264029 91989
rect 264063 91961 264091 91989
rect 250377 86147 250405 86175
rect 250439 86147 250467 86175
rect 250501 86147 250529 86175
rect 250563 86147 250591 86175
rect 250377 86085 250405 86113
rect 250439 86085 250467 86113
rect 250501 86085 250529 86113
rect 250563 86085 250591 86113
rect 250377 86023 250405 86051
rect 250439 86023 250467 86051
rect 250501 86023 250529 86051
rect 250563 86023 250591 86051
rect 250377 85961 250405 85989
rect 250439 85961 250467 85989
rect 250501 85961 250529 85989
rect 250563 85961 250591 85989
rect 261699 86147 261727 86175
rect 261761 86147 261789 86175
rect 261699 86085 261727 86113
rect 261761 86085 261789 86113
rect 261699 86023 261727 86051
rect 261761 86023 261789 86051
rect 261699 85961 261727 85989
rect 261761 85961 261789 85989
rect 254019 83147 254047 83175
rect 254081 83147 254109 83175
rect 254019 83085 254047 83113
rect 254081 83085 254109 83113
rect 254019 83023 254047 83051
rect 254081 83023 254109 83051
rect 254019 82961 254047 82989
rect 254081 82961 254109 82989
rect 263877 83147 263905 83175
rect 263939 83147 263967 83175
rect 264001 83147 264029 83175
rect 264063 83147 264091 83175
rect 263877 83085 263905 83113
rect 263939 83085 263967 83113
rect 264001 83085 264029 83113
rect 264063 83085 264091 83113
rect 263877 83023 263905 83051
rect 263939 83023 263967 83051
rect 264001 83023 264029 83051
rect 264063 83023 264091 83051
rect 263877 82961 263905 82989
rect 263939 82961 263967 82989
rect 264001 82961 264029 82989
rect 264063 82961 264091 82989
rect 250377 77147 250405 77175
rect 250439 77147 250467 77175
rect 250501 77147 250529 77175
rect 250563 77147 250591 77175
rect 250377 77085 250405 77113
rect 250439 77085 250467 77113
rect 250501 77085 250529 77113
rect 250563 77085 250591 77113
rect 250377 77023 250405 77051
rect 250439 77023 250467 77051
rect 250501 77023 250529 77051
rect 250563 77023 250591 77051
rect 250377 76961 250405 76989
rect 250439 76961 250467 76989
rect 250501 76961 250529 76989
rect 250563 76961 250591 76989
rect 261699 77147 261727 77175
rect 261761 77147 261789 77175
rect 261699 77085 261727 77113
rect 261761 77085 261789 77113
rect 261699 77023 261727 77051
rect 261761 77023 261789 77051
rect 261699 76961 261727 76989
rect 261761 76961 261789 76989
rect 254019 74147 254047 74175
rect 254081 74147 254109 74175
rect 254019 74085 254047 74113
rect 254081 74085 254109 74113
rect 254019 74023 254047 74051
rect 254081 74023 254109 74051
rect 254019 73961 254047 73989
rect 254081 73961 254109 73989
rect 263877 74147 263905 74175
rect 263939 74147 263967 74175
rect 264001 74147 264029 74175
rect 264063 74147 264091 74175
rect 263877 74085 263905 74113
rect 263939 74085 263967 74113
rect 264001 74085 264029 74113
rect 264063 74085 264091 74113
rect 263877 74023 263905 74051
rect 263939 74023 263967 74051
rect 264001 74023 264029 74051
rect 264063 74023 264091 74051
rect 263877 73961 263905 73989
rect 263939 73961 263967 73989
rect 264001 73961 264029 73989
rect 264063 73961 264091 73989
rect 250377 68147 250405 68175
rect 250439 68147 250467 68175
rect 250501 68147 250529 68175
rect 250563 68147 250591 68175
rect 250377 68085 250405 68113
rect 250439 68085 250467 68113
rect 250501 68085 250529 68113
rect 250563 68085 250591 68113
rect 250377 68023 250405 68051
rect 250439 68023 250467 68051
rect 250501 68023 250529 68051
rect 250563 68023 250591 68051
rect 250377 67961 250405 67989
rect 250439 67961 250467 67989
rect 250501 67961 250529 67989
rect 250563 67961 250591 67989
rect 261699 68147 261727 68175
rect 261761 68147 261789 68175
rect 261699 68085 261727 68113
rect 261761 68085 261789 68113
rect 261699 68023 261727 68051
rect 261761 68023 261789 68051
rect 261699 67961 261727 67989
rect 261761 67961 261789 67989
rect 254019 65147 254047 65175
rect 254081 65147 254109 65175
rect 254019 65085 254047 65113
rect 254081 65085 254109 65113
rect 254019 65023 254047 65051
rect 254081 65023 254109 65051
rect 254019 64961 254047 64989
rect 254081 64961 254109 64989
rect 263877 65147 263905 65175
rect 263939 65147 263967 65175
rect 264001 65147 264029 65175
rect 264063 65147 264091 65175
rect 263877 65085 263905 65113
rect 263939 65085 263967 65113
rect 264001 65085 264029 65113
rect 264063 65085 264091 65113
rect 263877 65023 263905 65051
rect 263939 65023 263967 65051
rect 264001 65023 264029 65051
rect 264063 65023 264091 65051
rect 263877 64961 263905 64989
rect 263939 64961 263967 64989
rect 264001 64961 264029 64989
rect 264063 64961 264091 64989
rect 250377 59147 250405 59175
rect 250439 59147 250467 59175
rect 250501 59147 250529 59175
rect 250563 59147 250591 59175
rect 250377 59085 250405 59113
rect 250439 59085 250467 59113
rect 250501 59085 250529 59113
rect 250563 59085 250591 59113
rect 250377 59023 250405 59051
rect 250439 59023 250467 59051
rect 250501 59023 250529 59051
rect 250563 59023 250591 59051
rect 250377 58961 250405 58989
rect 250439 58961 250467 58989
rect 250501 58961 250529 58989
rect 250563 58961 250591 58989
rect 261699 59147 261727 59175
rect 261761 59147 261789 59175
rect 261699 59085 261727 59113
rect 261761 59085 261789 59113
rect 261699 59023 261727 59051
rect 261761 59023 261789 59051
rect 261699 58961 261727 58989
rect 261761 58961 261789 58989
rect 254019 56147 254047 56175
rect 254081 56147 254109 56175
rect 254019 56085 254047 56113
rect 254081 56085 254109 56113
rect 254019 56023 254047 56051
rect 254081 56023 254109 56051
rect 254019 55961 254047 55989
rect 254081 55961 254109 55989
rect 263877 56147 263905 56175
rect 263939 56147 263967 56175
rect 264001 56147 264029 56175
rect 264063 56147 264091 56175
rect 263877 56085 263905 56113
rect 263939 56085 263967 56113
rect 264001 56085 264029 56113
rect 264063 56085 264091 56113
rect 263877 56023 263905 56051
rect 263939 56023 263967 56051
rect 264001 56023 264029 56051
rect 264063 56023 264091 56051
rect 263877 55961 263905 55989
rect 263939 55961 263967 55989
rect 264001 55961 264029 55989
rect 264063 55961 264091 55989
rect 250377 50147 250405 50175
rect 250439 50147 250467 50175
rect 250501 50147 250529 50175
rect 250563 50147 250591 50175
rect 250377 50085 250405 50113
rect 250439 50085 250467 50113
rect 250501 50085 250529 50113
rect 250563 50085 250591 50113
rect 250377 50023 250405 50051
rect 250439 50023 250467 50051
rect 250501 50023 250529 50051
rect 250563 50023 250591 50051
rect 250377 49961 250405 49989
rect 250439 49961 250467 49989
rect 250501 49961 250529 49989
rect 250563 49961 250591 49989
rect 261699 50147 261727 50175
rect 261761 50147 261789 50175
rect 261699 50085 261727 50113
rect 261761 50085 261789 50113
rect 261699 50023 261727 50051
rect 261761 50023 261789 50051
rect 261699 49961 261727 49989
rect 261761 49961 261789 49989
rect 254019 47147 254047 47175
rect 254081 47147 254109 47175
rect 254019 47085 254047 47113
rect 254081 47085 254109 47113
rect 254019 47023 254047 47051
rect 254081 47023 254109 47051
rect 254019 46961 254047 46989
rect 254081 46961 254109 46989
rect 263877 47147 263905 47175
rect 263939 47147 263967 47175
rect 264001 47147 264029 47175
rect 264063 47147 264091 47175
rect 263877 47085 263905 47113
rect 263939 47085 263967 47113
rect 264001 47085 264029 47113
rect 264063 47085 264091 47113
rect 263877 47023 263905 47051
rect 263939 47023 263967 47051
rect 264001 47023 264029 47051
rect 264063 47023 264091 47051
rect 263877 46961 263905 46989
rect 263939 46961 263967 46989
rect 264001 46961 264029 46989
rect 264063 46961 264091 46989
rect 250377 41147 250405 41175
rect 250439 41147 250467 41175
rect 250501 41147 250529 41175
rect 250563 41147 250591 41175
rect 250377 41085 250405 41113
rect 250439 41085 250467 41113
rect 250501 41085 250529 41113
rect 250563 41085 250591 41113
rect 250377 41023 250405 41051
rect 250439 41023 250467 41051
rect 250501 41023 250529 41051
rect 250563 41023 250591 41051
rect 250377 40961 250405 40989
rect 250439 40961 250467 40989
rect 250501 40961 250529 40989
rect 250563 40961 250591 40989
rect 261699 41147 261727 41175
rect 261761 41147 261789 41175
rect 261699 41085 261727 41113
rect 261761 41085 261789 41113
rect 261699 41023 261727 41051
rect 261761 41023 261789 41051
rect 261699 40961 261727 40989
rect 261761 40961 261789 40989
rect 254019 38147 254047 38175
rect 254081 38147 254109 38175
rect 254019 38085 254047 38113
rect 254081 38085 254109 38113
rect 254019 38023 254047 38051
rect 254081 38023 254109 38051
rect 254019 37961 254047 37989
rect 254081 37961 254109 37989
rect 263877 38147 263905 38175
rect 263939 38147 263967 38175
rect 264001 38147 264029 38175
rect 264063 38147 264091 38175
rect 263877 38085 263905 38113
rect 263939 38085 263967 38113
rect 264001 38085 264029 38113
rect 264063 38085 264091 38113
rect 263877 38023 263905 38051
rect 263939 38023 263967 38051
rect 264001 38023 264029 38051
rect 264063 38023 264091 38051
rect 263877 37961 263905 37989
rect 263939 37961 263967 37989
rect 264001 37961 264029 37989
rect 264063 37961 264091 37989
rect 250377 32147 250405 32175
rect 250439 32147 250467 32175
rect 250501 32147 250529 32175
rect 250563 32147 250591 32175
rect 250377 32085 250405 32113
rect 250439 32085 250467 32113
rect 250501 32085 250529 32113
rect 250563 32085 250591 32113
rect 250377 32023 250405 32051
rect 250439 32023 250467 32051
rect 250501 32023 250529 32051
rect 250563 32023 250591 32051
rect 250377 31961 250405 31989
rect 250439 31961 250467 31989
rect 250501 31961 250529 31989
rect 250563 31961 250591 31989
rect 261699 32147 261727 32175
rect 261761 32147 261789 32175
rect 261699 32085 261727 32113
rect 261761 32085 261789 32113
rect 261699 32023 261727 32051
rect 261761 32023 261789 32051
rect 261699 31961 261727 31989
rect 261761 31961 261789 31989
rect 254019 29147 254047 29175
rect 254081 29147 254109 29175
rect 254019 29085 254047 29113
rect 254081 29085 254109 29113
rect 254019 29023 254047 29051
rect 254081 29023 254109 29051
rect 254019 28961 254047 28989
rect 254081 28961 254109 28989
rect 263877 29147 263905 29175
rect 263939 29147 263967 29175
rect 264001 29147 264029 29175
rect 264063 29147 264091 29175
rect 263877 29085 263905 29113
rect 263939 29085 263967 29113
rect 264001 29085 264029 29113
rect 264063 29085 264091 29113
rect 263877 29023 263905 29051
rect 263939 29023 263967 29051
rect 264001 29023 264029 29051
rect 264063 29023 264091 29051
rect 263877 28961 263905 28989
rect 263939 28961 263967 28989
rect 264001 28961 264029 28989
rect 264063 28961 264091 28989
rect 250377 23147 250405 23175
rect 250439 23147 250467 23175
rect 250501 23147 250529 23175
rect 250563 23147 250591 23175
rect 250377 23085 250405 23113
rect 250439 23085 250467 23113
rect 250501 23085 250529 23113
rect 250563 23085 250591 23113
rect 250377 23023 250405 23051
rect 250439 23023 250467 23051
rect 250501 23023 250529 23051
rect 250563 23023 250591 23051
rect 250377 22961 250405 22989
rect 250439 22961 250467 22989
rect 250501 22961 250529 22989
rect 250563 22961 250591 22989
rect 261699 23147 261727 23175
rect 261761 23147 261789 23175
rect 261699 23085 261727 23113
rect 261761 23085 261789 23113
rect 261699 23023 261727 23051
rect 261761 23023 261789 23051
rect 261699 22961 261727 22989
rect 261761 22961 261789 22989
rect 254019 20147 254047 20175
rect 254081 20147 254109 20175
rect 254019 20085 254047 20113
rect 254081 20085 254109 20113
rect 254019 20023 254047 20051
rect 254081 20023 254109 20051
rect 254019 19961 254047 19989
rect 254081 19961 254109 19989
rect 263877 20147 263905 20175
rect 263939 20147 263967 20175
rect 264001 20147 264029 20175
rect 264063 20147 264091 20175
rect 263877 20085 263905 20113
rect 263939 20085 263967 20113
rect 264001 20085 264029 20113
rect 264063 20085 264091 20113
rect 263877 20023 263905 20051
rect 263939 20023 263967 20051
rect 264001 20023 264029 20051
rect 264063 20023 264091 20051
rect 263877 19961 263905 19989
rect 263939 19961 263967 19989
rect 264001 19961 264029 19989
rect 264063 19961 264091 19989
rect 250377 14147 250405 14175
rect 250439 14147 250467 14175
rect 250501 14147 250529 14175
rect 250563 14147 250591 14175
rect 250377 14085 250405 14113
rect 250439 14085 250467 14113
rect 250501 14085 250529 14113
rect 250563 14085 250591 14113
rect 250377 14023 250405 14051
rect 250439 14023 250467 14051
rect 250501 14023 250529 14051
rect 250563 14023 250591 14051
rect 250377 13961 250405 13989
rect 250439 13961 250467 13989
rect 250501 13961 250529 13989
rect 250563 13961 250591 13989
rect 261699 14147 261727 14175
rect 261761 14147 261789 14175
rect 261699 14085 261727 14113
rect 261761 14085 261789 14113
rect 261699 14023 261727 14051
rect 261761 14023 261789 14051
rect 261699 13961 261727 13989
rect 261761 13961 261789 13989
rect 254019 11147 254047 11175
rect 254081 11147 254109 11175
rect 254019 11085 254047 11113
rect 254081 11085 254109 11113
rect 254019 11023 254047 11051
rect 254081 11023 254109 11051
rect 254019 10961 254047 10989
rect 254081 10961 254109 10989
rect 263877 11147 263905 11175
rect 263939 11147 263967 11175
rect 264001 11147 264029 11175
rect 264063 11147 264091 11175
rect 263877 11085 263905 11113
rect 263939 11085 263967 11113
rect 264001 11085 264029 11113
rect 264063 11085 264091 11113
rect 263877 11023 263905 11051
rect 263939 11023 263967 11051
rect 264001 11023 264029 11051
rect 264063 11023 264091 11051
rect 263877 10961 263905 10989
rect 263939 10961 263967 10989
rect 264001 10961 264029 10989
rect 264063 10961 264091 10989
rect 250377 5147 250405 5175
rect 250439 5147 250467 5175
rect 250501 5147 250529 5175
rect 250563 5147 250591 5175
rect 250377 5085 250405 5113
rect 250439 5085 250467 5113
rect 250501 5085 250529 5113
rect 250563 5085 250591 5113
rect 250377 5023 250405 5051
rect 250439 5023 250467 5051
rect 250501 5023 250529 5051
rect 250563 5023 250591 5051
rect 250377 4961 250405 4989
rect 250439 4961 250467 4989
rect 250501 4961 250529 4989
rect 250563 4961 250591 4989
rect 261699 5147 261727 5175
rect 261761 5147 261789 5175
rect 261699 5085 261727 5113
rect 261761 5085 261789 5113
rect 261699 5023 261727 5051
rect 261761 5023 261789 5051
rect 261699 4961 261727 4989
rect 261761 4961 261789 4989
rect 250377 -588 250405 -560
rect 250439 -588 250467 -560
rect 250501 -588 250529 -560
rect 250563 -588 250591 -560
rect 250377 -650 250405 -622
rect 250439 -650 250467 -622
rect 250501 -650 250529 -622
rect 250563 -650 250591 -622
rect 250377 -712 250405 -684
rect 250439 -712 250467 -684
rect 250501 -712 250529 -684
rect 250563 -712 250591 -684
rect 250377 -774 250405 -746
rect 250439 -774 250467 -746
rect 250501 -774 250529 -746
rect 250563 -774 250591 -746
rect 263877 2147 263905 2175
rect 263939 2147 263967 2175
rect 264001 2147 264029 2175
rect 264063 2147 264091 2175
rect 263877 2085 263905 2113
rect 263939 2085 263967 2113
rect 264001 2085 264029 2113
rect 264063 2085 264091 2113
rect 263877 2023 263905 2051
rect 263939 2023 263967 2051
rect 264001 2023 264029 2051
rect 264063 2023 264091 2051
rect 263877 1961 263905 1989
rect 263939 1961 263967 1989
rect 264001 1961 264029 1989
rect 264063 1961 264091 1989
rect 263877 -108 263905 -80
rect 263939 -108 263967 -80
rect 264001 -108 264029 -80
rect 264063 -108 264091 -80
rect 263877 -170 263905 -142
rect 263939 -170 263967 -142
rect 264001 -170 264029 -142
rect 264063 -170 264091 -142
rect 263877 -232 263905 -204
rect 263939 -232 263967 -204
rect 264001 -232 264029 -204
rect 264063 -232 264091 -204
rect 263877 -294 263905 -266
rect 263939 -294 263967 -266
rect 264001 -294 264029 -266
rect 264063 -294 264091 -266
rect 265737 299058 265765 299086
rect 265799 299058 265827 299086
rect 265861 299058 265889 299086
rect 265923 299058 265951 299086
rect 265737 298996 265765 299024
rect 265799 298996 265827 299024
rect 265861 298996 265889 299024
rect 265923 298996 265951 299024
rect 265737 298934 265765 298962
rect 265799 298934 265827 298962
rect 265861 298934 265889 298962
rect 265923 298934 265951 298962
rect 265737 298872 265765 298900
rect 265799 298872 265827 298900
rect 265861 298872 265889 298900
rect 265923 298872 265951 298900
rect 265737 293147 265765 293175
rect 265799 293147 265827 293175
rect 265861 293147 265889 293175
rect 265923 293147 265951 293175
rect 265737 293085 265765 293113
rect 265799 293085 265827 293113
rect 265861 293085 265889 293113
rect 265923 293085 265951 293113
rect 265737 293023 265765 293051
rect 265799 293023 265827 293051
rect 265861 293023 265889 293051
rect 265923 293023 265951 293051
rect 265737 292961 265765 292989
rect 265799 292961 265827 292989
rect 265861 292961 265889 292989
rect 265923 292961 265951 292989
rect 265737 284147 265765 284175
rect 265799 284147 265827 284175
rect 265861 284147 265889 284175
rect 265923 284147 265951 284175
rect 265737 284085 265765 284113
rect 265799 284085 265827 284113
rect 265861 284085 265889 284113
rect 265923 284085 265951 284113
rect 265737 284023 265765 284051
rect 265799 284023 265827 284051
rect 265861 284023 265889 284051
rect 265923 284023 265951 284051
rect 265737 283961 265765 283989
rect 265799 283961 265827 283989
rect 265861 283961 265889 283989
rect 265923 283961 265951 283989
rect 265737 275147 265765 275175
rect 265799 275147 265827 275175
rect 265861 275147 265889 275175
rect 265923 275147 265951 275175
rect 265737 275085 265765 275113
rect 265799 275085 265827 275113
rect 265861 275085 265889 275113
rect 265923 275085 265951 275113
rect 265737 275023 265765 275051
rect 265799 275023 265827 275051
rect 265861 275023 265889 275051
rect 265923 275023 265951 275051
rect 265737 274961 265765 274989
rect 265799 274961 265827 274989
rect 265861 274961 265889 274989
rect 265923 274961 265951 274989
rect 265737 266147 265765 266175
rect 265799 266147 265827 266175
rect 265861 266147 265889 266175
rect 265923 266147 265951 266175
rect 265737 266085 265765 266113
rect 265799 266085 265827 266113
rect 265861 266085 265889 266113
rect 265923 266085 265951 266113
rect 265737 266023 265765 266051
rect 265799 266023 265827 266051
rect 265861 266023 265889 266051
rect 265923 266023 265951 266051
rect 265737 265961 265765 265989
rect 265799 265961 265827 265989
rect 265861 265961 265889 265989
rect 265923 265961 265951 265989
rect 265737 257147 265765 257175
rect 265799 257147 265827 257175
rect 265861 257147 265889 257175
rect 265923 257147 265951 257175
rect 265737 257085 265765 257113
rect 265799 257085 265827 257113
rect 265861 257085 265889 257113
rect 265923 257085 265951 257113
rect 265737 257023 265765 257051
rect 265799 257023 265827 257051
rect 265861 257023 265889 257051
rect 265923 257023 265951 257051
rect 265737 256961 265765 256989
rect 265799 256961 265827 256989
rect 265861 256961 265889 256989
rect 265923 256961 265951 256989
rect 265737 248147 265765 248175
rect 265799 248147 265827 248175
rect 265861 248147 265889 248175
rect 265923 248147 265951 248175
rect 265737 248085 265765 248113
rect 265799 248085 265827 248113
rect 265861 248085 265889 248113
rect 265923 248085 265951 248113
rect 265737 248023 265765 248051
rect 265799 248023 265827 248051
rect 265861 248023 265889 248051
rect 265923 248023 265951 248051
rect 265737 247961 265765 247989
rect 265799 247961 265827 247989
rect 265861 247961 265889 247989
rect 265923 247961 265951 247989
rect 265737 239147 265765 239175
rect 265799 239147 265827 239175
rect 265861 239147 265889 239175
rect 265923 239147 265951 239175
rect 265737 239085 265765 239113
rect 265799 239085 265827 239113
rect 265861 239085 265889 239113
rect 265923 239085 265951 239113
rect 265737 239023 265765 239051
rect 265799 239023 265827 239051
rect 265861 239023 265889 239051
rect 265923 239023 265951 239051
rect 265737 238961 265765 238989
rect 265799 238961 265827 238989
rect 265861 238961 265889 238989
rect 265923 238961 265951 238989
rect 265737 230147 265765 230175
rect 265799 230147 265827 230175
rect 265861 230147 265889 230175
rect 265923 230147 265951 230175
rect 265737 230085 265765 230113
rect 265799 230085 265827 230113
rect 265861 230085 265889 230113
rect 265923 230085 265951 230113
rect 265737 230023 265765 230051
rect 265799 230023 265827 230051
rect 265861 230023 265889 230051
rect 265923 230023 265951 230051
rect 265737 229961 265765 229989
rect 265799 229961 265827 229989
rect 265861 229961 265889 229989
rect 265923 229961 265951 229989
rect 265737 221147 265765 221175
rect 265799 221147 265827 221175
rect 265861 221147 265889 221175
rect 265923 221147 265951 221175
rect 265737 221085 265765 221113
rect 265799 221085 265827 221113
rect 265861 221085 265889 221113
rect 265923 221085 265951 221113
rect 265737 221023 265765 221051
rect 265799 221023 265827 221051
rect 265861 221023 265889 221051
rect 265923 221023 265951 221051
rect 265737 220961 265765 220989
rect 265799 220961 265827 220989
rect 265861 220961 265889 220989
rect 265923 220961 265951 220989
rect 265737 212147 265765 212175
rect 265799 212147 265827 212175
rect 265861 212147 265889 212175
rect 265923 212147 265951 212175
rect 265737 212085 265765 212113
rect 265799 212085 265827 212113
rect 265861 212085 265889 212113
rect 265923 212085 265951 212113
rect 265737 212023 265765 212051
rect 265799 212023 265827 212051
rect 265861 212023 265889 212051
rect 265923 212023 265951 212051
rect 265737 211961 265765 211989
rect 265799 211961 265827 211989
rect 265861 211961 265889 211989
rect 265923 211961 265951 211989
rect 265737 203147 265765 203175
rect 265799 203147 265827 203175
rect 265861 203147 265889 203175
rect 265923 203147 265951 203175
rect 265737 203085 265765 203113
rect 265799 203085 265827 203113
rect 265861 203085 265889 203113
rect 265923 203085 265951 203113
rect 265737 203023 265765 203051
rect 265799 203023 265827 203051
rect 265861 203023 265889 203051
rect 265923 203023 265951 203051
rect 265737 202961 265765 202989
rect 265799 202961 265827 202989
rect 265861 202961 265889 202989
rect 265923 202961 265951 202989
rect 265737 194147 265765 194175
rect 265799 194147 265827 194175
rect 265861 194147 265889 194175
rect 265923 194147 265951 194175
rect 265737 194085 265765 194113
rect 265799 194085 265827 194113
rect 265861 194085 265889 194113
rect 265923 194085 265951 194113
rect 265737 194023 265765 194051
rect 265799 194023 265827 194051
rect 265861 194023 265889 194051
rect 265923 194023 265951 194051
rect 265737 193961 265765 193989
rect 265799 193961 265827 193989
rect 265861 193961 265889 193989
rect 265923 193961 265951 193989
rect 265737 185147 265765 185175
rect 265799 185147 265827 185175
rect 265861 185147 265889 185175
rect 265923 185147 265951 185175
rect 265737 185085 265765 185113
rect 265799 185085 265827 185113
rect 265861 185085 265889 185113
rect 265923 185085 265951 185113
rect 265737 185023 265765 185051
rect 265799 185023 265827 185051
rect 265861 185023 265889 185051
rect 265923 185023 265951 185051
rect 265737 184961 265765 184989
rect 265799 184961 265827 184989
rect 265861 184961 265889 184989
rect 265923 184961 265951 184989
rect 265737 176147 265765 176175
rect 265799 176147 265827 176175
rect 265861 176147 265889 176175
rect 265923 176147 265951 176175
rect 265737 176085 265765 176113
rect 265799 176085 265827 176113
rect 265861 176085 265889 176113
rect 265923 176085 265951 176113
rect 265737 176023 265765 176051
rect 265799 176023 265827 176051
rect 265861 176023 265889 176051
rect 265923 176023 265951 176051
rect 265737 175961 265765 175989
rect 265799 175961 265827 175989
rect 265861 175961 265889 175989
rect 265923 175961 265951 175989
rect 279237 298578 279265 298606
rect 279299 298578 279327 298606
rect 279361 298578 279389 298606
rect 279423 298578 279451 298606
rect 279237 298516 279265 298544
rect 279299 298516 279327 298544
rect 279361 298516 279389 298544
rect 279423 298516 279451 298544
rect 279237 298454 279265 298482
rect 279299 298454 279327 298482
rect 279361 298454 279389 298482
rect 279423 298454 279451 298482
rect 279237 298392 279265 298420
rect 279299 298392 279327 298420
rect 279361 298392 279389 298420
rect 279423 298392 279451 298420
rect 279237 290147 279265 290175
rect 279299 290147 279327 290175
rect 279361 290147 279389 290175
rect 279423 290147 279451 290175
rect 279237 290085 279265 290113
rect 279299 290085 279327 290113
rect 279361 290085 279389 290113
rect 279423 290085 279451 290113
rect 279237 290023 279265 290051
rect 279299 290023 279327 290051
rect 279361 290023 279389 290051
rect 279423 290023 279451 290051
rect 279237 289961 279265 289989
rect 279299 289961 279327 289989
rect 279361 289961 279389 289989
rect 279423 289961 279451 289989
rect 279237 281147 279265 281175
rect 279299 281147 279327 281175
rect 279361 281147 279389 281175
rect 279423 281147 279451 281175
rect 279237 281085 279265 281113
rect 279299 281085 279327 281113
rect 279361 281085 279389 281113
rect 279423 281085 279451 281113
rect 279237 281023 279265 281051
rect 279299 281023 279327 281051
rect 279361 281023 279389 281051
rect 279423 281023 279451 281051
rect 279237 280961 279265 280989
rect 279299 280961 279327 280989
rect 279361 280961 279389 280989
rect 279423 280961 279451 280989
rect 279237 272147 279265 272175
rect 279299 272147 279327 272175
rect 279361 272147 279389 272175
rect 279423 272147 279451 272175
rect 279237 272085 279265 272113
rect 279299 272085 279327 272113
rect 279361 272085 279389 272113
rect 279423 272085 279451 272113
rect 279237 272023 279265 272051
rect 279299 272023 279327 272051
rect 279361 272023 279389 272051
rect 279423 272023 279451 272051
rect 279237 271961 279265 271989
rect 279299 271961 279327 271989
rect 279361 271961 279389 271989
rect 279423 271961 279451 271989
rect 279237 263147 279265 263175
rect 279299 263147 279327 263175
rect 279361 263147 279389 263175
rect 279423 263147 279451 263175
rect 279237 263085 279265 263113
rect 279299 263085 279327 263113
rect 279361 263085 279389 263113
rect 279423 263085 279451 263113
rect 279237 263023 279265 263051
rect 279299 263023 279327 263051
rect 279361 263023 279389 263051
rect 279423 263023 279451 263051
rect 279237 262961 279265 262989
rect 279299 262961 279327 262989
rect 279361 262961 279389 262989
rect 279423 262961 279451 262989
rect 279237 254147 279265 254175
rect 279299 254147 279327 254175
rect 279361 254147 279389 254175
rect 279423 254147 279451 254175
rect 279237 254085 279265 254113
rect 279299 254085 279327 254113
rect 279361 254085 279389 254113
rect 279423 254085 279451 254113
rect 279237 254023 279265 254051
rect 279299 254023 279327 254051
rect 279361 254023 279389 254051
rect 279423 254023 279451 254051
rect 279237 253961 279265 253989
rect 279299 253961 279327 253989
rect 279361 253961 279389 253989
rect 279423 253961 279451 253989
rect 279237 245147 279265 245175
rect 279299 245147 279327 245175
rect 279361 245147 279389 245175
rect 279423 245147 279451 245175
rect 279237 245085 279265 245113
rect 279299 245085 279327 245113
rect 279361 245085 279389 245113
rect 279423 245085 279451 245113
rect 279237 245023 279265 245051
rect 279299 245023 279327 245051
rect 279361 245023 279389 245051
rect 279423 245023 279451 245051
rect 279237 244961 279265 244989
rect 279299 244961 279327 244989
rect 279361 244961 279389 244989
rect 279423 244961 279451 244989
rect 279237 236147 279265 236175
rect 279299 236147 279327 236175
rect 279361 236147 279389 236175
rect 279423 236147 279451 236175
rect 279237 236085 279265 236113
rect 279299 236085 279327 236113
rect 279361 236085 279389 236113
rect 279423 236085 279451 236113
rect 279237 236023 279265 236051
rect 279299 236023 279327 236051
rect 279361 236023 279389 236051
rect 279423 236023 279451 236051
rect 279237 235961 279265 235989
rect 279299 235961 279327 235989
rect 279361 235961 279389 235989
rect 279423 235961 279451 235989
rect 279237 227147 279265 227175
rect 279299 227147 279327 227175
rect 279361 227147 279389 227175
rect 279423 227147 279451 227175
rect 279237 227085 279265 227113
rect 279299 227085 279327 227113
rect 279361 227085 279389 227113
rect 279423 227085 279451 227113
rect 279237 227023 279265 227051
rect 279299 227023 279327 227051
rect 279361 227023 279389 227051
rect 279423 227023 279451 227051
rect 279237 226961 279265 226989
rect 279299 226961 279327 226989
rect 279361 226961 279389 226989
rect 279423 226961 279451 226989
rect 279237 218147 279265 218175
rect 279299 218147 279327 218175
rect 279361 218147 279389 218175
rect 279423 218147 279451 218175
rect 279237 218085 279265 218113
rect 279299 218085 279327 218113
rect 279361 218085 279389 218113
rect 279423 218085 279451 218113
rect 279237 218023 279265 218051
rect 279299 218023 279327 218051
rect 279361 218023 279389 218051
rect 279423 218023 279451 218051
rect 279237 217961 279265 217989
rect 279299 217961 279327 217989
rect 279361 217961 279389 217989
rect 279423 217961 279451 217989
rect 279237 209147 279265 209175
rect 279299 209147 279327 209175
rect 279361 209147 279389 209175
rect 279423 209147 279451 209175
rect 279237 209085 279265 209113
rect 279299 209085 279327 209113
rect 279361 209085 279389 209113
rect 279423 209085 279451 209113
rect 279237 209023 279265 209051
rect 279299 209023 279327 209051
rect 279361 209023 279389 209051
rect 279423 209023 279451 209051
rect 279237 208961 279265 208989
rect 279299 208961 279327 208989
rect 279361 208961 279389 208989
rect 279423 208961 279451 208989
rect 279237 200147 279265 200175
rect 279299 200147 279327 200175
rect 279361 200147 279389 200175
rect 279423 200147 279451 200175
rect 279237 200085 279265 200113
rect 279299 200085 279327 200113
rect 279361 200085 279389 200113
rect 279423 200085 279451 200113
rect 279237 200023 279265 200051
rect 279299 200023 279327 200051
rect 279361 200023 279389 200051
rect 279423 200023 279451 200051
rect 279237 199961 279265 199989
rect 279299 199961 279327 199989
rect 279361 199961 279389 199989
rect 279423 199961 279451 199989
rect 279237 191147 279265 191175
rect 279299 191147 279327 191175
rect 279361 191147 279389 191175
rect 279423 191147 279451 191175
rect 279237 191085 279265 191113
rect 279299 191085 279327 191113
rect 279361 191085 279389 191113
rect 279423 191085 279451 191113
rect 279237 191023 279265 191051
rect 279299 191023 279327 191051
rect 279361 191023 279389 191051
rect 279423 191023 279451 191051
rect 279237 190961 279265 190989
rect 279299 190961 279327 190989
rect 279361 190961 279389 190989
rect 279423 190961 279451 190989
rect 279237 182147 279265 182175
rect 279299 182147 279327 182175
rect 279361 182147 279389 182175
rect 279423 182147 279451 182175
rect 279237 182085 279265 182113
rect 279299 182085 279327 182113
rect 279361 182085 279389 182113
rect 279423 182085 279451 182113
rect 279237 182023 279265 182051
rect 279299 182023 279327 182051
rect 279361 182023 279389 182051
rect 279423 182023 279451 182051
rect 279237 181961 279265 181989
rect 279299 181961 279327 181989
rect 279361 181961 279389 181989
rect 279423 181961 279451 181989
rect 269379 173147 269407 173175
rect 269441 173147 269469 173175
rect 269379 173085 269407 173113
rect 269441 173085 269469 173113
rect 269379 173023 269407 173051
rect 269441 173023 269469 173051
rect 269379 172961 269407 172989
rect 269441 172961 269469 172989
rect 279237 173147 279265 173175
rect 279299 173147 279327 173175
rect 279361 173147 279389 173175
rect 279423 173147 279451 173175
rect 279237 173085 279265 173113
rect 279299 173085 279327 173113
rect 279361 173085 279389 173113
rect 279423 173085 279451 173113
rect 279237 173023 279265 173051
rect 279299 173023 279327 173051
rect 279361 173023 279389 173051
rect 279423 173023 279451 173051
rect 279237 172961 279265 172989
rect 279299 172961 279327 172989
rect 279361 172961 279389 172989
rect 279423 172961 279451 172989
rect 265737 167147 265765 167175
rect 265799 167147 265827 167175
rect 265861 167147 265889 167175
rect 265923 167147 265951 167175
rect 265737 167085 265765 167113
rect 265799 167085 265827 167113
rect 265861 167085 265889 167113
rect 265923 167085 265951 167113
rect 265737 167023 265765 167051
rect 265799 167023 265827 167051
rect 265861 167023 265889 167051
rect 265923 167023 265951 167051
rect 265737 166961 265765 166989
rect 265799 166961 265827 166989
rect 265861 166961 265889 166989
rect 265923 166961 265951 166989
rect 277059 167147 277087 167175
rect 277121 167147 277149 167175
rect 277059 167085 277087 167113
rect 277121 167085 277149 167113
rect 277059 167023 277087 167051
rect 277121 167023 277149 167051
rect 277059 166961 277087 166989
rect 277121 166961 277149 166989
rect 269379 164147 269407 164175
rect 269441 164147 269469 164175
rect 269379 164085 269407 164113
rect 269441 164085 269469 164113
rect 269379 164023 269407 164051
rect 269441 164023 269469 164051
rect 269379 163961 269407 163989
rect 269441 163961 269469 163989
rect 279237 164147 279265 164175
rect 279299 164147 279327 164175
rect 279361 164147 279389 164175
rect 279423 164147 279451 164175
rect 279237 164085 279265 164113
rect 279299 164085 279327 164113
rect 279361 164085 279389 164113
rect 279423 164085 279451 164113
rect 279237 164023 279265 164051
rect 279299 164023 279327 164051
rect 279361 164023 279389 164051
rect 279423 164023 279451 164051
rect 279237 163961 279265 163989
rect 279299 163961 279327 163989
rect 279361 163961 279389 163989
rect 279423 163961 279451 163989
rect 265737 158147 265765 158175
rect 265799 158147 265827 158175
rect 265861 158147 265889 158175
rect 265923 158147 265951 158175
rect 265737 158085 265765 158113
rect 265799 158085 265827 158113
rect 265861 158085 265889 158113
rect 265923 158085 265951 158113
rect 265737 158023 265765 158051
rect 265799 158023 265827 158051
rect 265861 158023 265889 158051
rect 265923 158023 265951 158051
rect 265737 157961 265765 157989
rect 265799 157961 265827 157989
rect 265861 157961 265889 157989
rect 265923 157961 265951 157989
rect 277059 158147 277087 158175
rect 277121 158147 277149 158175
rect 277059 158085 277087 158113
rect 277121 158085 277149 158113
rect 277059 158023 277087 158051
rect 277121 158023 277149 158051
rect 277059 157961 277087 157989
rect 277121 157961 277149 157989
rect 269379 155147 269407 155175
rect 269441 155147 269469 155175
rect 269379 155085 269407 155113
rect 269441 155085 269469 155113
rect 269379 155023 269407 155051
rect 269441 155023 269469 155051
rect 269379 154961 269407 154989
rect 269441 154961 269469 154989
rect 279237 155147 279265 155175
rect 279299 155147 279327 155175
rect 279361 155147 279389 155175
rect 279423 155147 279451 155175
rect 279237 155085 279265 155113
rect 279299 155085 279327 155113
rect 279361 155085 279389 155113
rect 279423 155085 279451 155113
rect 279237 155023 279265 155051
rect 279299 155023 279327 155051
rect 279361 155023 279389 155051
rect 279423 155023 279451 155051
rect 279237 154961 279265 154989
rect 279299 154961 279327 154989
rect 279361 154961 279389 154989
rect 279423 154961 279451 154989
rect 265737 149147 265765 149175
rect 265799 149147 265827 149175
rect 265861 149147 265889 149175
rect 265923 149147 265951 149175
rect 265737 149085 265765 149113
rect 265799 149085 265827 149113
rect 265861 149085 265889 149113
rect 265923 149085 265951 149113
rect 265737 149023 265765 149051
rect 265799 149023 265827 149051
rect 265861 149023 265889 149051
rect 265923 149023 265951 149051
rect 265737 148961 265765 148989
rect 265799 148961 265827 148989
rect 265861 148961 265889 148989
rect 265923 148961 265951 148989
rect 277059 149147 277087 149175
rect 277121 149147 277149 149175
rect 277059 149085 277087 149113
rect 277121 149085 277149 149113
rect 277059 149023 277087 149051
rect 277121 149023 277149 149051
rect 277059 148961 277087 148989
rect 277121 148961 277149 148989
rect 269379 146147 269407 146175
rect 269441 146147 269469 146175
rect 269379 146085 269407 146113
rect 269441 146085 269469 146113
rect 269379 146023 269407 146051
rect 269441 146023 269469 146051
rect 269379 145961 269407 145989
rect 269441 145961 269469 145989
rect 279237 146147 279265 146175
rect 279299 146147 279327 146175
rect 279361 146147 279389 146175
rect 279423 146147 279451 146175
rect 279237 146085 279265 146113
rect 279299 146085 279327 146113
rect 279361 146085 279389 146113
rect 279423 146085 279451 146113
rect 279237 146023 279265 146051
rect 279299 146023 279327 146051
rect 279361 146023 279389 146051
rect 279423 146023 279451 146051
rect 279237 145961 279265 145989
rect 279299 145961 279327 145989
rect 279361 145961 279389 145989
rect 279423 145961 279451 145989
rect 265737 140147 265765 140175
rect 265799 140147 265827 140175
rect 265861 140147 265889 140175
rect 265923 140147 265951 140175
rect 265737 140085 265765 140113
rect 265799 140085 265827 140113
rect 265861 140085 265889 140113
rect 265923 140085 265951 140113
rect 265737 140023 265765 140051
rect 265799 140023 265827 140051
rect 265861 140023 265889 140051
rect 265923 140023 265951 140051
rect 265737 139961 265765 139989
rect 265799 139961 265827 139989
rect 265861 139961 265889 139989
rect 265923 139961 265951 139989
rect 277059 140147 277087 140175
rect 277121 140147 277149 140175
rect 277059 140085 277087 140113
rect 277121 140085 277149 140113
rect 277059 140023 277087 140051
rect 277121 140023 277149 140051
rect 277059 139961 277087 139989
rect 277121 139961 277149 139989
rect 269379 137147 269407 137175
rect 269441 137147 269469 137175
rect 269379 137085 269407 137113
rect 269441 137085 269469 137113
rect 269379 137023 269407 137051
rect 269441 137023 269469 137051
rect 269379 136961 269407 136989
rect 269441 136961 269469 136989
rect 279237 137147 279265 137175
rect 279299 137147 279327 137175
rect 279361 137147 279389 137175
rect 279423 137147 279451 137175
rect 279237 137085 279265 137113
rect 279299 137085 279327 137113
rect 279361 137085 279389 137113
rect 279423 137085 279451 137113
rect 279237 137023 279265 137051
rect 279299 137023 279327 137051
rect 279361 137023 279389 137051
rect 279423 137023 279451 137051
rect 279237 136961 279265 136989
rect 279299 136961 279327 136989
rect 279361 136961 279389 136989
rect 279423 136961 279451 136989
rect 265737 131147 265765 131175
rect 265799 131147 265827 131175
rect 265861 131147 265889 131175
rect 265923 131147 265951 131175
rect 265737 131085 265765 131113
rect 265799 131085 265827 131113
rect 265861 131085 265889 131113
rect 265923 131085 265951 131113
rect 265737 131023 265765 131051
rect 265799 131023 265827 131051
rect 265861 131023 265889 131051
rect 265923 131023 265951 131051
rect 265737 130961 265765 130989
rect 265799 130961 265827 130989
rect 265861 130961 265889 130989
rect 265923 130961 265951 130989
rect 277059 131147 277087 131175
rect 277121 131147 277149 131175
rect 277059 131085 277087 131113
rect 277121 131085 277149 131113
rect 277059 131023 277087 131051
rect 277121 131023 277149 131051
rect 277059 130961 277087 130989
rect 277121 130961 277149 130989
rect 269379 128147 269407 128175
rect 269441 128147 269469 128175
rect 269379 128085 269407 128113
rect 269441 128085 269469 128113
rect 269379 128023 269407 128051
rect 269441 128023 269469 128051
rect 269379 127961 269407 127989
rect 269441 127961 269469 127989
rect 279237 128147 279265 128175
rect 279299 128147 279327 128175
rect 279361 128147 279389 128175
rect 279423 128147 279451 128175
rect 279237 128085 279265 128113
rect 279299 128085 279327 128113
rect 279361 128085 279389 128113
rect 279423 128085 279451 128113
rect 279237 128023 279265 128051
rect 279299 128023 279327 128051
rect 279361 128023 279389 128051
rect 279423 128023 279451 128051
rect 279237 127961 279265 127989
rect 279299 127961 279327 127989
rect 279361 127961 279389 127989
rect 279423 127961 279451 127989
rect 265737 122147 265765 122175
rect 265799 122147 265827 122175
rect 265861 122147 265889 122175
rect 265923 122147 265951 122175
rect 265737 122085 265765 122113
rect 265799 122085 265827 122113
rect 265861 122085 265889 122113
rect 265923 122085 265951 122113
rect 265737 122023 265765 122051
rect 265799 122023 265827 122051
rect 265861 122023 265889 122051
rect 265923 122023 265951 122051
rect 265737 121961 265765 121989
rect 265799 121961 265827 121989
rect 265861 121961 265889 121989
rect 265923 121961 265951 121989
rect 277059 122147 277087 122175
rect 277121 122147 277149 122175
rect 277059 122085 277087 122113
rect 277121 122085 277149 122113
rect 277059 122023 277087 122051
rect 277121 122023 277149 122051
rect 277059 121961 277087 121989
rect 277121 121961 277149 121989
rect 269379 119147 269407 119175
rect 269441 119147 269469 119175
rect 269379 119085 269407 119113
rect 269441 119085 269469 119113
rect 269379 119023 269407 119051
rect 269441 119023 269469 119051
rect 269379 118961 269407 118989
rect 269441 118961 269469 118989
rect 279237 119147 279265 119175
rect 279299 119147 279327 119175
rect 279361 119147 279389 119175
rect 279423 119147 279451 119175
rect 279237 119085 279265 119113
rect 279299 119085 279327 119113
rect 279361 119085 279389 119113
rect 279423 119085 279451 119113
rect 279237 119023 279265 119051
rect 279299 119023 279327 119051
rect 279361 119023 279389 119051
rect 279423 119023 279451 119051
rect 279237 118961 279265 118989
rect 279299 118961 279327 118989
rect 279361 118961 279389 118989
rect 279423 118961 279451 118989
rect 265737 113147 265765 113175
rect 265799 113147 265827 113175
rect 265861 113147 265889 113175
rect 265923 113147 265951 113175
rect 265737 113085 265765 113113
rect 265799 113085 265827 113113
rect 265861 113085 265889 113113
rect 265923 113085 265951 113113
rect 265737 113023 265765 113051
rect 265799 113023 265827 113051
rect 265861 113023 265889 113051
rect 265923 113023 265951 113051
rect 265737 112961 265765 112989
rect 265799 112961 265827 112989
rect 265861 112961 265889 112989
rect 265923 112961 265951 112989
rect 277059 113147 277087 113175
rect 277121 113147 277149 113175
rect 277059 113085 277087 113113
rect 277121 113085 277149 113113
rect 277059 113023 277087 113051
rect 277121 113023 277149 113051
rect 277059 112961 277087 112989
rect 277121 112961 277149 112989
rect 269379 110147 269407 110175
rect 269441 110147 269469 110175
rect 269379 110085 269407 110113
rect 269441 110085 269469 110113
rect 269379 110023 269407 110051
rect 269441 110023 269469 110051
rect 269379 109961 269407 109989
rect 269441 109961 269469 109989
rect 279237 110147 279265 110175
rect 279299 110147 279327 110175
rect 279361 110147 279389 110175
rect 279423 110147 279451 110175
rect 279237 110085 279265 110113
rect 279299 110085 279327 110113
rect 279361 110085 279389 110113
rect 279423 110085 279451 110113
rect 279237 110023 279265 110051
rect 279299 110023 279327 110051
rect 279361 110023 279389 110051
rect 279423 110023 279451 110051
rect 279237 109961 279265 109989
rect 279299 109961 279327 109989
rect 279361 109961 279389 109989
rect 279423 109961 279451 109989
rect 265737 104147 265765 104175
rect 265799 104147 265827 104175
rect 265861 104147 265889 104175
rect 265923 104147 265951 104175
rect 265737 104085 265765 104113
rect 265799 104085 265827 104113
rect 265861 104085 265889 104113
rect 265923 104085 265951 104113
rect 265737 104023 265765 104051
rect 265799 104023 265827 104051
rect 265861 104023 265889 104051
rect 265923 104023 265951 104051
rect 265737 103961 265765 103989
rect 265799 103961 265827 103989
rect 265861 103961 265889 103989
rect 265923 103961 265951 103989
rect 277059 104147 277087 104175
rect 277121 104147 277149 104175
rect 277059 104085 277087 104113
rect 277121 104085 277149 104113
rect 277059 104023 277087 104051
rect 277121 104023 277149 104051
rect 277059 103961 277087 103989
rect 277121 103961 277149 103989
rect 269379 101147 269407 101175
rect 269441 101147 269469 101175
rect 269379 101085 269407 101113
rect 269441 101085 269469 101113
rect 269379 101023 269407 101051
rect 269441 101023 269469 101051
rect 269379 100961 269407 100989
rect 269441 100961 269469 100989
rect 279237 101147 279265 101175
rect 279299 101147 279327 101175
rect 279361 101147 279389 101175
rect 279423 101147 279451 101175
rect 279237 101085 279265 101113
rect 279299 101085 279327 101113
rect 279361 101085 279389 101113
rect 279423 101085 279451 101113
rect 279237 101023 279265 101051
rect 279299 101023 279327 101051
rect 279361 101023 279389 101051
rect 279423 101023 279451 101051
rect 279237 100961 279265 100989
rect 279299 100961 279327 100989
rect 279361 100961 279389 100989
rect 279423 100961 279451 100989
rect 265737 95147 265765 95175
rect 265799 95147 265827 95175
rect 265861 95147 265889 95175
rect 265923 95147 265951 95175
rect 265737 95085 265765 95113
rect 265799 95085 265827 95113
rect 265861 95085 265889 95113
rect 265923 95085 265951 95113
rect 265737 95023 265765 95051
rect 265799 95023 265827 95051
rect 265861 95023 265889 95051
rect 265923 95023 265951 95051
rect 265737 94961 265765 94989
rect 265799 94961 265827 94989
rect 265861 94961 265889 94989
rect 265923 94961 265951 94989
rect 277059 95147 277087 95175
rect 277121 95147 277149 95175
rect 277059 95085 277087 95113
rect 277121 95085 277149 95113
rect 277059 95023 277087 95051
rect 277121 95023 277149 95051
rect 277059 94961 277087 94989
rect 277121 94961 277149 94989
rect 269379 92147 269407 92175
rect 269441 92147 269469 92175
rect 269379 92085 269407 92113
rect 269441 92085 269469 92113
rect 269379 92023 269407 92051
rect 269441 92023 269469 92051
rect 269379 91961 269407 91989
rect 269441 91961 269469 91989
rect 279237 92147 279265 92175
rect 279299 92147 279327 92175
rect 279361 92147 279389 92175
rect 279423 92147 279451 92175
rect 279237 92085 279265 92113
rect 279299 92085 279327 92113
rect 279361 92085 279389 92113
rect 279423 92085 279451 92113
rect 279237 92023 279265 92051
rect 279299 92023 279327 92051
rect 279361 92023 279389 92051
rect 279423 92023 279451 92051
rect 279237 91961 279265 91989
rect 279299 91961 279327 91989
rect 279361 91961 279389 91989
rect 279423 91961 279451 91989
rect 265737 86147 265765 86175
rect 265799 86147 265827 86175
rect 265861 86147 265889 86175
rect 265923 86147 265951 86175
rect 265737 86085 265765 86113
rect 265799 86085 265827 86113
rect 265861 86085 265889 86113
rect 265923 86085 265951 86113
rect 265737 86023 265765 86051
rect 265799 86023 265827 86051
rect 265861 86023 265889 86051
rect 265923 86023 265951 86051
rect 265737 85961 265765 85989
rect 265799 85961 265827 85989
rect 265861 85961 265889 85989
rect 265923 85961 265951 85989
rect 277059 86147 277087 86175
rect 277121 86147 277149 86175
rect 277059 86085 277087 86113
rect 277121 86085 277149 86113
rect 277059 86023 277087 86051
rect 277121 86023 277149 86051
rect 277059 85961 277087 85989
rect 277121 85961 277149 85989
rect 269379 83147 269407 83175
rect 269441 83147 269469 83175
rect 269379 83085 269407 83113
rect 269441 83085 269469 83113
rect 269379 83023 269407 83051
rect 269441 83023 269469 83051
rect 269379 82961 269407 82989
rect 269441 82961 269469 82989
rect 279237 83147 279265 83175
rect 279299 83147 279327 83175
rect 279361 83147 279389 83175
rect 279423 83147 279451 83175
rect 279237 83085 279265 83113
rect 279299 83085 279327 83113
rect 279361 83085 279389 83113
rect 279423 83085 279451 83113
rect 279237 83023 279265 83051
rect 279299 83023 279327 83051
rect 279361 83023 279389 83051
rect 279423 83023 279451 83051
rect 279237 82961 279265 82989
rect 279299 82961 279327 82989
rect 279361 82961 279389 82989
rect 279423 82961 279451 82989
rect 265737 77147 265765 77175
rect 265799 77147 265827 77175
rect 265861 77147 265889 77175
rect 265923 77147 265951 77175
rect 265737 77085 265765 77113
rect 265799 77085 265827 77113
rect 265861 77085 265889 77113
rect 265923 77085 265951 77113
rect 265737 77023 265765 77051
rect 265799 77023 265827 77051
rect 265861 77023 265889 77051
rect 265923 77023 265951 77051
rect 265737 76961 265765 76989
rect 265799 76961 265827 76989
rect 265861 76961 265889 76989
rect 265923 76961 265951 76989
rect 277059 77147 277087 77175
rect 277121 77147 277149 77175
rect 277059 77085 277087 77113
rect 277121 77085 277149 77113
rect 277059 77023 277087 77051
rect 277121 77023 277149 77051
rect 277059 76961 277087 76989
rect 277121 76961 277149 76989
rect 269379 74147 269407 74175
rect 269441 74147 269469 74175
rect 269379 74085 269407 74113
rect 269441 74085 269469 74113
rect 269379 74023 269407 74051
rect 269441 74023 269469 74051
rect 269379 73961 269407 73989
rect 269441 73961 269469 73989
rect 279237 74147 279265 74175
rect 279299 74147 279327 74175
rect 279361 74147 279389 74175
rect 279423 74147 279451 74175
rect 279237 74085 279265 74113
rect 279299 74085 279327 74113
rect 279361 74085 279389 74113
rect 279423 74085 279451 74113
rect 279237 74023 279265 74051
rect 279299 74023 279327 74051
rect 279361 74023 279389 74051
rect 279423 74023 279451 74051
rect 279237 73961 279265 73989
rect 279299 73961 279327 73989
rect 279361 73961 279389 73989
rect 279423 73961 279451 73989
rect 265737 68147 265765 68175
rect 265799 68147 265827 68175
rect 265861 68147 265889 68175
rect 265923 68147 265951 68175
rect 265737 68085 265765 68113
rect 265799 68085 265827 68113
rect 265861 68085 265889 68113
rect 265923 68085 265951 68113
rect 265737 68023 265765 68051
rect 265799 68023 265827 68051
rect 265861 68023 265889 68051
rect 265923 68023 265951 68051
rect 265737 67961 265765 67989
rect 265799 67961 265827 67989
rect 265861 67961 265889 67989
rect 265923 67961 265951 67989
rect 277059 68147 277087 68175
rect 277121 68147 277149 68175
rect 277059 68085 277087 68113
rect 277121 68085 277149 68113
rect 277059 68023 277087 68051
rect 277121 68023 277149 68051
rect 277059 67961 277087 67989
rect 277121 67961 277149 67989
rect 269379 65147 269407 65175
rect 269441 65147 269469 65175
rect 269379 65085 269407 65113
rect 269441 65085 269469 65113
rect 269379 65023 269407 65051
rect 269441 65023 269469 65051
rect 269379 64961 269407 64989
rect 269441 64961 269469 64989
rect 279237 65147 279265 65175
rect 279299 65147 279327 65175
rect 279361 65147 279389 65175
rect 279423 65147 279451 65175
rect 279237 65085 279265 65113
rect 279299 65085 279327 65113
rect 279361 65085 279389 65113
rect 279423 65085 279451 65113
rect 279237 65023 279265 65051
rect 279299 65023 279327 65051
rect 279361 65023 279389 65051
rect 279423 65023 279451 65051
rect 279237 64961 279265 64989
rect 279299 64961 279327 64989
rect 279361 64961 279389 64989
rect 279423 64961 279451 64989
rect 265737 59147 265765 59175
rect 265799 59147 265827 59175
rect 265861 59147 265889 59175
rect 265923 59147 265951 59175
rect 265737 59085 265765 59113
rect 265799 59085 265827 59113
rect 265861 59085 265889 59113
rect 265923 59085 265951 59113
rect 265737 59023 265765 59051
rect 265799 59023 265827 59051
rect 265861 59023 265889 59051
rect 265923 59023 265951 59051
rect 265737 58961 265765 58989
rect 265799 58961 265827 58989
rect 265861 58961 265889 58989
rect 265923 58961 265951 58989
rect 277059 59147 277087 59175
rect 277121 59147 277149 59175
rect 277059 59085 277087 59113
rect 277121 59085 277149 59113
rect 277059 59023 277087 59051
rect 277121 59023 277149 59051
rect 277059 58961 277087 58989
rect 277121 58961 277149 58989
rect 269379 56147 269407 56175
rect 269441 56147 269469 56175
rect 269379 56085 269407 56113
rect 269441 56085 269469 56113
rect 269379 56023 269407 56051
rect 269441 56023 269469 56051
rect 269379 55961 269407 55989
rect 269441 55961 269469 55989
rect 279237 56147 279265 56175
rect 279299 56147 279327 56175
rect 279361 56147 279389 56175
rect 279423 56147 279451 56175
rect 279237 56085 279265 56113
rect 279299 56085 279327 56113
rect 279361 56085 279389 56113
rect 279423 56085 279451 56113
rect 279237 56023 279265 56051
rect 279299 56023 279327 56051
rect 279361 56023 279389 56051
rect 279423 56023 279451 56051
rect 279237 55961 279265 55989
rect 279299 55961 279327 55989
rect 279361 55961 279389 55989
rect 279423 55961 279451 55989
rect 265737 50147 265765 50175
rect 265799 50147 265827 50175
rect 265861 50147 265889 50175
rect 265923 50147 265951 50175
rect 265737 50085 265765 50113
rect 265799 50085 265827 50113
rect 265861 50085 265889 50113
rect 265923 50085 265951 50113
rect 265737 50023 265765 50051
rect 265799 50023 265827 50051
rect 265861 50023 265889 50051
rect 265923 50023 265951 50051
rect 265737 49961 265765 49989
rect 265799 49961 265827 49989
rect 265861 49961 265889 49989
rect 265923 49961 265951 49989
rect 277059 50147 277087 50175
rect 277121 50147 277149 50175
rect 277059 50085 277087 50113
rect 277121 50085 277149 50113
rect 277059 50023 277087 50051
rect 277121 50023 277149 50051
rect 277059 49961 277087 49989
rect 277121 49961 277149 49989
rect 269379 47147 269407 47175
rect 269441 47147 269469 47175
rect 269379 47085 269407 47113
rect 269441 47085 269469 47113
rect 269379 47023 269407 47051
rect 269441 47023 269469 47051
rect 269379 46961 269407 46989
rect 269441 46961 269469 46989
rect 279237 47147 279265 47175
rect 279299 47147 279327 47175
rect 279361 47147 279389 47175
rect 279423 47147 279451 47175
rect 279237 47085 279265 47113
rect 279299 47085 279327 47113
rect 279361 47085 279389 47113
rect 279423 47085 279451 47113
rect 279237 47023 279265 47051
rect 279299 47023 279327 47051
rect 279361 47023 279389 47051
rect 279423 47023 279451 47051
rect 279237 46961 279265 46989
rect 279299 46961 279327 46989
rect 279361 46961 279389 46989
rect 279423 46961 279451 46989
rect 265737 41147 265765 41175
rect 265799 41147 265827 41175
rect 265861 41147 265889 41175
rect 265923 41147 265951 41175
rect 265737 41085 265765 41113
rect 265799 41085 265827 41113
rect 265861 41085 265889 41113
rect 265923 41085 265951 41113
rect 265737 41023 265765 41051
rect 265799 41023 265827 41051
rect 265861 41023 265889 41051
rect 265923 41023 265951 41051
rect 265737 40961 265765 40989
rect 265799 40961 265827 40989
rect 265861 40961 265889 40989
rect 265923 40961 265951 40989
rect 277059 41147 277087 41175
rect 277121 41147 277149 41175
rect 277059 41085 277087 41113
rect 277121 41085 277149 41113
rect 277059 41023 277087 41051
rect 277121 41023 277149 41051
rect 277059 40961 277087 40989
rect 277121 40961 277149 40989
rect 269379 38147 269407 38175
rect 269441 38147 269469 38175
rect 269379 38085 269407 38113
rect 269441 38085 269469 38113
rect 269379 38023 269407 38051
rect 269441 38023 269469 38051
rect 269379 37961 269407 37989
rect 269441 37961 269469 37989
rect 279237 38147 279265 38175
rect 279299 38147 279327 38175
rect 279361 38147 279389 38175
rect 279423 38147 279451 38175
rect 279237 38085 279265 38113
rect 279299 38085 279327 38113
rect 279361 38085 279389 38113
rect 279423 38085 279451 38113
rect 279237 38023 279265 38051
rect 279299 38023 279327 38051
rect 279361 38023 279389 38051
rect 279423 38023 279451 38051
rect 279237 37961 279265 37989
rect 279299 37961 279327 37989
rect 279361 37961 279389 37989
rect 279423 37961 279451 37989
rect 265737 32147 265765 32175
rect 265799 32147 265827 32175
rect 265861 32147 265889 32175
rect 265923 32147 265951 32175
rect 265737 32085 265765 32113
rect 265799 32085 265827 32113
rect 265861 32085 265889 32113
rect 265923 32085 265951 32113
rect 265737 32023 265765 32051
rect 265799 32023 265827 32051
rect 265861 32023 265889 32051
rect 265923 32023 265951 32051
rect 265737 31961 265765 31989
rect 265799 31961 265827 31989
rect 265861 31961 265889 31989
rect 265923 31961 265951 31989
rect 277059 32147 277087 32175
rect 277121 32147 277149 32175
rect 277059 32085 277087 32113
rect 277121 32085 277149 32113
rect 277059 32023 277087 32051
rect 277121 32023 277149 32051
rect 277059 31961 277087 31989
rect 277121 31961 277149 31989
rect 269379 29147 269407 29175
rect 269441 29147 269469 29175
rect 269379 29085 269407 29113
rect 269441 29085 269469 29113
rect 269379 29023 269407 29051
rect 269441 29023 269469 29051
rect 269379 28961 269407 28989
rect 269441 28961 269469 28989
rect 279237 29147 279265 29175
rect 279299 29147 279327 29175
rect 279361 29147 279389 29175
rect 279423 29147 279451 29175
rect 279237 29085 279265 29113
rect 279299 29085 279327 29113
rect 279361 29085 279389 29113
rect 279423 29085 279451 29113
rect 279237 29023 279265 29051
rect 279299 29023 279327 29051
rect 279361 29023 279389 29051
rect 279423 29023 279451 29051
rect 279237 28961 279265 28989
rect 279299 28961 279327 28989
rect 279361 28961 279389 28989
rect 279423 28961 279451 28989
rect 265737 23147 265765 23175
rect 265799 23147 265827 23175
rect 265861 23147 265889 23175
rect 265923 23147 265951 23175
rect 265737 23085 265765 23113
rect 265799 23085 265827 23113
rect 265861 23085 265889 23113
rect 265923 23085 265951 23113
rect 265737 23023 265765 23051
rect 265799 23023 265827 23051
rect 265861 23023 265889 23051
rect 265923 23023 265951 23051
rect 265737 22961 265765 22989
rect 265799 22961 265827 22989
rect 265861 22961 265889 22989
rect 265923 22961 265951 22989
rect 277059 23147 277087 23175
rect 277121 23147 277149 23175
rect 277059 23085 277087 23113
rect 277121 23085 277149 23113
rect 277059 23023 277087 23051
rect 277121 23023 277149 23051
rect 277059 22961 277087 22989
rect 277121 22961 277149 22989
rect 269379 20147 269407 20175
rect 269441 20147 269469 20175
rect 269379 20085 269407 20113
rect 269441 20085 269469 20113
rect 269379 20023 269407 20051
rect 269441 20023 269469 20051
rect 269379 19961 269407 19989
rect 269441 19961 269469 19989
rect 279237 20147 279265 20175
rect 279299 20147 279327 20175
rect 279361 20147 279389 20175
rect 279423 20147 279451 20175
rect 279237 20085 279265 20113
rect 279299 20085 279327 20113
rect 279361 20085 279389 20113
rect 279423 20085 279451 20113
rect 279237 20023 279265 20051
rect 279299 20023 279327 20051
rect 279361 20023 279389 20051
rect 279423 20023 279451 20051
rect 279237 19961 279265 19989
rect 279299 19961 279327 19989
rect 279361 19961 279389 19989
rect 279423 19961 279451 19989
rect 265737 14147 265765 14175
rect 265799 14147 265827 14175
rect 265861 14147 265889 14175
rect 265923 14147 265951 14175
rect 265737 14085 265765 14113
rect 265799 14085 265827 14113
rect 265861 14085 265889 14113
rect 265923 14085 265951 14113
rect 265737 14023 265765 14051
rect 265799 14023 265827 14051
rect 265861 14023 265889 14051
rect 265923 14023 265951 14051
rect 265737 13961 265765 13989
rect 265799 13961 265827 13989
rect 265861 13961 265889 13989
rect 265923 13961 265951 13989
rect 277059 14147 277087 14175
rect 277121 14147 277149 14175
rect 277059 14085 277087 14113
rect 277121 14085 277149 14113
rect 277059 14023 277087 14051
rect 277121 14023 277149 14051
rect 277059 13961 277087 13989
rect 277121 13961 277149 13989
rect 269379 11147 269407 11175
rect 269441 11147 269469 11175
rect 269379 11085 269407 11113
rect 269441 11085 269469 11113
rect 269379 11023 269407 11051
rect 269441 11023 269469 11051
rect 269379 10961 269407 10989
rect 269441 10961 269469 10989
rect 279237 11147 279265 11175
rect 279299 11147 279327 11175
rect 279361 11147 279389 11175
rect 279423 11147 279451 11175
rect 279237 11085 279265 11113
rect 279299 11085 279327 11113
rect 279361 11085 279389 11113
rect 279423 11085 279451 11113
rect 279237 11023 279265 11051
rect 279299 11023 279327 11051
rect 279361 11023 279389 11051
rect 279423 11023 279451 11051
rect 279237 10961 279265 10989
rect 279299 10961 279327 10989
rect 279361 10961 279389 10989
rect 279423 10961 279451 10989
rect 265737 5147 265765 5175
rect 265799 5147 265827 5175
rect 265861 5147 265889 5175
rect 265923 5147 265951 5175
rect 265737 5085 265765 5113
rect 265799 5085 265827 5113
rect 265861 5085 265889 5113
rect 265923 5085 265951 5113
rect 265737 5023 265765 5051
rect 265799 5023 265827 5051
rect 265861 5023 265889 5051
rect 265923 5023 265951 5051
rect 265737 4961 265765 4989
rect 265799 4961 265827 4989
rect 265861 4961 265889 4989
rect 265923 4961 265951 4989
rect 277059 5147 277087 5175
rect 277121 5147 277149 5175
rect 277059 5085 277087 5113
rect 277121 5085 277149 5113
rect 277059 5023 277087 5051
rect 277121 5023 277149 5051
rect 277059 4961 277087 4989
rect 277121 4961 277149 4989
rect 265737 -588 265765 -560
rect 265799 -588 265827 -560
rect 265861 -588 265889 -560
rect 265923 -588 265951 -560
rect 265737 -650 265765 -622
rect 265799 -650 265827 -622
rect 265861 -650 265889 -622
rect 265923 -650 265951 -622
rect 265737 -712 265765 -684
rect 265799 -712 265827 -684
rect 265861 -712 265889 -684
rect 265923 -712 265951 -684
rect 265737 -774 265765 -746
rect 265799 -774 265827 -746
rect 265861 -774 265889 -746
rect 265923 -774 265951 -746
rect 279237 2147 279265 2175
rect 279299 2147 279327 2175
rect 279361 2147 279389 2175
rect 279423 2147 279451 2175
rect 279237 2085 279265 2113
rect 279299 2085 279327 2113
rect 279361 2085 279389 2113
rect 279423 2085 279451 2113
rect 279237 2023 279265 2051
rect 279299 2023 279327 2051
rect 279361 2023 279389 2051
rect 279423 2023 279451 2051
rect 279237 1961 279265 1989
rect 279299 1961 279327 1989
rect 279361 1961 279389 1989
rect 279423 1961 279451 1989
rect 279237 -108 279265 -80
rect 279299 -108 279327 -80
rect 279361 -108 279389 -80
rect 279423 -108 279451 -80
rect 279237 -170 279265 -142
rect 279299 -170 279327 -142
rect 279361 -170 279389 -142
rect 279423 -170 279451 -142
rect 279237 -232 279265 -204
rect 279299 -232 279327 -204
rect 279361 -232 279389 -204
rect 279423 -232 279451 -204
rect 279237 -294 279265 -266
rect 279299 -294 279327 -266
rect 279361 -294 279389 -266
rect 279423 -294 279451 -266
rect 281097 299058 281125 299086
rect 281159 299058 281187 299086
rect 281221 299058 281249 299086
rect 281283 299058 281311 299086
rect 281097 298996 281125 299024
rect 281159 298996 281187 299024
rect 281221 298996 281249 299024
rect 281283 298996 281311 299024
rect 281097 298934 281125 298962
rect 281159 298934 281187 298962
rect 281221 298934 281249 298962
rect 281283 298934 281311 298962
rect 281097 298872 281125 298900
rect 281159 298872 281187 298900
rect 281221 298872 281249 298900
rect 281283 298872 281311 298900
rect 281097 293147 281125 293175
rect 281159 293147 281187 293175
rect 281221 293147 281249 293175
rect 281283 293147 281311 293175
rect 281097 293085 281125 293113
rect 281159 293085 281187 293113
rect 281221 293085 281249 293113
rect 281283 293085 281311 293113
rect 281097 293023 281125 293051
rect 281159 293023 281187 293051
rect 281221 293023 281249 293051
rect 281283 293023 281311 293051
rect 281097 292961 281125 292989
rect 281159 292961 281187 292989
rect 281221 292961 281249 292989
rect 281283 292961 281311 292989
rect 281097 284147 281125 284175
rect 281159 284147 281187 284175
rect 281221 284147 281249 284175
rect 281283 284147 281311 284175
rect 281097 284085 281125 284113
rect 281159 284085 281187 284113
rect 281221 284085 281249 284113
rect 281283 284085 281311 284113
rect 281097 284023 281125 284051
rect 281159 284023 281187 284051
rect 281221 284023 281249 284051
rect 281283 284023 281311 284051
rect 281097 283961 281125 283989
rect 281159 283961 281187 283989
rect 281221 283961 281249 283989
rect 281283 283961 281311 283989
rect 281097 275147 281125 275175
rect 281159 275147 281187 275175
rect 281221 275147 281249 275175
rect 281283 275147 281311 275175
rect 281097 275085 281125 275113
rect 281159 275085 281187 275113
rect 281221 275085 281249 275113
rect 281283 275085 281311 275113
rect 281097 275023 281125 275051
rect 281159 275023 281187 275051
rect 281221 275023 281249 275051
rect 281283 275023 281311 275051
rect 281097 274961 281125 274989
rect 281159 274961 281187 274989
rect 281221 274961 281249 274989
rect 281283 274961 281311 274989
rect 281097 266147 281125 266175
rect 281159 266147 281187 266175
rect 281221 266147 281249 266175
rect 281283 266147 281311 266175
rect 281097 266085 281125 266113
rect 281159 266085 281187 266113
rect 281221 266085 281249 266113
rect 281283 266085 281311 266113
rect 281097 266023 281125 266051
rect 281159 266023 281187 266051
rect 281221 266023 281249 266051
rect 281283 266023 281311 266051
rect 281097 265961 281125 265989
rect 281159 265961 281187 265989
rect 281221 265961 281249 265989
rect 281283 265961 281311 265989
rect 281097 257147 281125 257175
rect 281159 257147 281187 257175
rect 281221 257147 281249 257175
rect 281283 257147 281311 257175
rect 281097 257085 281125 257113
rect 281159 257085 281187 257113
rect 281221 257085 281249 257113
rect 281283 257085 281311 257113
rect 281097 257023 281125 257051
rect 281159 257023 281187 257051
rect 281221 257023 281249 257051
rect 281283 257023 281311 257051
rect 281097 256961 281125 256989
rect 281159 256961 281187 256989
rect 281221 256961 281249 256989
rect 281283 256961 281311 256989
rect 281097 248147 281125 248175
rect 281159 248147 281187 248175
rect 281221 248147 281249 248175
rect 281283 248147 281311 248175
rect 281097 248085 281125 248113
rect 281159 248085 281187 248113
rect 281221 248085 281249 248113
rect 281283 248085 281311 248113
rect 281097 248023 281125 248051
rect 281159 248023 281187 248051
rect 281221 248023 281249 248051
rect 281283 248023 281311 248051
rect 281097 247961 281125 247989
rect 281159 247961 281187 247989
rect 281221 247961 281249 247989
rect 281283 247961 281311 247989
rect 281097 239147 281125 239175
rect 281159 239147 281187 239175
rect 281221 239147 281249 239175
rect 281283 239147 281311 239175
rect 281097 239085 281125 239113
rect 281159 239085 281187 239113
rect 281221 239085 281249 239113
rect 281283 239085 281311 239113
rect 281097 239023 281125 239051
rect 281159 239023 281187 239051
rect 281221 239023 281249 239051
rect 281283 239023 281311 239051
rect 281097 238961 281125 238989
rect 281159 238961 281187 238989
rect 281221 238961 281249 238989
rect 281283 238961 281311 238989
rect 281097 230147 281125 230175
rect 281159 230147 281187 230175
rect 281221 230147 281249 230175
rect 281283 230147 281311 230175
rect 281097 230085 281125 230113
rect 281159 230085 281187 230113
rect 281221 230085 281249 230113
rect 281283 230085 281311 230113
rect 281097 230023 281125 230051
rect 281159 230023 281187 230051
rect 281221 230023 281249 230051
rect 281283 230023 281311 230051
rect 281097 229961 281125 229989
rect 281159 229961 281187 229989
rect 281221 229961 281249 229989
rect 281283 229961 281311 229989
rect 281097 221147 281125 221175
rect 281159 221147 281187 221175
rect 281221 221147 281249 221175
rect 281283 221147 281311 221175
rect 281097 221085 281125 221113
rect 281159 221085 281187 221113
rect 281221 221085 281249 221113
rect 281283 221085 281311 221113
rect 281097 221023 281125 221051
rect 281159 221023 281187 221051
rect 281221 221023 281249 221051
rect 281283 221023 281311 221051
rect 281097 220961 281125 220989
rect 281159 220961 281187 220989
rect 281221 220961 281249 220989
rect 281283 220961 281311 220989
rect 281097 212147 281125 212175
rect 281159 212147 281187 212175
rect 281221 212147 281249 212175
rect 281283 212147 281311 212175
rect 281097 212085 281125 212113
rect 281159 212085 281187 212113
rect 281221 212085 281249 212113
rect 281283 212085 281311 212113
rect 281097 212023 281125 212051
rect 281159 212023 281187 212051
rect 281221 212023 281249 212051
rect 281283 212023 281311 212051
rect 281097 211961 281125 211989
rect 281159 211961 281187 211989
rect 281221 211961 281249 211989
rect 281283 211961 281311 211989
rect 281097 203147 281125 203175
rect 281159 203147 281187 203175
rect 281221 203147 281249 203175
rect 281283 203147 281311 203175
rect 281097 203085 281125 203113
rect 281159 203085 281187 203113
rect 281221 203085 281249 203113
rect 281283 203085 281311 203113
rect 281097 203023 281125 203051
rect 281159 203023 281187 203051
rect 281221 203023 281249 203051
rect 281283 203023 281311 203051
rect 281097 202961 281125 202989
rect 281159 202961 281187 202989
rect 281221 202961 281249 202989
rect 281283 202961 281311 202989
rect 281097 194147 281125 194175
rect 281159 194147 281187 194175
rect 281221 194147 281249 194175
rect 281283 194147 281311 194175
rect 281097 194085 281125 194113
rect 281159 194085 281187 194113
rect 281221 194085 281249 194113
rect 281283 194085 281311 194113
rect 281097 194023 281125 194051
rect 281159 194023 281187 194051
rect 281221 194023 281249 194051
rect 281283 194023 281311 194051
rect 281097 193961 281125 193989
rect 281159 193961 281187 193989
rect 281221 193961 281249 193989
rect 281283 193961 281311 193989
rect 281097 185147 281125 185175
rect 281159 185147 281187 185175
rect 281221 185147 281249 185175
rect 281283 185147 281311 185175
rect 281097 185085 281125 185113
rect 281159 185085 281187 185113
rect 281221 185085 281249 185113
rect 281283 185085 281311 185113
rect 281097 185023 281125 185051
rect 281159 185023 281187 185051
rect 281221 185023 281249 185051
rect 281283 185023 281311 185051
rect 281097 184961 281125 184989
rect 281159 184961 281187 184989
rect 281221 184961 281249 184989
rect 281283 184961 281311 184989
rect 281097 176147 281125 176175
rect 281159 176147 281187 176175
rect 281221 176147 281249 176175
rect 281283 176147 281311 176175
rect 281097 176085 281125 176113
rect 281159 176085 281187 176113
rect 281221 176085 281249 176113
rect 281283 176085 281311 176113
rect 281097 176023 281125 176051
rect 281159 176023 281187 176051
rect 281221 176023 281249 176051
rect 281283 176023 281311 176051
rect 281097 175961 281125 175989
rect 281159 175961 281187 175989
rect 281221 175961 281249 175989
rect 281283 175961 281311 175989
rect 294597 298578 294625 298606
rect 294659 298578 294687 298606
rect 294721 298578 294749 298606
rect 294783 298578 294811 298606
rect 294597 298516 294625 298544
rect 294659 298516 294687 298544
rect 294721 298516 294749 298544
rect 294783 298516 294811 298544
rect 294597 298454 294625 298482
rect 294659 298454 294687 298482
rect 294721 298454 294749 298482
rect 294783 298454 294811 298482
rect 294597 298392 294625 298420
rect 294659 298392 294687 298420
rect 294721 298392 294749 298420
rect 294783 298392 294811 298420
rect 294597 290147 294625 290175
rect 294659 290147 294687 290175
rect 294721 290147 294749 290175
rect 294783 290147 294811 290175
rect 294597 290085 294625 290113
rect 294659 290085 294687 290113
rect 294721 290085 294749 290113
rect 294783 290085 294811 290113
rect 294597 290023 294625 290051
rect 294659 290023 294687 290051
rect 294721 290023 294749 290051
rect 294783 290023 294811 290051
rect 294597 289961 294625 289989
rect 294659 289961 294687 289989
rect 294721 289961 294749 289989
rect 294783 289961 294811 289989
rect 294597 281147 294625 281175
rect 294659 281147 294687 281175
rect 294721 281147 294749 281175
rect 294783 281147 294811 281175
rect 294597 281085 294625 281113
rect 294659 281085 294687 281113
rect 294721 281085 294749 281113
rect 294783 281085 294811 281113
rect 294597 281023 294625 281051
rect 294659 281023 294687 281051
rect 294721 281023 294749 281051
rect 294783 281023 294811 281051
rect 294597 280961 294625 280989
rect 294659 280961 294687 280989
rect 294721 280961 294749 280989
rect 294783 280961 294811 280989
rect 294597 272147 294625 272175
rect 294659 272147 294687 272175
rect 294721 272147 294749 272175
rect 294783 272147 294811 272175
rect 294597 272085 294625 272113
rect 294659 272085 294687 272113
rect 294721 272085 294749 272113
rect 294783 272085 294811 272113
rect 294597 272023 294625 272051
rect 294659 272023 294687 272051
rect 294721 272023 294749 272051
rect 294783 272023 294811 272051
rect 294597 271961 294625 271989
rect 294659 271961 294687 271989
rect 294721 271961 294749 271989
rect 294783 271961 294811 271989
rect 294597 263147 294625 263175
rect 294659 263147 294687 263175
rect 294721 263147 294749 263175
rect 294783 263147 294811 263175
rect 294597 263085 294625 263113
rect 294659 263085 294687 263113
rect 294721 263085 294749 263113
rect 294783 263085 294811 263113
rect 294597 263023 294625 263051
rect 294659 263023 294687 263051
rect 294721 263023 294749 263051
rect 294783 263023 294811 263051
rect 294597 262961 294625 262989
rect 294659 262961 294687 262989
rect 294721 262961 294749 262989
rect 294783 262961 294811 262989
rect 294597 254147 294625 254175
rect 294659 254147 294687 254175
rect 294721 254147 294749 254175
rect 294783 254147 294811 254175
rect 294597 254085 294625 254113
rect 294659 254085 294687 254113
rect 294721 254085 294749 254113
rect 294783 254085 294811 254113
rect 294597 254023 294625 254051
rect 294659 254023 294687 254051
rect 294721 254023 294749 254051
rect 294783 254023 294811 254051
rect 294597 253961 294625 253989
rect 294659 253961 294687 253989
rect 294721 253961 294749 253989
rect 294783 253961 294811 253989
rect 294597 245147 294625 245175
rect 294659 245147 294687 245175
rect 294721 245147 294749 245175
rect 294783 245147 294811 245175
rect 294597 245085 294625 245113
rect 294659 245085 294687 245113
rect 294721 245085 294749 245113
rect 294783 245085 294811 245113
rect 294597 245023 294625 245051
rect 294659 245023 294687 245051
rect 294721 245023 294749 245051
rect 294783 245023 294811 245051
rect 294597 244961 294625 244989
rect 294659 244961 294687 244989
rect 294721 244961 294749 244989
rect 294783 244961 294811 244989
rect 294597 236147 294625 236175
rect 294659 236147 294687 236175
rect 294721 236147 294749 236175
rect 294783 236147 294811 236175
rect 294597 236085 294625 236113
rect 294659 236085 294687 236113
rect 294721 236085 294749 236113
rect 294783 236085 294811 236113
rect 294597 236023 294625 236051
rect 294659 236023 294687 236051
rect 294721 236023 294749 236051
rect 294783 236023 294811 236051
rect 294597 235961 294625 235989
rect 294659 235961 294687 235989
rect 294721 235961 294749 235989
rect 294783 235961 294811 235989
rect 294597 227147 294625 227175
rect 294659 227147 294687 227175
rect 294721 227147 294749 227175
rect 294783 227147 294811 227175
rect 294597 227085 294625 227113
rect 294659 227085 294687 227113
rect 294721 227085 294749 227113
rect 294783 227085 294811 227113
rect 294597 227023 294625 227051
rect 294659 227023 294687 227051
rect 294721 227023 294749 227051
rect 294783 227023 294811 227051
rect 294597 226961 294625 226989
rect 294659 226961 294687 226989
rect 294721 226961 294749 226989
rect 294783 226961 294811 226989
rect 294597 218147 294625 218175
rect 294659 218147 294687 218175
rect 294721 218147 294749 218175
rect 294783 218147 294811 218175
rect 294597 218085 294625 218113
rect 294659 218085 294687 218113
rect 294721 218085 294749 218113
rect 294783 218085 294811 218113
rect 294597 218023 294625 218051
rect 294659 218023 294687 218051
rect 294721 218023 294749 218051
rect 294783 218023 294811 218051
rect 294597 217961 294625 217989
rect 294659 217961 294687 217989
rect 294721 217961 294749 217989
rect 294783 217961 294811 217989
rect 294597 209147 294625 209175
rect 294659 209147 294687 209175
rect 294721 209147 294749 209175
rect 294783 209147 294811 209175
rect 294597 209085 294625 209113
rect 294659 209085 294687 209113
rect 294721 209085 294749 209113
rect 294783 209085 294811 209113
rect 294597 209023 294625 209051
rect 294659 209023 294687 209051
rect 294721 209023 294749 209051
rect 294783 209023 294811 209051
rect 294597 208961 294625 208989
rect 294659 208961 294687 208989
rect 294721 208961 294749 208989
rect 294783 208961 294811 208989
rect 294597 200147 294625 200175
rect 294659 200147 294687 200175
rect 294721 200147 294749 200175
rect 294783 200147 294811 200175
rect 294597 200085 294625 200113
rect 294659 200085 294687 200113
rect 294721 200085 294749 200113
rect 294783 200085 294811 200113
rect 294597 200023 294625 200051
rect 294659 200023 294687 200051
rect 294721 200023 294749 200051
rect 294783 200023 294811 200051
rect 294597 199961 294625 199989
rect 294659 199961 294687 199989
rect 294721 199961 294749 199989
rect 294783 199961 294811 199989
rect 294597 191147 294625 191175
rect 294659 191147 294687 191175
rect 294721 191147 294749 191175
rect 294783 191147 294811 191175
rect 294597 191085 294625 191113
rect 294659 191085 294687 191113
rect 294721 191085 294749 191113
rect 294783 191085 294811 191113
rect 294597 191023 294625 191051
rect 294659 191023 294687 191051
rect 294721 191023 294749 191051
rect 294783 191023 294811 191051
rect 294597 190961 294625 190989
rect 294659 190961 294687 190989
rect 294721 190961 294749 190989
rect 294783 190961 294811 190989
rect 294597 182147 294625 182175
rect 294659 182147 294687 182175
rect 294721 182147 294749 182175
rect 294783 182147 294811 182175
rect 294597 182085 294625 182113
rect 294659 182085 294687 182113
rect 294721 182085 294749 182113
rect 294783 182085 294811 182113
rect 294597 182023 294625 182051
rect 294659 182023 294687 182051
rect 294721 182023 294749 182051
rect 294783 182023 294811 182051
rect 294597 181961 294625 181989
rect 294659 181961 294687 181989
rect 294721 181961 294749 181989
rect 294783 181961 294811 181989
rect 284739 173147 284767 173175
rect 284801 173147 284829 173175
rect 284739 173085 284767 173113
rect 284801 173085 284829 173113
rect 284739 173023 284767 173051
rect 284801 173023 284829 173051
rect 284739 172961 284767 172989
rect 284801 172961 284829 172989
rect 281097 167147 281125 167175
rect 281159 167147 281187 167175
rect 281221 167147 281249 167175
rect 281283 167147 281311 167175
rect 281097 167085 281125 167113
rect 281159 167085 281187 167113
rect 281221 167085 281249 167113
rect 281283 167085 281311 167113
rect 281097 167023 281125 167051
rect 281159 167023 281187 167051
rect 281221 167023 281249 167051
rect 281283 167023 281311 167051
rect 281097 166961 281125 166989
rect 281159 166961 281187 166989
rect 281221 166961 281249 166989
rect 281283 166961 281311 166989
rect 284739 164147 284767 164175
rect 284801 164147 284829 164175
rect 284739 164085 284767 164113
rect 284801 164085 284829 164113
rect 284739 164023 284767 164051
rect 284801 164023 284829 164051
rect 284739 163961 284767 163989
rect 284801 163961 284829 163989
rect 281097 158147 281125 158175
rect 281159 158147 281187 158175
rect 281221 158147 281249 158175
rect 281283 158147 281311 158175
rect 281097 158085 281125 158113
rect 281159 158085 281187 158113
rect 281221 158085 281249 158113
rect 281283 158085 281311 158113
rect 281097 158023 281125 158051
rect 281159 158023 281187 158051
rect 281221 158023 281249 158051
rect 281283 158023 281311 158051
rect 281097 157961 281125 157989
rect 281159 157961 281187 157989
rect 281221 157961 281249 157989
rect 281283 157961 281311 157989
rect 294597 173147 294625 173175
rect 294659 173147 294687 173175
rect 294721 173147 294749 173175
rect 294783 173147 294811 173175
rect 294597 173085 294625 173113
rect 294659 173085 294687 173113
rect 294721 173085 294749 173113
rect 294783 173085 294811 173113
rect 294597 173023 294625 173051
rect 294659 173023 294687 173051
rect 294721 173023 294749 173051
rect 294783 173023 294811 173051
rect 294597 172961 294625 172989
rect 294659 172961 294687 172989
rect 294721 172961 294749 172989
rect 294783 172961 294811 172989
rect 284739 155147 284767 155175
rect 284801 155147 284829 155175
rect 284739 155085 284767 155113
rect 284801 155085 284829 155113
rect 284739 155023 284767 155051
rect 284801 155023 284829 155051
rect 284739 154961 284767 154989
rect 284801 154961 284829 154989
rect 281097 149147 281125 149175
rect 281159 149147 281187 149175
rect 281221 149147 281249 149175
rect 281283 149147 281311 149175
rect 281097 149085 281125 149113
rect 281159 149085 281187 149113
rect 281221 149085 281249 149113
rect 281283 149085 281311 149113
rect 281097 149023 281125 149051
rect 281159 149023 281187 149051
rect 281221 149023 281249 149051
rect 281283 149023 281311 149051
rect 281097 148961 281125 148989
rect 281159 148961 281187 148989
rect 281221 148961 281249 148989
rect 281283 148961 281311 148989
rect 284739 146147 284767 146175
rect 284801 146147 284829 146175
rect 284739 146085 284767 146113
rect 284801 146085 284829 146113
rect 284739 146023 284767 146051
rect 284801 146023 284829 146051
rect 284739 145961 284767 145989
rect 284801 145961 284829 145989
rect 281097 140147 281125 140175
rect 281159 140147 281187 140175
rect 281221 140147 281249 140175
rect 281283 140147 281311 140175
rect 281097 140085 281125 140113
rect 281159 140085 281187 140113
rect 281221 140085 281249 140113
rect 281283 140085 281311 140113
rect 281097 140023 281125 140051
rect 281159 140023 281187 140051
rect 281221 140023 281249 140051
rect 281283 140023 281311 140051
rect 281097 139961 281125 139989
rect 281159 139961 281187 139989
rect 281221 139961 281249 139989
rect 281283 139961 281311 139989
rect 284739 137147 284767 137175
rect 284801 137147 284829 137175
rect 284739 137085 284767 137113
rect 284801 137085 284829 137113
rect 284739 137023 284767 137051
rect 284801 137023 284829 137051
rect 284739 136961 284767 136989
rect 284801 136961 284829 136989
rect 294597 164147 294625 164175
rect 294659 164147 294687 164175
rect 294721 164147 294749 164175
rect 294783 164147 294811 164175
rect 294597 164085 294625 164113
rect 294659 164085 294687 164113
rect 294721 164085 294749 164113
rect 294783 164085 294811 164113
rect 294597 164023 294625 164051
rect 294659 164023 294687 164051
rect 294721 164023 294749 164051
rect 294783 164023 294811 164051
rect 294597 163961 294625 163989
rect 294659 163961 294687 163989
rect 294721 163961 294749 163989
rect 294783 163961 294811 163989
rect 281097 131147 281125 131175
rect 281159 131147 281187 131175
rect 281221 131147 281249 131175
rect 281283 131147 281311 131175
rect 281097 131085 281125 131113
rect 281159 131085 281187 131113
rect 281221 131085 281249 131113
rect 281283 131085 281311 131113
rect 281097 131023 281125 131051
rect 281159 131023 281187 131051
rect 281221 131023 281249 131051
rect 281283 131023 281311 131051
rect 281097 130961 281125 130989
rect 281159 130961 281187 130989
rect 281221 130961 281249 130989
rect 281283 130961 281311 130989
rect 284739 128147 284767 128175
rect 284801 128147 284829 128175
rect 284739 128085 284767 128113
rect 284801 128085 284829 128113
rect 284739 128023 284767 128051
rect 284801 128023 284829 128051
rect 284739 127961 284767 127989
rect 284801 127961 284829 127989
rect 281097 122147 281125 122175
rect 281159 122147 281187 122175
rect 281221 122147 281249 122175
rect 281283 122147 281311 122175
rect 281097 122085 281125 122113
rect 281159 122085 281187 122113
rect 281221 122085 281249 122113
rect 281283 122085 281311 122113
rect 281097 122023 281125 122051
rect 281159 122023 281187 122051
rect 281221 122023 281249 122051
rect 281283 122023 281311 122051
rect 281097 121961 281125 121989
rect 281159 121961 281187 121989
rect 281221 121961 281249 121989
rect 281283 121961 281311 121989
rect 284739 119147 284767 119175
rect 284801 119147 284829 119175
rect 284739 119085 284767 119113
rect 284801 119085 284829 119113
rect 284739 119023 284767 119051
rect 284801 119023 284829 119051
rect 284739 118961 284767 118989
rect 284801 118961 284829 118989
rect 294597 155147 294625 155175
rect 294659 155147 294687 155175
rect 294721 155147 294749 155175
rect 294783 155147 294811 155175
rect 294597 155085 294625 155113
rect 294659 155085 294687 155113
rect 294721 155085 294749 155113
rect 294783 155085 294811 155113
rect 294597 155023 294625 155051
rect 294659 155023 294687 155051
rect 294721 155023 294749 155051
rect 294783 155023 294811 155051
rect 294597 154961 294625 154989
rect 294659 154961 294687 154989
rect 294721 154961 294749 154989
rect 294783 154961 294811 154989
rect 294597 146147 294625 146175
rect 294659 146147 294687 146175
rect 294721 146147 294749 146175
rect 294783 146147 294811 146175
rect 294597 146085 294625 146113
rect 294659 146085 294687 146113
rect 294721 146085 294749 146113
rect 294783 146085 294811 146113
rect 294597 146023 294625 146051
rect 294659 146023 294687 146051
rect 294721 146023 294749 146051
rect 294783 146023 294811 146051
rect 294597 145961 294625 145989
rect 294659 145961 294687 145989
rect 294721 145961 294749 145989
rect 294783 145961 294811 145989
rect 294597 137147 294625 137175
rect 294659 137147 294687 137175
rect 294721 137147 294749 137175
rect 294783 137147 294811 137175
rect 294597 137085 294625 137113
rect 294659 137085 294687 137113
rect 294721 137085 294749 137113
rect 294783 137085 294811 137113
rect 294597 137023 294625 137051
rect 294659 137023 294687 137051
rect 294721 137023 294749 137051
rect 294783 137023 294811 137051
rect 294597 136961 294625 136989
rect 294659 136961 294687 136989
rect 294721 136961 294749 136989
rect 294783 136961 294811 136989
rect 294597 128147 294625 128175
rect 294659 128147 294687 128175
rect 294721 128147 294749 128175
rect 294783 128147 294811 128175
rect 294597 128085 294625 128113
rect 294659 128085 294687 128113
rect 294721 128085 294749 128113
rect 294783 128085 294811 128113
rect 294597 128023 294625 128051
rect 294659 128023 294687 128051
rect 294721 128023 294749 128051
rect 294783 128023 294811 128051
rect 294597 127961 294625 127989
rect 294659 127961 294687 127989
rect 294721 127961 294749 127989
rect 294783 127961 294811 127989
rect 281097 113147 281125 113175
rect 281159 113147 281187 113175
rect 281221 113147 281249 113175
rect 281283 113147 281311 113175
rect 281097 113085 281125 113113
rect 281159 113085 281187 113113
rect 281221 113085 281249 113113
rect 281283 113085 281311 113113
rect 281097 113023 281125 113051
rect 281159 113023 281187 113051
rect 281221 113023 281249 113051
rect 281283 113023 281311 113051
rect 281097 112961 281125 112989
rect 281159 112961 281187 112989
rect 281221 112961 281249 112989
rect 281283 112961 281311 112989
rect 284739 110147 284767 110175
rect 284801 110147 284829 110175
rect 284739 110085 284767 110113
rect 284801 110085 284829 110113
rect 284739 110023 284767 110051
rect 284801 110023 284829 110051
rect 284739 109961 284767 109989
rect 284801 109961 284829 109989
rect 281097 104147 281125 104175
rect 281159 104147 281187 104175
rect 281221 104147 281249 104175
rect 281283 104147 281311 104175
rect 281097 104085 281125 104113
rect 281159 104085 281187 104113
rect 281221 104085 281249 104113
rect 281283 104085 281311 104113
rect 281097 104023 281125 104051
rect 281159 104023 281187 104051
rect 281221 104023 281249 104051
rect 281283 104023 281311 104051
rect 281097 103961 281125 103989
rect 281159 103961 281187 103989
rect 281221 103961 281249 103989
rect 281283 103961 281311 103989
rect 284739 101147 284767 101175
rect 284801 101147 284829 101175
rect 284739 101085 284767 101113
rect 284801 101085 284829 101113
rect 284739 101023 284767 101051
rect 284801 101023 284829 101051
rect 284739 100961 284767 100989
rect 284801 100961 284829 100989
rect 294597 119147 294625 119175
rect 294659 119147 294687 119175
rect 294721 119147 294749 119175
rect 294783 119147 294811 119175
rect 294597 119085 294625 119113
rect 294659 119085 294687 119113
rect 294721 119085 294749 119113
rect 294783 119085 294811 119113
rect 294597 119023 294625 119051
rect 294659 119023 294687 119051
rect 294721 119023 294749 119051
rect 294783 119023 294811 119051
rect 294597 118961 294625 118989
rect 294659 118961 294687 118989
rect 294721 118961 294749 118989
rect 294783 118961 294811 118989
rect 294597 110147 294625 110175
rect 294659 110147 294687 110175
rect 294721 110147 294749 110175
rect 294783 110147 294811 110175
rect 294597 110085 294625 110113
rect 294659 110085 294687 110113
rect 294721 110085 294749 110113
rect 294783 110085 294811 110113
rect 294597 110023 294625 110051
rect 294659 110023 294687 110051
rect 294721 110023 294749 110051
rect 294783 110023 294811 110051
rect 294597 109961 294625 109989
rect 294659 109961 294687 109989
rect 294721 109961 294749 109989
rect 294783 109961 294811 109989
rect 294597 101147 294625 101175
rect 294659 101147 294687 101175
rect 294721 101147 294749 101175
rect 294783 101147 294811 101175
rect 294597 101085 294625 101113
rect 294659 101085 294687 101113
rect 294721 101085 294749 101113
rect 294783 101085 294811 101113
rect 294597 101023 294625 101051
rect 294659 101023 294687 101051
rect 294721 101023 294749 101051
rect 294783 101023 294811 101051
rect 294597 100961 294625 100989
rect 294659 100961 294687 100989
rect 294721 100961 294749 100989
rect 294783 100961 294811 100989
rect 281097 95147 281125 95175
rect 281159 95147 281187 95175
rect 281221 95147 281249 95175
rect 281283 95147 281311 95175
rect 281097 95085 281125 95113
rect 281159 95085 281187 95113
rect 281221 95085 281249 95113
rect 281283 95085 281311 95113
rect 281097 95023 281125 95051
rect 281159 95023 281187 95051
rect 281221 95023 281249 95051
rect 281283 95023 281311 95051
rect 281097 94961 281125 94989
rect 281159 94961 281187 94989
rect 281221 94961 281249 94989
rect 281283 94961 281311 94989
rect 284739 92147 284767 92175
rect 284801 92147 284829 92175
rect 284739 92085 284767 92113
rect 284801 92085 284829 92113
rect 284739 92023 284767 92051
rect 284801 92023 284829 92051
rect 284739 91961 284767 91989
rect 284801 91961 284829 91989
rect 281097 86147 281125 86175
rect 281159 86147 281187 86175
rect 281221 86147 281249 86175
rect 281283 86147 281311 86175
rect 281097 86085 281125 86113
rect 281159 86085 281187 86113
rect 281221 86085 281249 86113
rect 281283 86085 281311 86113
rect 281097 86023 281125 86051
rect 281159 86023 281187 86051
rect 281221 86023 281249 86051
rect 281283 86023 281311 86051
rect 281097 85961 281125 85989
rect 281159 85961 281187 85989
rect 281221 85961 281249 85989
rect 281283 85961 281311 85989
rect 284739 83147 284767 83175
rect 284801 83147 284829 83175
rect 284739 83085 284767 83113
rect 284801 83085 284829 83113
rect 284739 83023 284767 83051
rect 284801 83023 284829 83051
rect 284739 82961 284767 82989
rect 284801 82961 284829 82989
rect 281097 77147 281125 77175
rect 281159 77147 281187 77175
rect 281221 77147 281249 77175
rect 281283 77147 281311 77175
rect 281097 77085 281125 77113
rect 281159 77085 281187 77113
rect 281221 77085 281249 77113
rect 281283 77085 281311 77113
rect 281097 77023 281125 77051
rect 281159 77023 281187 77051
rect 281221 77023 281249 77051
rect 281283 77023 281311 77051
rect 281097 76961 281125 76989
rect 281159 76961 281187 76989
rect 281221 76961 281249 76989
rect 281283 76961 281311 76989
rect 294597 92147 294625 92175
rect 294659 92147 294687 92175
rect 294721 92147 294749 92175
rect 294783 92147 294811 92175
rect 294597 92085 294625 92113
rect 294659 92085 294687 92113
rect 294721 92085 294749 92113
rect 294783 92085 294811 92113
rect 294597 92023 294625 92051
rect 294659 92023 294687 92051
rect 294721 92023 294749 92051
rect 294783 92023 294811 92051
rect 294597 91961 294625 91989
rect 294659 91961 294687 91989
rect 294721 91961 294749 91989
rect 294783 91961 294811 91989
rect 294597 83147 294625 83175
rect 294659 83147 294687 83175
rect 294721 83147 294749 83175
rect 294783 83147 294811 83175
rect 294597 83085 294625 83113
rect 294659 83085 294687 83113
rect 294721 83085 294749 83113
rect 294783 83085 294811 83113
rect 294597 83023 294625 83051
rect 294659 83023 294687 83051
rect 294721 83023 294749 83051
rect 294783 83023 294811 83051
rect 294597 82961 294625 82989
rect 294659 82961 294687 82989
rect 294721 82961 294749 82989
rect 294783 82961 294811 82989
rect 284739 74147 284767 74175
rect 284801 74147 284829 74175
rect 284739 74085 284767 74113
rect 284801 74085 284829 74113
rect 284739 74023 284767 74051
rect 284801 74023 284829 74051
rect 284739 73961 284767 73989
rect 284801 73961 284829 73989
rect 294597 74147 294625 74175
rect 294659 74147 294687 74175
rect 294721 74147 294749 74175
rect 294783 74147 294811 74175
rect 294597 74085 294625 74113
rect 294659 74085 294687 74113
rect 294721 74085 294749 74113
rect 294783 74085 294811 74113
rect 294597 74023 294625 74051
rect 294659 74023 294687 74051
rect 294721 74023 294749 74051
rect 294783 74023 294811 74051
rect 294597 73961 294625 73989
rect 294659 73961 294687 73989
rect 294721 73961 294749 73989
rect 294783 73961 294811 73989
rect 281097 68147 281125 68175
rect 281159 68147 281187 68175
rect 281221 68147 281249 68175
rect 281283 68147 281311 68175
rect 281097 68085 281125 68113
rect 281159 68085 281187 68113
rect 281221 68085 281249 68113
rect 281283 68085 281311 68113
rect 281097 68023 281125 68051
rect 281159 68023 281187 68051
rect 281221 68023 281249 68051
rect 281283 68023 281311 68051
rect 281097 67961 281125 67989
rect 281159 67961 281187 67989
rect 281221 67961 281249 67989
rect 281283 67961 281311 67989
rect 284739 65147 284767 65175
rect 284801 65147 284829 65175
rect 284739 65085 284767 65113
rect 284801 65085 284829 65113
rect 284739 65023 284767 65051
rect 284801 65023 284829 65051
rect 284739 64961 284767 64989
rect 284801 64961 284829 64989
rect 281097 59147 281125 59175
rect 281159 59147 281187 59175
rect 281221 59147 281249 59175
rect 281283 59147 281311 59175
rect 281097 59085 281125 59113
rect 281159 59085 281187 59113
rect 281221 59085 281249 59113
rect 281283 59085 281311 59113
rect 281097 59023 281125 59051
rect 281159 59023 281187 59051
rect 281221 59023 281249 59051
rect 281283 59023 281311 59051
rect 281097 58961 281125 58989
rect 281159 58961 281187 58989
rect 281221 58961 281249 58989
rect 281283 58961 281311 58989
rect 294597 65147 294625 65175
rect 294659 65147 294687 65175
rect 294721 65147 294749 65175
rect 294783 65147 294811 65175
rect 294597 65085 294625 65113
rect 294659 65085 294687 65113
rect 294721 65085 294749 65113
rect 294783 65085 294811 65113
rect 294597 65023 294625 65051
rect 294659 65023 294687 65051
rect 294721 65023 294749 65051
rect 294783 65023 294811 65051
rect 294597 64961 294625 64989
rect 294659 64961 294687 64989
rect 294721 64961 294749 64989
rect 294783 64961 294811 64989
rect 284739 56147 284767 56175
rect 284801 56147 284829 56175
rect 284739 56085 284767 56113
rect 284801 56085 284829 56113
rect 284739 56023 284767 56051
rect 284801 56023 284829 56051
rect 284739 55961 284767 55989
rect 284801 55961 284829 55989
rect 296457 299058 296485 299086
rect 296519 299058 296547 299086
rect 296581 299058 296609 299086
rect 296643 299058 296671 299086
rect 296457 298996 296485 299024
rect 296519 298996 296547 299024
rect 296581 298996 296609 299024
rect 296643 298996 296671 299024
rect 296457 298934 296485 298962
rect 296519 298934 296547 298962
rect 296581 298934 296609 298962
rect 296643 298934 296671 298962
rect 296457 298872 296485 298900
rect 296519 298872 296547 298900
rect 296581 298872 296609 298900
rect 296643 298872 296671 298900
rect 298728 299058 298756 299086
rect 298790 299058 298818 299086
rect 298852 299058 298880 299086
rect 298914 299058 298942 299086
rect 298728 298996 298756 299024
rect 298790 298996 298818 299024
rect 298852 298996 298880 299024
rect 298914 298996 298942 299024
rect 298728 298934 298756 298962
rect 298790 298934 298818 298962
rect 298852 298934 298880 298962
rect 298914 298934 298942 298962
rect 298728 298872 298756 298900
rect 298790 298872 298818 298900
rect 298852 298872 298880 298900
rect 298914 298872 298942 298900
rect 296457 293147 296485 293175
rect 296519 293147 296547 293175
rect 296581 293147 296609 293175
rect 296643 293147 296671 293175
rect 296457 293085 296485 293113
rect 296519 293085 296547 293113
rect 296581 293085 296609 293113
rect 296643 293085 296671 293113
rect 296457 293023 296485 293051
rect 296519 293023 296547 293051
rect 296581 293023 296609 293051
rect 296643 293023 296671 293051
rect 296457 292961 296485 292989
rect 296519 292961 296547 292989
rect 296581 292961 296609 292989
rect 296643 292961 296671 292989
rect 296457 284147 296485 284175
rect 296519 284147 296547 284175
rect 296581 284147 296609 284175
rect 296643 284147 296671 284175
rect 296457 284085 296485 284113
rect 296519 284085 296547 284113
rect 296581 284085 296609 284113
rect 296643 284085 296671 284113
rect 296457 284023 296485 284051
rect 296519 284023 296547 284051
rect 296581 284023 296609 284051
rect 296643 284023 296671 284051
rect 296457 283961 296485 283989
rect 296519 283961 296547 283989
rect 296581 283961 296609 283989
rect 296643 283961 296671 283989
rect 296457 275147 296485 275175
rect 296519 275147 296547 275175
rect 296581 275147 296609 275175
rect 296643 275147 296671 275175
rect 296457 275085 296485 275113
rect 296519 275085 296547 275113
rect 296581 275085 296609 275113
rect 296643 275085 296671 275113
rect 296457 275023 296485 275051
rect 296519 275023 296547 275051
rect 296581 275023 296609 275051
rect 296643 275023 296671 275051
rect 296457 274961 296485 274989
rect 296519 274961 296547 274989
rect 296581 274961 296609 274989
rect 296643 274961 296671 274989
rect 296457 266147 296485 266175
rect 296519 266147 296547 266175
rect 296581 266147 296609 266175
rect 296643 266147 296671 266175
rect 296457 266085 296485 266113
rect 296519 266085 296547 266113
rect 296581 266085 296609 266113
rect 296643 266085 296671 266113
rect 296457 266023 296485 266051
rect 296519 266023 296547 266051
rect 296581 266023 296609 266051
rect 296643 266023 296671 266051
rect 296457 265961 296485 265989
rect 296519 265961 296547 265989
rect 296581 265961 296609 265989
rect 296643 265961 296671 265989
rect 296457 257147 296485 257175
rect 296519 257147 296547 257175
rect 296581 257147 296609 257175
rect 296643 257147 296671 257175
rect 296457 257085 296485 257113
rect 296519 257085 296547 257113
rect 296581 257085 296609 257113
rect 296643 257085 296671 257113
rect 296457 257023 296485 257051
rect 296519 257023 296547 257051
rect 296581 257023 296609 257051
rect 296643 257023 296671 257051
rect 296457 256961 296485 256989
rect 296519 256961 296547 256989
rect 296581 256961 296609 256989
rect 296643 256961 296671 256989
rect 296457 248147 296485 248175
rect 296519 248147 296547 248175
rect 296581 248147 296609 248175
rect 296643 248147 296671 248175
rect 296457 248085 296485 248113
rect 296519 248085 296547 248113
rect 296581 248085 296609 248113
rect 296643 248085 296671 248113
rect 296457 248023 296485 248051
rect 296519 248023 296547 248051
rect 296581 248023 296609 248051
rect 296643 248023 296671 248051
rect 296457 247961 296485 247989
rect 296519 247961 296547 247989
rect 296581 247961 296609 247989
rect 296643 247961 296671 247989
rect 296457 239147 296485 239175
rect 296519 239147 296547 239175
rect 296581 239147 296609 239175
rect 296643 239147 296671 239175
rect 296457 239085 296485 239113
rect 296519 239085 296547 239113
rect 296581 239085 296609 239113
rect 296643 239085 296671 239113
rect 296457 239023 296485 239051
rect 296519 239023 296547 239051
rect 296581 239023 296609 239051
rect 296643 239023 296671 239051
rect 296457 238961 296485 238989
rect 296519 238961 296547 238989
rect 296581 238961 296609 238989
rect 296643 238961 296671 238989
rect 296457 230147 296485 230175
rect 296519 230147 296547 230175
rect 296581 230147 296609 230175
rect 296643 230147 296671 230175
rect 296457 230085 296485 230113
rect 296519 230085 296547 230113
rect 296581 230085 296609 230113
rect 296643 230085 296671 230113
rect 296457 230023 296485 230051
rect 296519 230023 296547 230051
rect 296581 230023 296609 230051
rect 296643 230023 296671 230051
rect 296457 229961 296485 229989
rect 296519 229961 296547 229989
rect 296581 229961 296609 229989
rect 296643 229961 296671 229989
rect 296457 221147 296485 221175
rect 296519 221147 296547 221175
rect 296581 221147 296609 221175
rect 296643 221147 296671 221175
rect 296457 221085 296485 221113
rect 296519 221085 296547 221113
rect 296581 221085 296609 221113
rect 296643 221085 296671 221113
rect 296457 221023 296485 221051
rect 296519 221023 296547 221051
rect 296581 221023 296609 221051
rect 296643 221023 296671 221051
rect 296457 220961 296485 220989
rect 296519 220961 296547 220989
rect 296581 220961 296609 220989
rect 296643 220961 296671 220989
rect 296457 212147 296485 212175
rect 296519 212147 296547 212175
rect 296581 212147 296609 212175
rect 296643 212147 296671 212175
rect 296457 212085 296485 212113
rect 296519 212085 296547 212113
rect 296581 212085 296609 212113
rect 296643 212085 296671 212113
rect 296457 212023 296485 212051
rect 296519 212023 296547 212051
rect 296581 212023 296609 212051
rect 296643 212023 296671 212051
rect 296457 211961 296485 211989
rect 296519 211961 296547 211989
rect 296581 211961 296609 211989
rect 296643 211961 296671 211989
rect 296457 203147 296485 203175
rect 296519 203147 296547 203175
rect 296581 203147 296609 203175
rect 296643 203147 296671 203175
rect 296457 203085 296485 203113
rect 296519 203085 296547 203113
rect 296581 203085 296609 203113
rect 296643 203085 296671 203113
rect 296457 203023 296485 203051
rect 296519 203023 296547 203051
rect 296581 203023 296609 203051
rect 296643 203023 296671 203051
rect 296457 202961 296485 202989
rect 296519 202961 296547 202989
rect 296581 202961 296609 202989
rect 296643 202961 296671 202989
rect 296457 194147 296485 194175
rect 296519 194147 296547 194175
rect 296581 194147 296609 194175
rect 296643 194147 296671 194175
rect 296457 194085 296485 194113
rect 296519 194085 296547 194113
rect 296581 194085 296609 194113
rect 296643 194085 296671 194113
rect 296457 194023 296485 194051
rect 296519 194023 296547 194051
rect 296581 194023 296609 194051
rect 296643 194023 296671 194051
rect 296457 193961 296485 193989
rect 296519 193961 296547 193989
rect 296581 193961 296609 193989
rect 296643 193961 296671 193989
rect 296457 185147 296485 185175
rect 296519 185147 296547 185175
rect 296581 185147 296609 185175
rect 296643 185147 296671 185175
rect 296457 185085 296485 185113
rect 296519 185085 296547 185113
rect 296581 185085 296609 185113
rect 296643 185085 296671 185113
rect 296457 185023 296485 185051
rect 296519 185023 296547 185051
rect 296581 185023 296609 185051
rect 296643 185023 296671 185051
rect 296457 184961 296485 184989
rect 296519 184961 296547 184989
rect 296581 184961 296609 184989
rect 296643 184961 296671 184989
rect 296457 176147 296485 176175
rect 296519 176147 296547 176175
rect 296581 176147 296609 176175
rect 296643 176147 296671 176175
rect 296457 176085 296485 176113
rect 296519 176085 296547 176113
rect 296581 176085 296609 176113
rect 296643 176085 296671 176113
rect 296457 176023 296485 176051
rect 296519 176023 296547 176051
rect 296581 176023 296609 176051
rect 296643 176023 296671 176051
rect 296457 175961 296485 175989
rect 296519 175961 296547 175989
rect 296581 175961 296609 175989
rect 296643 175961 296671 175989
rect 296457 167147 296485 167175
rect 296519 167147 296547 167175
rect 296581 167147 296609 167175
rect 296643 167147 296671 167175
rect 296457 167085 296485 167113
rect 296519 167085 296547 167113
rect 296581 167085 296609 167113
rect 296643 167085 296671 167113
rect 296457 167023 296485 167051
rect 296519 167023 296547 167051
rect 296581 167023 296609 167051
rect 296643 167023 296671 167051
rect 296457 166961 296485 166989
rect 296519 166961 296547 166989
rect 296581 166961 296609 166989
rect 296643 166961 296671 166989
rect 296457 158147 296485 158175
rect 296519 158147 296547 158175
rect 296581 158147 296609 158175
rect 296643 158147 296671 158175
rect 296457 158085 296485 158113
rect 296519 158085 296547 158113
rect 296581 158085 296609 158113
rect 296643 158085 296671 158113
rect 296457 158023 296485 158051
rect 296519 158023 296547 158051
rect 296581 158023 296609 158051
rect 296643 158023 296671 158051
rect 296457 157961 296485 157989
rect 296519 157961 296547 157989
rect 296581 157961 296609 157989
rect 296643 157961 296671 157989
rect 296457 149147 296485 149175
rect 296519 149147 296547 149175
rect 296581 149147 296609 149175
rect 296643 149147 296671 149175
rect 296457 149085 296485 149113
rect 296519 149085 296547 149113
rect 296581 149085 296609 149113
rect 296643 149085 296671 149113
rect 296457 149023 296485 149051
rect 296519 149023 296547 149051
rect 296581 149023 296609 149051
rect 296643 149023 296671 149051
rect 296457 148961 296485 148989
rect 296519 148961 296547 148989
rect 296581 148961 296609 148989
rect 296643 148961 296671 148989
rect 296457 140147 296485 140175
rect 296519 140147 296547 140175
rect 296581 140147 296609 140175
rect 296643 140147 296671 140175
rect 296457 140085 296485 140113
rect 296519 140085 296547 140113
rect 296581 140085 296609 140113
rect 296643 140085 296671 140113
rect 296457 140023 296485 140051
rect 296519 140023 296547 140051
rect 296581 140023 296609 140051
rect 296643 140023 296671 140051
rect 296457 139961 296485 139989
rect 296519 139961 296547 139989
rect 296581 139961 296609 139989
rect 296643 139961 296671 139989
rect 296457 131147 296485 131175
rect 296519 131147 296547 131175
rect 296581 131147 296609 131175
rect 296643 131147 296671 131175
rect 296457 131085 296485 131113
rect 296519 131085 296547 131113
rect 296581 131085 296609 131113
rect 296643 131085 296671 131113
rect 296457 131023 296485 131051
rect 296519 131023 296547 131051
rect 296581 131023 296609 131051
rect 296643 131023 296671 131051
rect 296457 130961 296485 130989
rect 296519 130961 296547 130989
rect 296581 130961 296609 130989
rect 296643 130961 296671 130989
rect 296457 122147 296485 122175
rect 296519 122147 296547 122175
rect 296581 122147 296609 122175
rect 296643 122147 296671 122175
rect 296457 122085 296485 122113
rect 296519 122085 296547 122113
rect 296581 122085 296609 122113
rect 296643 122085 296671 122113
rect 296457 122023 296485 122051
rect 296519 122023 296547 122051
rect 296581 122023 296609 122051
rect 296643 122023 296671 122051
rect 296457 121961 296485 121989
rect 296519 121961 296547 121989
rect 296581 121961 296609 121989
rect 296643 121961 296671 121989
rect 296457 113147 296485 113175
rect 296519 113147 296547 113175
rect 296581 113147 296609 113175
rect 296643 113147 296671 113175
rect 296457 113085 296485 113113
rect 296519 113085 296547 113113
rect 296581 113085 296609 113113
rect 296643 113085 296671 113113
rect 296457 113023 296485 113051
rect 296519 113023 296547 113051
rect 296581 113023 296609 113051
rect 296643 113023 296671 113051
rect 296457 112961 296485 112989
rect 296519 112961 296547 112989
rect 296581 112961 296609 112989
rect 296643 112961 296671 112989
rect 296457 104147 296485 104175
rect 296519 104147 296547 104175
rect 296581 104147 296609 104175
rect 296643 104147 296671 104175
rect 296457 104085 296485 104113
rect 296519 104085 296547 104113
rect 296581 104085 296609 104113
rect 296643 104085 296671 104113
rect 296457 104023 296485 104051
rect 296519 104023 296547 104051
rect 296581 104023 296609 104051
rect 296643 104023 296671 104051
rect 296457 103961 296485 103989
rect 296519 103961 296547 103989
rect 296581 103961 296609 103989
rect 296643 103961 296671 103989
rect 296457 95147 296485 95175
rect 296519 95147 296547 95175
rect 296581 95147 296609 95175
rect 296643 95147 296671 95175
rect 296457 95085 296485 95113
rect 296519 95085 296547 95113
rect 296581 95085 296609 95113
rect 296643 95085 296671 95113
rect 296457 95023 296485 95051
rect 296519 95023 296547 95051
rect 296581 95023 296609 95051
rect 296643 95023 296671 95051
rect 296457 94961 296485 94989
rect 296519 94961 296547 94989
rect 296581 94961 296609 94989
rect 296643 94961 296671 94989
rect 296457 86147 296485 86175
rect 296519 86147 296547 86175
rect 296581 86147 296609 86175
rect 296643 86147 296671 86175
rect 296457 86085 296485 86113
rect 296519 86085 296547 86113
rect 296581 86085 296609 86113
rect 296643 86085 296671 86113
rect 296457 86023 296485 86051
rect 296519 86023 296547 86051
rect 296581 86023 296609 86051
rect 296643 86023 296671 86051
rect 296457 85961 296485 85989
rect 296519 85961 296547 85989
rect 296581 85961 296609 85989
rect 296643 85961 296671 85989
rect 296457 77147 296485 77175
rect 296519 77147 296547 77175
rect 296581 77147 296609 77175
rect 296643 77147 296671 77175
rect 296457 77085 296485 77113
rect 296519 77085 296547 77113
rect 296581 77085 296609 77113
rect 296643 77085 296671 77113
rect 296457 77023 296485 77051
rect 296519 77023 296547 77051
rect 296581 77023 296609 77051
rect 296643 77023 296671 77051
rect 296457 76961 296485 76989
rect 296519 76961 296547 76989
rect 296581 76961 296609 76989
rect 296643 76961 296671 76989
rect 296457 68147 296485 68175
rect 296519 68147 296547 68175
rect 296581 68147 296609 68175
rect 296643 68147 296671 68175
rect 296457 68085 296485 68113
rect 296519 68085 296547 68113
rect 296581 68085 296609 68113
rect 296643 68085 296671 68113
rect 296457 68023 296485 68051
rect 296519 68023 296547 68051
rect 296581 68023 296609 68051
rect 296643 68023 296671 68051
rect 296457 67961 296485 67989
rect 296519 67961 296547 67989
rect 296581 67961 296609 67989
rect 296643 67961 296671 67989
rect 296457 59147 296485 59175
rect 296519 59147 296547 59175
rect 296581 59147 296609 59175
rect 296643 59147 296671 59175
rect 296457 59085 296485 59113
rect 296519 59085 296547 59113
rect 296581 59085 296609 59113
rect 296643 59085 296671 59113
rect 296457 59023 296485 59051
rect 296519 59023 296547 59051
rect 296581 59023 296609 59051
rect 296643 59023 296671 59051
rect 296457 58961 296485 58989
rect 296519 58961 296547 58989
rect 296581 58961 296609 58989
rect 296643 58961 296671 58989
rect 294597 56147 294625 56175
rect 294659 56147 294687 56175
rect 294721 56147 294749 56175
rect 294783 56147 294811 56175
rect 294597 56085 294625 56113
rect 294659 56085 294687 56113
rect 294721 56085 294749 56113
rect 294783 56085 294811 56113
rect 294597 56023 294625 56051
rect 294659 56023 294687 56051
rect 294721 56023 294749 56051
rect 294783 56023 294811 56051
rect 294597 55961 294625 55989
rect 294659 55961 294687 55989
rect 294721 55961 294749 55989
rect 294783 55961 294811 55989
rect 281097 50147 281125 50175
rect 281159 50147 281187 50175
rect 281221 50147 281249 50175
rect 281283 50147 281311 50175
rect 281097 50085 281125 50113
rect 281159 50085 281187 50113
rect 281221 50085 281249 50113
rect 281283 50085 281311 50113
rect 281097 50023 281125 50051
rect 281159 50023 281187 50051
rect 281221 50023 281249 50051
rect 281283 50023 281311 50051
rect 281097 49961 281125 49989
rect 281159 49961 281187 49989
rect 281221 49961 281249 49989
rect 281283 49961 281311 49989
rect 284739 47147 284767 47175
rect 284801 47147 284829 47175
rect 284739 47085 284767 47113
rect 284801 47085 284829 47113
rect 284739 47023 284767 47051
rect 284801 47023 284829 47051
rect 284739 46961 284767 46989
rect 284801 46961 284829 46989
rect 296457 50147 296485 50175
rect 296519 50147 296547 50175
rect 296581 50147 296609 50175
rect 296643 50147 296671 50175
rect 296457 50085 296485 50113
rect 296519 50085 296547 50113
rect 296581 50085 296609 50113
rect 296643 50085 296671 50113
rect 296457 50023 296485 50051
rect 296519 50023 296547 50051
rect 296581 50023 296609 50051
rect 296643 50023 296671 50051
rect 296457 49961 296485 49989
rect 296519 49961 296547 49989
rect 296581 49961 296609 49989
rect 296643 49961 296671 49989
rect 294597 47147 294625 47175
rect 294659 47147 294687 47175
rect 294721 47147 294749 47175
rect 294783 47147 294811 47175
rect 294597 47085 294625 47113
rect 294659 47085 294687 47113
rect 294721 47085 294749 47113
rect 294783 47085 294811 47113
rect 294597 47023 294625 47051
rect 294659 47023 294687 47051
rect 294721 47023 294749 47051
rect 294783 47023 294811 47051
rect 294597 46961 294625 46989
rect 294659 46961 294687 46989
rect 294721 46961 294749 46989
rect 294783 46961 294811 46989
rect 281097 41147 281125 41175
rect 281159 41147 281187 41175
rect 281221 41147 281249 41175
rect 281283 41147 281311 41175
rect 281097 41085 281125 41113
rect 281159 41085 281187 41113
rect 281221 41085 281249 41113
rect 281283 41085 281311 41113
rect 281097 41023 281125 41051
rect 281159 41023 281187 41051
rect 281221 41023 281249 41051
rect 281283 41023 281311 41051
rect 281097 40961 281125 40989
rect 281159 40961 281187 40989
rect 281221 40961 281249 40989
rect 281283 40961 281311 40989
rect 284739 38147 284767 38175
rect 284801 38147 284829 38175
rect 284739 38085 284767 38113
rect 284801 38085 284829 38113
rect 284739 38023 284767 38051
rect 284801 38023 284829 38051
rect 284739 37961 284767 37989
rect 284801 37961 284829 37989
rect 294597 38147 294625 38175
rect 294659 38147 294687 38175
rect 294721 38147 294749 38175
rect 294783 38147 294811 38175
rect 294597 38085 294625 38113
rect 294659 38085 294687 38113
rect 294721 38085 294749 38113
rect 294783 38085 294811 38113
rect 294597 38023 294625 38051
rect 294659 38023 294687 38051
rect 294721 38023 294749 38051
rect 294783 38023 294811 38051
rect 294597 37961 294625 37989
rect 294659 37961 294687 37989
rect 294721 37961 294749 37989
rect 294783 37961 294811 37989
rect 281097 32147 281125 32175
rect 281159 32147 281187 32175
rect 281221 32147 281249 32175
rect 281283 32147 281311 32175
rect 281097 32085 281125 32113
rect 281159 32085 281187 32113
rect 281221 32085 281249 32113
rect 281283 32085 281311 32113
rect 281097 32023 281125 32051
rect 281159 32023 281187 32051
rect 281221 32023 281249 32051
rect 281283 32023 281311 32051
rect 281097 31961 281125 31989
rect 281159 31961 281187 31989
rect 281221 31961 281249 31989
rect 281283 31961 281311 31989
rect 284739 29147 284767 29175
rect 284801 29147 284829 29175
rect 284739 29085 284767 29113
rect 284801 29085 284829 29113
rect 284739 29023 284767 29051
rect 284801 29023 284829 29051
rect 284739 28961 284767 28989
rect 284801 28961 284829 28989
rect 294597 29147 294625 29175
rect 294659 29147 294687 29175
rect 294721 29147 294749 29175
rect 294783 29147 294811 29175
rect 294597 29085 294625 29113
rect 294659 29085 294687 29113
rect 294721 29085 294749 29113
rect 294783 29085 294811 29113
rect 294597 29023 294625 29051
rect 294659 29023 294687 29051
rect 294721 29023 294749 29051
rect 294783 29023 294811 29051
rect 294597 28961 294625 28989
rect 294659 28961 294687 28989
rect 294721 28961 294749 28989
rect 294783 28961 294811 28989
rect 281097 23147 281125 23175
rect 281159 23147 281187 23175
rect 281221 23147 281249 23175
rect 281283 23147 281311 23175
rect 281097 23085 281125 23113
rect 281159 23085 281187 23113
rect 281221 23085 281249 23113
rect 281283 23085 281311 23113
rect 281097 23023 281125 23051
rect 281159 23023 281187 23051
rect 281221 23023 281249 23051
rect 281283 23023 281311 23051
rect 281097 22961 281125 22989
rect 281159 22961 281187 22989
rect 281221 22961 281249 22989
rect 281283 22961 281311 22989
rect 284739 20147 284767 20175
rect 284801 20147 284829 20175
rect 284739 20085 284767 20113
rect 284801 20085 284829 20113
rect 284739 20023 284767 20051
rect 284801 20023 284829 20051
rect 284739 19961 284767 19989
rect 284801 19961 284829 19989
rect 294597 20147 294625 20175
rect 294659 20147 294687 20175
rect 294721 20147 294749 20175
rect 294783 20147 294811 20175
rect 294597 20085 294625 20113
rect 294659 20085 294687 20113
rect 294721 20085 294749 20113
rect 294783 20085 294811 20113
rect 294597 20023 294625 20051
rect 294659 20023 294687 20051
rect 294721 20023 294749 20051
rect 294783 20023 294811 20051
rect 294597 19961 294625 19989
rect 294659 19961 294687 19989
rect 294721 19961 294749 19989
rect 294783 19961 294811 19989
rect 281097 14147 281125 14175
rect 281159 14147 281187 14175
rect 281221 14147 281249 14175
rect 281283 14147 281311 14175
rect 281097 14085 281125 14113
rect 281159 14085 281187 14113
rect 281221 14085 281249 14113
rect 281283 14085 281311 14113
rect 281097 14023 281125 14051
rect 281159 14023 281187 14051
rect 281221 14023 281249 14051
rect 281283 14023 281311 14051
rect 281097 13961 281125 13989
rect 281159 13961 281187 13989
rect 281221 13961 281249 13989
rect 281283 13961 281311 13989
rect 284739 11147 284767 11175
rect 284801 11147 284829 11175
rect 284739 11085 284767 11113
rect 284801 11085 284829 11113
rect 284739 11023 284767 11051
rect 284801 11023 284829 11051
rect 284739 10961 284767 10989
rect 284801 10961 284829 10989
rect 294597 11147 294625 11175
rect 294659 11147 294687 11175
rect 294721 11147 294749 11175
rect 294783 11147 294811 11175
rect 294597 11085 294625 11113
rect 294659 11085 294687 11113
rect 294721 11085 294749 11113
rect 294783 11085 294811 11113
rect 294597 11023 294625 11051
rect 294659 11023 294687 11051
rect 294721 11023 294749 11051
rect 294783 11023 294811 11051
rect 294597 10961 294625 10989
rect 294659 10961 294687 10989
rect 294721 10961 294749 10989
rect 294783 10961 294811 10989
rect 281097 5147 281125 5175
rect 281159 5147 281187 5175
rect 281221 5147 281249 5175
rect 281283 5147 281311 5175
rect 281097 5085 281125 5113
rect 281159 5085 281187 5113
rect 281221 5085 281249 5113
rect 281283 5085 281311 5113
rect 281097 5023 281125 5051
rect 281159 5023 281187 5051
rect 281221 5023 281249 5051
rect 281283 5023 281311 5051
rect 281097 4961 281125 4989
rect 281159 4961 281187 4989
rect 281221 4961 281249 4989
rect 281283 4961 281311 4989
rect 281097 -588 281125 -560
rect 281159 -588 281187 -560
rect 281221 -588 281249 -560
rect 281283 -588 281311 -560
rect 281097 -650 281125 -622
rect 281159 -650 281187 -622
rect 281221 -650 281249 -622
rect 281283 -650 281311 -622
rect 281097 -712 281125 -684
rect 281159 -712 281187 -684
rect 281221 -712 281249 -684
rect 281283 -712 281311 -684
rect 281097 -774 281125 -746
rect 281159 -774 281187 -746
rect 281221 -774 281249 -746
rect 281283 -774 281311 -746
rect 296457 41147 296485 41175
rect 296519 41147 296547 41175
rect 296581 41147 296609 41175
rect 296643 41147 296671 41175
rect 296457 41085 296485 41113
rect 296519 41085 296547 41113
rect 296581 41085 296609 41113
rect 296643 41085 296671 41113
rect 296457 41023 296485 41051
rect 296519 41023 296547 41051
rect 296581 41023 296609 41051
rect 296643 41023 296671 41051
rect 296457 40961 296485 40989
rect 296519 40961 296547 40989
rect 296581 40961 296609 40989
rect 296643 40961 296671 40989
rect 296457 32147 296485 32175
rect 296519 32147 296547 32175
rect 296581 32147 296609 32175
rect 296643 32147 296671 32175
rect 296457 32085 296485 32113
rect 296519 32085 296547 32113
rect 296581 32085 296609 32113
rect 296643 32085 296671 32113
rect 296457 32023 296485 32051
rect 296519 32023 296547 32051
rect 296581 32023 296609 32051
rect 296643 32023 296671 32051
rect 296457 31961 296485 31989
rect 296519 31961 296547 31989
rect 296581 31961 296609 31989
rect 296643 31961 296671 31989
rect 296457 23147 296485 23175
rect 296519 23147 296547 23175
rect 296581 23147 296609 23175
rect 296643 23147 296671 23175
rect 296457 23085 296485 23113
rect 296519 23085 296547 23113
rect 296581 23085 296609 23113
rect 296643 23085 296671 23113
rect 296457 23023 296485 23051
rect 296519 23023 296547 23051
rect 296581 23023 296609 23051
rect 296643 23023 296671 23051
rect 296457 22961 296485 22989
rect 296519 22961 296547 22989
rect 296581 22961 296609 22989
rect 296643 22961 296671 22989
rect 296457 14147 296485 14175
rect 296519 14147 296547 14175
rect 296581 14147 296609 14175
rect 296643 14147 296671 14175
rect 296457 14085 296485 14113
rect 296519 14085 296547 14113
rect 296581 14085 296609 14113
rect 296643 14085 296671 14113
rect 296457 14023 296485 14051
rect 296519 14023 296547 14051
rect 296581 14023 296609 14051
rect 296643 14023 296671 14051
rect 296457 13961 296485 13989
rect 296519 13961 296547 13989
rect 296581 13961 296609 13989
rect 296643 13961 296671 13989
rect 296457 5147 296485 5175
rect 296519 5147 296547 5175
rect 296581 5147 296609 5175
rect 296643 5147 296671 5175
rect 296457 5085 296485 5113
rect 296519 5085 296547 5113
rect 296581 5085 296609 5113
rect 296643 5085 296671 5113
rect 296457 5023 296485 5051
rect 296519 5023 296547 5051
rect 296581 5023 296609 5051
rect 296643 5023 296671 5051
rect 296457 4961 296485 4989
rect 296519 4961 296547 4989
rect 296581 4961 296609 4989
rect 296643 4961 296671 4989
rect 294597 2147 294625 2175
rect 294659 2147 294687 2175
rect 294721 2147 294749 2175
rect 294783 2147 294811 2175
rect 294597 2085 294625 2113
rect 294659 2085 294687 2113
rect 294721 2085 294749 2113
rect 294783 2085 294811 2113
rect 294597 2023 294625 2051
rect 294659 2023 294687 2051
rect 294721 2023 294749 2051
rect 294783 2023 294811 2051
rect 294597 1961 294625 1989
rect 294659 1961 294687 1989
rect 294721 1961 294749 1989
rect 294783 1961 294811 1989
rect 294597 -108 294625 -80
rect 294659 -108 294687 -80
rect 294721 -108 294749 -80
rect 294783 -108 294811 -80
rect 294597 -170 294625 -142
rect 294659 -170 294687 -142
rect 294721 -170 294749 -142
rect 294783 -170 294811 -142
rect 294597 -232 294625 -204
rect 294659 -232 294687 -204
rect 294721 -232 294749 -204
rect 294783 -232 294811 -204
rect 294597 -294 294625 -266
rect 294659 -294 294687 -266
rect 294721 -294 294749 -266
rect 294783 -294 294811 -266
rect 298248 298578 298276 298606
rect 298310 298578 298338 298606
rect 298372 298578 298400 298606
rect 298434 298578 298462 298606
rect 298248 298516 298276 298544
rect 298310 298516 298338 298544
rect 298372 298516 298400 298544
rect 298434 298516 298462 298544
rect 298248 298454 298276 298482
rect 298310 298454 298338 298482
rect 298372 298454 298400 298482
rect 298434 298454 298462 298482
rect 298248 298392 298276 298420
rect 298310 298392 298338 298420
rect 298372 298392 298400 298420
rect 298434 298392 298462 298420
rect 298248 290147 298276 290175
rect 298310 290147 298338 290175
rect 298372 290147 298400 290175
rect 298434 290147 298462 290175
rect 298248 290085 298276 290113
rect 298310 290085 298338 290113
rect 298372 290085 298400 290113
rect 298434 290085 298462 290113
rect 298248 290023 298276 290051
rect 298310 290023 298338 290051
rect 298372 290023 298400 290051
rect 298434 290023 298462 290051
rect 298248 289961 298276 289989
rect 298310 289961 298338 289989
rect 298372 289961 298400 289989
rect 298434 289961 298462 289989
rect 298248 281147 298276 281175
rect 298310 281147 298338 281175
rect 298372 281147 298400 281175
rect 298434 281147 298462 281175
rect 298248 281085 298276 281113
rect 298310 281085 298338 281113
rect 298372 281085 298400 281113
rect 298434 281085 298462 281113
rect 298248 281023 298276 281051
rect 298310 281023 298338 281051
rect 298372 281023 298400 281051
rect 298434 281023 298462 281051
rect 298248 280961 298276 280989
rect 298310 280961 298338 280989
rect 298372 280961 298400 280989
rect 298434 280961 298462 280989
rect 298248 272147 298276 272175
rect 298310 272147 298338 272175
rect 298372 272147 298400 272175
rect 298434 272147 298462 272175
rect 298248 272085 298276 272113
rect 298310 272085 298338 272113
rect 298372 272085 298400 272113
rect 298434 272085 298462 272113
rect 298248 272023 298276 272051
rect 298310 272023 298338 272051
rect 298372 272023 298400 272051
rect 298434 272023 298462 272051
rect 298248 271961 298276 271989
rect 298310 271961 298338 271989
rect 298372 271961 298400 271989
rect 298434 271961 298462 271989
rect 298248 263147 298276 263175
rect 298310 263147 298338 263175
rect 298372 263147 298400 263175
rect 298434 263147 298462 263175
rect 298248 263085 298276 263113
rect 298310 263085 298338 263113
rect 298372 263085 298400 263113
rect 298434 263085 298462 263113
rect 298248 263023 298276 263051
rect 298310 263023 298338 263051
rect 298372 263023 298400 263051
rect 298434 263023 298462 263051
rect 298248 262961 298276 262989
rect 298310 262961 298338 262989
rect 298372 262961 298400 262989
rect 298434 262961 298462 262989
rect 298248 254147 298276 254175
rect 298310 254147 298338 254175
rect 298372 254147 298400 254175
rect 298434 254147 298462 254175
rect 298248 254085 298276 254113
rect 298310 254085 298338 254113
rect 298372 254085 298400 254113
rect 298434 254085 298462 254113
rect 298248 254023 298276 254051
rect 298310 254023 298338 254051
rect 298372 254023 298400 254051
rect 298434 254023 298462 254051
rect 298248 253961 298276 253989
rect 298310 253961 298338 253989
rect 298372 253961 298400 253989
rect 298434 253961 298462 253989
rect 298248 245147 298276 245175
rect 298310 245147 298338 245175
rect 298372 245147 298400 245175
rect 298434 245147 298462 245175
rect 298248 245085 298276 245113
rect 298310 245085 298338 245113
rect 298372 245085 298400 245113
rect 298434 245085 298462 245113
rect 298248 245023 298276 245051
rect 298310 245023 298338 245051
rect 298372 245023 298400 245051
rect 298434 245023 298462 245051
rect 298248 244961 298276 244989
rect 298310 244961 298338 244989
rect 298372 244961 298400 244989
rect 298434 244961 298462 244989
rect 298248 236147 298276 236175
rect 298310 236147 298338 236175
rect 298372 236147 298400 236175
rect 298434 236147 298462 236175
rect 298248 236085 298276 236113
rect 298310 236085 298338 236113
rect 298372 236085 298400 236113
rect 298434 236085 298462 236113
rect 298248 236023 298276 236051
rect 298310 236023 298338 236051
rect 298372 236023 298400 236051
rect 298434 236023 298462 236051
rect 298248 235961 298276 235989
rect 298310 235961 298338 235989
rect 298372 235961 298400 235989
rect 298434 235961 298462 235989
rect 298248 227147 298276 227175
rect 298310 227147 298338 227175
rect 298372 227147 298400 227175
rect 298434 227147 298462 227175
rect 298248 227085 298276 227113
rect 298310 227085 298338 227113
rect 298372 227085 298400 227113
rect 298434 227085 298462 227113
rect 298248 227023 298276 227051
rect 298310 227023 298338 227051
rect 298372 227023 298400 227051
rect 298434 227023 298462 227051
rect 298248 226961 298276 226989
rect 298310 226961 298338 226989
rect 298372 226961 298400 226989
rect 298434 226961 298462 226989
rect 298248 218147 298276 218175
rect 298310 218147 298338 218175
rect 298372 218147 298400 218175
rect 298434 218147 298462 218175
rect 298248 218085 298276 218113
rect 298310 218085 298338 218113
rect 298372 218085 298400 218113
rect 298434 218085 298462 218113
rect 298248 218023 298276 218051
rect 298310 218023 298338 218051
rect 298372 218023 298400 218051
rect 298434 218023 298462 218051
rect 298248 217961 298276 217989
rect 298310 217961 298338 217989
rect 298372 217961 298400 217989
rect 298434 217961 298462 217989
rect 298248 209147 298276 209175
rect 298310 209147 298338 209175
rect 298372 209147 298400 209175
rect 298434 209147 298462 209175
rect 298248 209085 298276 209113
rect 298310 209085 298338 209113
rect 298372 209085 298400 209113
rect 298434 209085 298462 209113
rect 298248 209023 298276 209051
rect 298310 209023 298338 209051
rect 298372 209023 298400 209051
rect 298434 209023 298462 209051
rect 298248 208961 298276 208989
rect 298310 208961 298338 208989
rect 298372 208961 298400 208989
rect 298434 208961 298462 208989
rect 298248 200147 298276 200175
rect 298310 200147 298338 200175
rect 298372 200147 298400 200175
rect 298434 200147 298462 200175
rect 298248 200085 298276 200113
rect 298310 200085 298338 200113
rect 298372 200085 298400 200113
rect 298434 200085 298462 200113
rect 298248 200023 298276 200051
rect 298310 200023 298338 200051
rect 298372 200023 298400 200051
rect 298434 200023 298462 200051
rect 298248 199961 298276 199989
rect 298310 199961 298338 199989
rect 298372 199961 298400 199989
rect 298434 199961 298462 199989
rect 298248 191147 298276 191175
rect 298310 191147 298338 191175
rect 298372 191147 298400 191175
rect 298434 191147 298462 191175
rect 298248 191085 298276 191113
rect 298310 191085 298338 191113
rect 298372 191085 298400 191113
rect 298434 191085 298462 191113
rect 298248 191023 298276 191051
rect 298310 191023 298338 191051
rect 298372 191023 298400 191051
rect 298434 191023 298462 191051
rect 298248 190961 298276 190989
rect 298310 190961 298338 190989
rect 298372 190961 298400 190989
rect 298434 190961 298462 190989
rect 298248 182147 298276 182175
rect 298310 182147 298338 182175
rect 298372 182147 298400 182175
rect 298434 182147 298462 182175
rect 298248 182085 298276 182113
rect 298310 182085 298338 182113
rect 298372 182085 298400 182113
rect 298434 182085 298462 182113
rect 298248 182023 298276 182051
rect 298310 182023 298338 182051
rect 298372 182023 298400 182051
rect 298434 182023 298462 182051
rect 298248 181961 298276 181989
rect 298310 181961 298338 181989
rect 298372 181961 298400 181989
rect 298434 181961 298462 181989
rect 298248 173147 298276 173175
rect 298310 173147 298338 173175
rect 298372 173147 298400 173175
rect 298434 173147 298462 173175
rect 298248 173085 298276 173113
rect 298310 173085 298338 173113
rect 298372 173085 298400 173113
rect 298434 173085 298462 173113
rect 298248 173023 298276 173051
rect 298310 173023 298338 173051
rect 298372 173023 298400 173051
rect 298434 173023 298462 173051
rect 298248 172961 298276 172989
rect 298310 172961 298338 172989
rect 298372 172961 298400 172989
rect 298434 172961 298462 172989
rect 298248 164147 298276 164175
rect 298310 164147 298338 164175
rect 298372 164147 298400 164175
rect 298434 164147 298462 164175
rect 298248 164085 298276 164113
rect 298310 164085 298338 164113
rect 298372 164085 298400 164113
rect 298434 164085 298462 164113
rect 298248 164023 298276 164051
rect 298310 164023 298338 164051
rect 298372 164023 298400 164051
rect 298434 164023 298462 164051
rect 298248 163961 298276 163989
rect 298310 163961 298338 163989
rect 298372 163961 298400 163989
rect 298434 163961 298462 163989
rect 298248 155147 298276 155175
rect 298310 155147 298338 155175
rect 298372 155147 298400 155175
rect 298434 155147 298462 155175
rect 298248 155085 298276 155113
rect 298310 155085 298338 155113
rect 298372 155085 298400 155113
rect 298434 155085 298462 155113
rect 298248 155023 298276 155051
rect 298310 155023 298338 155051
rect 298372 155023 298400 155051
rect 298434 155023 298462 155051
rect 298248 154961 298276 154989
rect 298310 154961 298338 154989
rect 298372 154961 298400 154989
rect 298434 154961 298462 154989
rect 298248 146147 298276 146175
rect 298310 146147 298338 146175
rect 298372 146147 298400 146175
rect 298434 146147 298462 146175
rect 298248 146085 298276 146113
rect 298310 146085 298338 146113
rect 298372 146085 298400 146113
rect 298434 146085 298462 146113
rect 298248 146023 298276 146051
rect 298310 146023 298338 146051
rect 298372 146023 298400 146051
rect 298434 146023 298462 146051
rect 298248 145961 298276 145989
rect 298310 145961 298338 145989
rect 298372 145961 298400 145989
rect 298434 145961 298462 145989
rect 298248 137147 298276 137175
rect 298310 137147 298338 137175
rect 298372 137147 298400 137175
rect 298434 137147 298462 137175
rect 298248 137085 298276 137113
rect 298310 137085 298338 137113
rect 298372 137085 298400 137113
rect 298434 137085 298462 137113
rect 298248 137023 298276 137051
rect 298310 137023 298338 137051
rect 298372 137023 298400 137051
rect 298434 137023 298462 137051
rect 298248 136961 298276 136989
rect 298310 136961 298338 136989
rect 298372 136961 298400 136989
rect 298434 136961 298462 136989
rect 298248 128147 298276 128175
rect 298310 128147 298338 128175
rect 298372 128147 298400 128175
rect 298434 128147 298462 128175
rect 298248 128085 298276 128113
rect 298310 128085 298338 128113
rect 298372 128085 298400 128113
rect 298434 128085 298462 128113
rect 298248 128023 298276 128051
rect 298310 128023 298338 128051
rect 298372 128023 298400 128051
rect 298434 128023 298462 128051
rect 298248 127961 298276 127989
rect 298310 127961 298338 127989
rect 298372 127961 298400 127989
rect 298434 127961 298462 127989
rect 298248 119147 298276 119175
rect 298310 119147 298338 119175
rect 298372 119147 298400 119175
rect 298434 119147 298462 119175
rect 298248 119085 298276 119113
rect 298310 119085 298338 119113
rect 298372 119085 298400 119113
rect 298434 119085 298462 119113
rect 298248 119023 298276 119051
rect 298310 119023 298338 119051
rect 298372 119023 298400 119051
rect 298434 119023 298462 119051
rect 298248 118961 298276 118989
rect 298310 118961 298338 118989
rect 298372 118961 298400 118989
rect 298434 118961 298462 118989
rect 298248 110147 298276 110175
rect 298310 110147 298338 110175
rect 298372 110147 298400 110175
rect 298434 110147 298462 110175
rect 298248 110085 298276 110113
rect 298310 110085 298338 110113
rect 298372 110085 298400 110113
rect 298434 110085 298462 110113
rect 298248 110023 298276 110051
rect 298310 110023 298338 110051
rect 298372 110023 298400 110051
rect 298434 110023 298462 110051
rect 298248 109961 298276 109989
rect 298310 109961 298338 109989
rect 298372 109961 298400 109989
rect 298434 109961 298462 109989
rect 298248 101147 298276 101175
rect 298310 101147 298338 101175
rect 298372 101147 298400 101175
rect 298434 101147 298462 101175
rect 298248 101085 298276 101113
rect 298310 101085 298338 101113
rect 298372 101085 298400 101113
rect 298434 101085 298462 101113
rect 298248 101023 298276 101051
rect 298310 101023 298338 101051
rect 298372 101023 298400 101051
rect 298434 101023 298462 101051
rect 298248 100961 298276 100989
rect 298310 100961 298338 100989
rect 298372 100961 298400 100989
rect 298434 100961 298462 100989
rect 298248 92147 298276 92175
rect 298310 92147 298338 92175
rect 298372 92147 298400 92175
rect 298434 92147 298462 92175
rect 298248 92085 298276 92113
rect 298310 92085 298338 92113
rect 298372 92085 298400 92113
rect 298434 92085 298462 92113
rect 298248 92023 298276 92051
rect 298310 92023 298338 92051
rect 298372 92023 298400 92051
rect 298434 92023 298462 92051
rect 298248 91961 298276 91989
rect 298310 91961 298338 91989
rect 298372 91961 298400 91989
rect 298434 91961 298462 91989
rect 298248 83147 298276 83175
rect 298310 83147 298338 83175
rect 298372 83147 298400 83175
rect 298434 83147 298462 83175
rect 298248 83085 298276 83113
rect 298310 83085 298338 83113
rect 298372 83085 298400 83113
rect 298434 83085 298462 83113
rect 298248 83023 298276 83051
rect 298310 83023 298338 83051
rect 298372 83023 298400 83051
rect 298434 83023 298462 83051
rect 298248 82961 298276 82989
rect 298310 82961 298338 82989
rect 298372 82961 298400 82989
rect 298434 82961 298462 82989
rect 298248 74147 298276 74175
rect 298310 74147 298338 74175
rect 298372 74147 298400 74175
rect 298434 74147 298462 74175
rect 298248 74085 298276 74113
rect 298310 74085 298338 74113
rect 298372 74085 298400 74113
rect 298434 74085 298462 74113
rect 298248 74023 298276 74051
rect 298310 74023 298338 74051
rect 298372 74023 298400 74051
rect 298434 74023 298462 74051
rect 298248 73961 298276 73989
rect 298310 73961 298338 73989
rect 298372 73961 298400 73989
rect 298434 73961 298462 73989
rect 298248 65147 298276 65175
rect 298310 65147 298338 65175
rect 298372 65147 298400 65175
rect 298434 65147 298462 65175
rect 298248 65085 298276 65113
rect 298310 65085 298338 65113
rect 298372 65085 298400 65113
rect 298434 65085 298462 65113
rect 298248 65023 298276 65051
rect 298310 65023 298338 65051
rect 298372 65023 298400 65051
rect 298434 65023 298462 65051
rect 298248 64961 298276 64989
rect 298310 64961 298338 64989
rect 298372 64961 298400 64989
rect 298434 64961 298462 64989
rect 298248 56147 298276 56175
rect 298310 56147 298338 56175
rect 298372 56147 298400 56175
rect 298434 56147 298462 56175
rect 298248 56085 298276 56113
rect 298310 56085 298338 56113
rect 298372 56085 298400 56113
rect 298434 56085 298462 56113
rect 298248 56023 298276 56051
rect 298310 56023 298338 56051
rect 298372 56023 298400 56051
rect 298434 56023 298462 56051
rect 298248 55961 298276 55989
rect 298310 55961 298338 55989
rect 298372 55961 298400 55989
rect 298434 55961 298462 55989
rect 298248 47147 298276 47175
rect 298310 47147 298338 47175
rect 298372 47147 298400 47175
rect 298434 47147 298462 47175
rect 298248 47085 298276 47113
rect 298310 47085 298338 47113
rect 298372 47085 298400 47113
rect 298434 47085 298462 47113
rect 298248 47023 298276 47051
rect 298310 47023 298338 47051
rect 298372 47023 298400 47051
rect 298434 47023 298462 47051
rect 298248 46961 298276 46989
rect 298310 46961 298338 46989
rect 298372 46961 298400 46989
rect 298434 46961 298462 46989
rect 298248 38147 298276 38175
rect 298310 38147 298338 38175
rect 298372 38147 298400 38175
rect 298434 38147 298462 38175
rect 298248 38085 298276 38113
rect 298310 38085 298338 38113
rect 298372 38085 298400 38113
rect 298434 38085 298462 38113
rect 298248 38023 298276 38051
rect 298310 38023 298338 38051
rect 298372 38023 298400 38051
rect 298434 38023 298462 38051
rect 298248 37961 298276 37989
rect 298310 37961 298338 37989
rect 298372 37961 298400 37989
rect 298434 37961 298462 37989
rect 298248 29147 298276 29175
rect 298310 29147 298338 29175
rect 298372 29147 298400 29175
rect 298434 29147 298462 29175
rect 298248 29085 298276 29113
rect 298310 29085 298338 29113
rect 298372 29085 298400 29113
rect 298434 29085 298462 29113
rect 298248 29023 298276 29051
rect 298310 29023 298338 29051
rect 298372 29023 298400 29051
rect 298434 29023 298462 29051
rect 298248 28961 298276 28989
rect 298310 28961 298338 28989
rect 298372 28961 298400 28989
rect 298434 28961 298462 28989
rect 298248 20147 298276 20175
rect 298310 20147 298338 20175
rect 298372 20147 298400 20175
rect 298434 20147 298462 20175
rect 298248 20085 298276 20113
rect 298310 20085 298338 20113
rect 298372 20085 298400 20113
rect 298434 20085 298462 20113
rect 298248 20023 298276 20051
rect 298310 20023 298338 20051
rect 298372 20023 298400 20051
rect 298434 20023 298462 20051
rect 298248 19961 298276 19989
rect 298310 19961 298338 19989
rect 298372 19961 298400 19989
rect 298434 19961 298462 19989
rect 298248 11147 298276 11175
rect 298310 11147 298338 11175
rect 298372 11147 298400 11175
rect 298434 11147 298462 11175
rect 298248 11085 298276 11113
rect 298310 11085 298338 11113
rect 298372 11085 298400 11113
rect 298434 11085 298462 11113
rect 298248 11023 298276 11051
rect 298310 11023 298338 11051
rect 298372 11023 298400 11051
rect 298434 11023 298462 11051
rect 298248 10961 298276 10989
rect 298310 10961 298338 10989
rect 298372 10961 298400 10989
rect 298434 10961 298462 10989
rect 298248 2147 298276 2175
rect 298310 2147 298338 2175
rect 298372 2147 298400 2175
rect 298434 2147 298462 2175
rect 298248 2085 298276 2113
rect 298310 2085 298338 2113
rect 298372 2085 298400 2113
rect 298434 2085 298462 2113
rect 298248 2023 298276 2051
rect 298310 2023 298338 2051
rect 298372 2023 298400 2051
rect 298434 2023 298462 2051
rect 298248 1961 298276 1989
rect 298310 1961 298338 1989
rect 298372 1961 298400 1989
rect 298434 1961 298462 1989
rect 298248 -108 298276 -80
rect 298310 -108 298338 -80
rect 298372 -108 298400 -80
rect 298434 -108 298462 -80
rect 298248 -170 298276 -142
rect 298310 -170 298338 -142
rect 298372 -170 298400 -142
rect 298434 -170 298462 -142
rect 298248 -232 298276 -204
rect 298310 -232 298338 -204
rect 298372 -232 298400 -204
rect 298434 -232 298462 -204
rect 298248 -294 298276 -266
rect 298310 -294 298338 -266
rect 298372 -294 298400 -266
rect 298434 -294 298462 -266
rect 298728 293147 298756 293175
rect 298790 293147 298818 293175
rect 298852 293147 298880 293175
rect 298914 293147 298942 293175
rect 298728 293085 298756 293113
rect 298790 293085 298818 293113
rect 298852 293085 298880 293113
rect 298914 293085 298942 293113
rect 298728 293023 298756 293051
rect 298790 293023 298818 293051
rect 298852 293023 298880 293051
rect 298914 293023 298942 293051
rect 298728 292961 298756 292989
rect 298790 292961 298818 292989
rect 298852 292961 298880 292989
rect 298914 292961 298942 292989
rect 298728 284147 298756 284175
rect 298790 284147 298818 284175
rect 298852 284147 298880 284175
rect 298914 284147 298942 284175
rect 298728 284085 298756 284113
rect 298790 284085 298818 284113
rect 298852 284085 298880 284113
rect 298914 284085 298942 284113
rect 298728 284023 298756 284051
rect 298790 284023 298818 284051
rect 298852 284023 298880 284051
rect 298914 284023 298942 284051
rect 298728 283961 298756 283989
rect 298790 283961 298818 283989
rect 298852 283961 298880 283989
rect 298914 283961 298942 283989
rect 298728 275147 298756 275175
rect 298790 275147 298818 275175
rect 298852 275147 298880 275175
rect 298914 275147 298942 275175
rect 298728 275085 298756 275113
rect 298790 275085 298818 275113
rect 298852 275085 298880 275113
rect 298914 275085 298942 275113
rect 298728 275023 298756 275051
rect 298790 275023 298818 275051
rect 298852 275023 298880 275051
rect 298914 275023 298942 275051
rect 298728 274961 298756 274989
rect 298790 274961 298818 274989
rect 298852 274961 298880 274989
rect 298914 274961 298942 274989
rect 298728 266147 298756 266175
rect 298790 266147 298818 266175
rect 298852 266147 298880 266175
rect 298914 266147 298942 266175
rect 298728 266085 298756 266113
rect 298790 266085 298818 266113
rect 298852 266085 298880 266113
rect 298914 266085 298942 266113
rect 298728 266023 298756 266051
rect 298790 266023 298818 266051
rect 298852 266023 298880 266051
rect 298914 266023 298942 266051
rect 298728 265961 298756 265989
rect 298790 265961 298818 265989
rect 298852 265961 298880 265989
rect 298914 265961 298942 265989
rect 298728 257147 298756 257175
rect 298790 257147 298818 257175
rect 298852 257147 298880 257175
rect 298914 257147 298942 257175
rect 298728 257085 298756 257113
rect 298790 257085 298818 257113
rect 298852 257085 298880 257113
rect 298914 257085 298942 257113
rect 298728 257023 298756 257051
rect 298790 257023 298818 257051
rect 298852 257023 298880 257051
rect 298914 257023 298942 257051
rect 298728 256961 298756 256989
rect 298790 256961 298818 256989
rect 298852 256961 298880 256989
rect 298914 256961 298942 256989
rect 298728 248147 298756 248175
rect 298790 248147 298818 248175
rect 298852 248147 298880 248175
rect 298914 248147 298942 248175
rect 298728 248085 298756 248113
rect 298790 248085 298818 248113
rect 298852 248085 298880 248113
rect 298914 248085 298942 248113
rect 298728 248023 298756 248051
rect 298790 248023 298818 248051
rect 298852 248023 298880 248051
rect 298914 248023 298942 248051
rect 298728 247961 298756 247989
rect 298790 247961 298818 247989
rect 298852 247961 298880 247989
rect 298914 247961 298942 247989
rect 298728 239147 298756 239175
rect 298790 239147 298818 239175
rect 298852 239147 298880 239175
rect 298914 239147 298942 239175
rect 298728 239085 298756 239113
rect 298790 239085 298818 239113
rect 298852 239085 298880 239113
rect 298914 239085 298942 239113
rect 298728 239023 298756 239051
rect 298790 239023 298818 239051
rect 298852 239023 298880 239051
rect 298914 239023 298942 239051
rect 298728 238961 298756 238989
rect 298790 238961 298818 238989
rect 298852 238961 298880 238989
rect 298914 238961 298942 238989
rect 298728 230147 298756 230175
rect 298790 230147 298818 230175
rect 298852 230147 298880 230175
rect 298914 230147 298942 230175
rect 298728 230085 298756 230113
rect 298790 230085 298818 230113
rect 298852 230085 298880 230113
rect 298914 230085 298942 230113
rect 298728 230023 298756 230051
rect 298790 230023 298818 230051
rect 298852 230023 298880 230051
rect 298914 230023 298942 230051
rect 298728 229961 298756 229989
rect 298790 229961 298818 229989
rect 298852 229961 298880 229989
rect 298914 229961 298942 229989
rect 298728 221147 298756 221175
rect 298790 221147 298818 221175
rect 298852 221147 298880 221175
rect 298914 221147 298942 221175
rect 298728 221085 298756 221113
rect 298790 221085 298818 221113
rect 298852 221085 298880 221113
rect 298914 221085 298942 221113
rect 298728 221023 298756 221051
rect 298790 221023 298818 221051
rect 298852 221023 298880 221051
rect 298914 221023 298942 221051
rect 298728 220961 298756 220989
rect 298790 220961 298818 220989
rect 298852 220961 298880 220989
rect 298914 220961 298942 220989
rect 298728 212147 298756 212175
rect 298790 212147 298818 212175
rect 298852 212147 298880 212175
rect 298914 212147 298942 212175
rect 298728 212085 298756 212113
rect 298790 212085 298818 212113
rect 298852 212085 298880 212113
rect 298914 212085 298942 212113
rect 298728 212023 298756 212051
rect 298790 212023 298818 212051
rect 298852 212023 298880 212051
rect 298914 212023 298942 212051
rect 298728 211961 298756 211989
rect 298790 211961 298818 211989
rect 298852 211961 298880 211989
rect 298914 211961 298942 211989
rect 298728 203147 298756 203175
rect 298790 203147 298818 203175
rect 298852 203147 298880 203175
rect 298914 203147 298942 203175
rect 298728 203085 298756 203113
rect 298790 203085 298818 203113
rect 298852 203085 298880 203113
rect 298914 203085 298942 203113
rect 298728 203023 298756 203051
rect 298790 203023 298818 203051
rect 298852 203023 298880 203051
rect 298914 203023 298942 203051
rect 298728 202961 298756 202989
rect 298790 202961 298818 202989
rect 298852 202961 298880 202989
rect 298914 202961 298942 202989
rect 298728 194147 298756 194175
rect 298790 194147 298818 194175
rect 298852 194147 298880 194175
rect 298914 194147 298942 194175
rect 298728 194085 298756 194113
rect 298790 194085 298818 194113
rect 298852 194085 298880 194113
rect 298914 194085 298942 194113
rect 298728 194023 298756 194051
rect 298790 194023 298818 194051
rect 298852 194023 298880 194051
rect 298914 194023 298942 194051
rect 298728 193961 298756 193989
rect 298790 193961 298818 193989
rect 298852 193961 298880 193989
rect 298914 193961 298942 193989
rect 298728 185147 298756 185175
rect 298790 185147 298818 185175
rect 298852 185147 298880 185175
rect 298914 185147 298942 185175
rect 298728 185085 298756 185113
rect 298790 185085 298818 185113
rect 298852 185085 298880 185113
rect 298914 185085 298942 185113
rect 298728 185023 298756 185051
rect 298790 185023 298818 185051
rect 298852 185023 298880 185051
rect 298914 185023 298942 185051
rect 298728 184961 298756 184989
rect 298790 184961 298818 184989
rect 298852 184961 298880 184989
rect 298914 184961 298942 184989
rect 298728 176147 298756 176175
rect 298790 176147 298818 176175
rect 298852 176147 298880 176175
rect 298914 176147 298942 176175
rect 298728 176085 298756 176113
rect 298790 176085 298818 176113
rect 298852 176085 298880 176113
rect 298914 176085 298942 176113
rect 298728 176023 298756 176051
rect 298790 176023 298818 176051
rect 298852 176023 298880 176051
rect 298914 176023 298942 176051
rect 298728 175961 298756 175989
rect 298790 175961 298818 175989
rect 298852 175961 298880 175989
rect 298914 175961 298942 175989
rect 298728 167147 298756 167175
rect 298790 167147 298818 167175
rect 298852 167147 298880 167175
rect 298914 167147 298942 167175
rect 298728 167085 298756 167113
rect 298790 167085 298818 167113
rect 298852 167085 298880 167113
rect 298914 167085 298942 167113
rect 298728 167023 298756 167051
rect 298790 167023 298818 167051
rect 298852 167023 298880 167051
rect 298914 167023 298942 167051
rect 298728 166961 298756 166989
rect 298790 166961 298818 166989
rect 298852 166961 298880 166989
rect 298914 166961 298942 166989
rect 298728 158147 298756 158175
rect 298790 158147 298818 158175
rect 298852 158147 298880 158175
rect 298914 158147 298942 158175
rect 298728 158085 298756 158113
rect 298790 158085 298818 158113
rect 298852 158085 298880 158113
rect 298914 158085 298942 158113
rect 298728 158023 298756 158051
rect 298790 158023 298818 158051
rect 298852 158023 298880 158051
rect 298914 158023 298942 158051
rect 298728 157961 298756 157989
rect 298790 157961 298818 157989
rect 298852 157961 298880 157989
rect 298914 157961 298942 157989
rect 298728 149147 298756 149175
rect 298790 149147 298818 149175
rect 298852 149147 298880 149175
rect 298914 149147 298942 149175
rect 298728 149085 298756 149113
rect 298790 149085 298818 149113
rect 298852 149085 298880 149113
rect 298914 149085 298942 149113
rect 298728 149023 298756 149051
rect 298790 149023 298818 149051
rect 298852 149023 298880 149051
rect 298914 149023 298942 149051
rect 298728 148961 298756 148989
rect 298790 148961 298818 148989
rect 298852 148961 298880 148989
rect 298914 148961 298942 148989
rect 298728 140147 298756 140175
rect 298790 140147 298818 140175
rect 298852 140147 298880 140175
rect 298914 140147 298942 140175
rect 298728 140085 298756 140113
rect 298790 140085 298818 140113
rect 298852 140085 298880 140113
rect 298914 140085 298942 140113
rect 298728 140023 298756 140051
rect 298790 140023 298818 140051
rect 298852 140023 298880 140051
rect 298914 140023 298942 140051
rect 298728 139961 298756 139989
rect 298790 139961 298818 139989
rect 298852 139961 298880 139989
rect 298914 139961 298942 139989
rect 298728 131147 298756 131175
rect 298790 131147 298818 131175
rect 298852 131147 298880 131175
rect 298914 131147 298942 131175
rect 298728 131085 298756 131113
rect 298790 131085 298818 131113
rect 298852 131085 298880 131113
rect 298914 131085 298942 131113
rect 298728 131023 298756 131051
rect 298790 131023 298818 131051
rect 298852 131023 298880 131051
rect 298914 131023 298942 131051
rect 298728 130961 298756 130989
rect 298790 130961 298818 130989
rect 298852 130961 298880 130989
rect 298914 130961 298942 130989
rect 298728 122147 298756 122175
rect 298790 122147 298818 122175
rect 298852 122147 298880 122175
rect 298914 122147 298942 122175
rect 298728 122085 298756 122113
rect 298790 122085 298818 122113
rect 298852 122085 298880 122113
rect 298914 122085 298942 122113
rect 298728 122023 298756 122051
rect 298790 122023 298818 122051
rect 298852 122023 298880 122051
rect 298914 122023 298942 122051
rect 298728 121961 298756 121989
rect 298790 121961 298818 121989
rect 298852 121961 298880 121989
rect 298914 121961 298942 121989
rect 298728 113147 298756 113175
rect 298790 113147 298818 113175
rect 298852 113147 298880 113175
rect 298914 113147 298942 113175
rect 298728 113085 298756 113113
rect 298790 113085 298818 113113
rect 298852 113085 298880 113113
rect 298914 113085 298942 113113
rect 298728 113023 298756 113051
rect 298790 113023 298818 113051
rect 298852 113023 298880 113051
rect 298914 113023 298942 113051
rect 298728 112961 298756 112989
rect 298790 112961 298818 112989
rect 298852 112961 298880 112989
rect 298914 112961 298942 112989
rect 298728 104147 298756 104175
rect 298790 104147 298818 104175
rect 298852 104147 298880 104175
rect 298914 104147 298942 104175
rect 298728 104085 298756 104113
rect 298790 104085 298818 104113
rect 298852 104085 298880 104113
rect 298914 104085 298942 104113
rect 298728 104023 298756 104051
rect 298790 104023 298818 104051
rect 298852 104023 298880 104051
rect 298914 104023 298942 104051
rect 298728 103961 298756 103989
rect 298790 103961 298818 103989
rect 298852 103961 298880 103989
rect 298914 103961 298942 103989
rect 298728 95147 298756 95175
rect 298790 95147 298818 95175
rect 298852 95147 298880 95175
rect 298914 95147 298942 95175
rect 298728 95085 298756 95113
rect 298790 95085 298818 95113
rect 298852 95085 298880 95113
rect 298914 95085 298942 95113
rect 298728 95023 298756 95051
rect 298790 95023 298818 95051
rect 298852 95023 298880 95051
rect 298914 95023 298942 95051
rect 298728 94961 298756 94989
rect 298790 94961 298818 94989
rect 298852 94961 298880 94989
rect 298914 94961 298942 94989
rect 298728 86147 298756 86175
rect 298790 86147 298818 86175
rect 298852 86147 298880 86175
rect 298914 86147 298942 86175
rect 298728 86085 298756 86113
rect 298790 86085 298818 86113
rect 298852 86085 298880 86113
rect 298914 86085 298942 86113
rect 298728 86023 298756 86051
rect 298790 86023 298818 86051
rect 298852 86023 298880 86051
rect 298914 86023 298942 86051
rect 298728 85961 298756 85989
rect 298790 85961 298818 85989
rect 298852 85961 298880 85989
rect 298914 85961 298942 85989
rect 298728 77147 298756 77175
rect 298790 77147 298818 77175
rect 298852 77147 298880 77175
rect 298914 77147 298942 77175
rect 298728 77085 298756 77113
rect 298790 77085 298818 77113
rect 298852 77085 298880 77113
rect 298914 77085 298942 77113
rect 298728 77023 298756 77051
rect 298790 77023 298818 77051
rect 298852 77023 298880 77051
rect 298914 77023 298942 77051
rect 298728 76961 298756 76989
rect 298790 76961 298818 76989
rect 298852 76961 298880 76989
rect 298914 76961 298942 76989
rect 298728 68147 298756 68175
rect 298790 68147 298818 68175
rect 298852 68147 298880 68175
rect 298914 68147 298942 68175
rect 298728 68085 298756 68113
rect 298790 68085 298818 68113
rect 298852 68085 298880 68113
rect 298914 68085 298942 68113
rect 298728 68023 298756 68051
rect 298790 68023 298818 68051
rect 298852 68023 298880 68051
rect 298914 68023 298942 68051
rect 298728 67961 298756 67989
rect 298790 67961 298818 67989
rect 298852 67961 298880 67989
rect 298914 67961 298942 67989
rect 298728 59147 298756 59175
rect 298790 59147 298818 59175
rect 298852 59147 298880 59175
rect 298914 59147 298942 59175
rect 298728 59085 298756 59113
rect 298790 59085 298818 59113
rect 298852 59085 298880 59113
rect 298914 59085 298942 59113
rect 298728 59023 298756 59051
rect 298790 59023 298818 59051
rect 298852 59023 298880 59051
rect 298914 59023 298942 59051
rect 298728 58961 298756 58989
rect 298790 58961 298818 58989
rect 298852 58961 298880 58989
rect 298914 58961 298942 58989
rect 298728 50147 298756 50175
rect 298790 50147 298818 50175
rect 298852 50147 298880 50175
rect 298914 50147 298942 50175
rect 298728 50085 298756 50113
rect 298790 50085 298818 50113
rect 298852 50085 298880 50113
rect 298914 50085 298942 50113
rect 298728 50023 298756 50051
rect 298790 50023 298818 50051
rect 298852 50023 298880 50051
rect 298914 50023 298942 50051
rect 298728 49961 298756 49989
rect 298790 49961 298818 49989
rect 298852 49961 298880 49989
rect 298914 49961 298942 49989
rect 298728 41147 298756 41175
rect 298790 41147 298818 41175
rect 298852 41147 298880 41175
rect 298914 41147 298942 41175
rect 298728 41085 298756 41113
rect 298790 41085 298818 41113
rect 298852 41085 298880 41113
rect 298914 41085 298942 41113
rect 298728 41023 298756 41051
rect 298790 41023 298818 41051
rect 298852 41023 298880 41051
rect 298914 41023 298942 41051
rect 298728 40961 298756 40989
rect 298790 40961 298818 40989
rect 298852 40961 298880 40989
rect 298914 40961 298942 40989
rect 298728 32147 298756 32175
rect 298790 32147 298818 32175
rect 298852 32147 298880 32175
rect 298914 32147 298942 32175
rect 298728 32085 298756 32113
rect 298790 32085 298818 32113
rect 298852 32085 298880 32113
rect 298914 32085 298942 32113
rect 298728 32023 298756 32051
rect 298790 32023 298818 32051
rect 298852 32023 298880 32051
rect 298914 32023 298942 32051
rect 298728 31961 298756 31989
rect 298790 31961 298818 31989
rect 298852 31961 298880 31989
rect 298914 31961 298942 31989
rect 298728 23147 298756 23175
rect 298790 23147 298818 23175
rect 298852 23147 298880 23175
rect 298914 23147 298942 23175
rect 298728 23085 298756 23113
rect 298790 23085 298818 23113
rect 298852 23085 298880 23113
rect 298914 23085 298942 23113
rect 298728 23023 298756 23051
rect 298790 23023 298818 23051
rect 298852 23023 298880 23051
rect 298914 23023 298942 23051
rect 298728 22961 298756 22989
rect 298790 22961 298818 22989
rect 298852 22961 298880 22989
rect 298914 22961 298942 22989
rect 298728 14147 298756 14175
rect 298790 14147 298818 14175
rect 298852 14147 298880 14175
rect 298914 14147 298942 14175
rect 298728 14085 298756 14113
rect 298790 14085 298818 14113
rect 298852 14085 298880 14113
rect 298914 14085 298942 14113
rect 298728 14023 298756 14051
rect 298790 14023 298818 14051
rect 298852 14023 298880 14051
rect 298914 14023 298942 14051
rect 298728 13961 298756 13989
rect 298790 13961 298818 13989
rect 298852 13961 298880 13989
rect 298914 13961 298942 13989
rect 298728 5147 298756 5175
rect 298790 5147 298818 5175
rect 298852 5147 298880 5175
rect 298914 5147 298942 5175
rect 298728 5085 298756 5113
rect 298790 5085 298818 5113
rect 298852 5085 298880 5113
rect 298914 5085 298942 5113
rect 298728 5023 298756 5051
rect 298790 5023 298818 5051
rect 298852 5023 298880 5051
rect 298914 5023 298942 5051
rect 298728 4961 298756 4989
rect 298790 4961 298818 4989
rect 298852 4961 298880 4989
rect 298914 4961 298942 4989
rect 296457 -588 296485 -560
rect 296519 -588 296547 -560
rect 296581 -588 296609 -560
rect 296643 -588 296671 -560
rect 296457 -650 296485 -622
rect 296519 -650 296547 -622
rect 296581 -650 296609 -622
rect 296643 -650 296671 -622
rect 296457 -712 296485 -684
rect 296519 -712 296547 -684
rect 296581 -712 296609 -684
rect 296643 -712 296671 -684
rect 296457 -774 296485 -746
rect 296519 -774 296547 -746
rect 296581 -774 296609 -746
rect 296643 -774 296671 -746
rect 298728 -588 298756 -560
rect 298790 -588 298818 -560
rect 298852 -588 298880 -560
rect 298914 -588 298942 -560
rect 298728 -650 298756 -622
rect 298790 -650 298818 -622
rect 298852 -650 298880 -622
rect 298914 -650 298942 -622
rect 298728 -712 298756 -684
rect 298790 -712 298818 -684
rect 298852 -712 298880 -684
rect 298914 -712 298942 -684
rect 298728 -774 298756 -746
rect 298790 -774 298818 -746
rect 298852 -774 298880 -746
rect 298914 -774 298942 -746
<< metal5 >>
rect -958 299086 298990 299134
rect -958 299058 -910 299086
rect -882 299058 -848 299086
rect -820 299058 -786 299086
rect -758 299058 -724 299086
rect -696 299058 4617 299086
rect 4645 299058 4679 299086
rect 4707 299058 4741 299086
rect 4769 299058 4803 299086
rect 4831 299058 19977 299086
rect 20005 299058 20039 299086
rect 20067 299058 20101 299086
rect 20129 299058 20163 299086
rect 20191 299058 35337 299086
rect 35365 299058 35399 299086
rect 35427 299058 35461 299086
rect 35489 299058 35523 299086
rect 35551 299058 50697 299086
rect 50725 299058 50759 299086
rect 50787 299058 50821 299086
rect 50849 299058 50883 299086
rect 50911 299058 66057 299086
rect 66085 299058 66119 299086
rect 66147 299058 66181 299086
rect 66209 299058 66243 299086
rect 66271 299058 81417 299086
rect 81445 299058 81479 299086
rect 81507 299058 81541 299086
rect 81569 299058 81603 299086
rect 81631 299058 96777 299086
rect 96805 299058 96839 299086
rect 96867 299058 96901 299086
rect 96929 299058 96963 299086
rect 96991 299058 112137 299086
rect 112165 299058 112199 299086
rect 112227 299058 112261 299086
rect 112289 299058 112323 299086
rect 112351 299058 127497 299086
rect 127525 299058 127559 299086
rect 127587 299058 127621 299086
rect 127649 299058 127683 299086
rect 127711 299058 142857 299086
rect 142885 299058 142919 299086
rect 142947 299058 142981 299086
rect 143009 299058 143043 299086
rect 143071 299058 158217 299086
rect 158245 299058 158279 299086
rect 158307 299058 158341 299086
rect 158369 299058 158403 299086
rect 158431 299058 173577 299086
rect 173605 299058 173639 299086
rect 173667 299058 173701 299086
rect 173729 299058 173763 299086
rect 173791 299058 188937 299086
rect 188965 299058 188999 299086
rect 189027 299058 189061 299086
rect 189089 299058 189123 299086
rect 189151 299058 204297 299086
rect 204325 299058 204359 299086
rect 204387 299058 204421 299086
rect 204449 299058 204483 299086
rect 204511 299058 219657 299086
rect 219685 299058 219719 299086
rect 219747 299058 219781 299086
rect 219809 299058 219843 299086
rect 219871 299058 235017 299086
rect 235045 299058 235079 299086
rect 235107 299058 235141 299086
rect 235169 299058 235203 299086
rect 235231 299058 250377 299086
rect 250405 299058 250439 299086
rect 250467 299058 250501 299086
rect 250529 299058 250563 299086
rect 250591 299058 265737 299086
rect 265765 299058 265799 299086
rect 265827 299058 265861 299086
rect 265889 299058 265923 299086
rect 265951 299058 281097 299086
rect 281125 299058 281159 299086
rect 281187 299058 281221 299086
rect 281249 299058 281283 299086
rect 281311 299058 296457 299086
rect 296485 299058 296519 299086
rect 296547 299058 296581 299086
rect 296609 299058 296643 299086
rect 296671 299058 298728 299086
rect 298756 299058 298790 299086
rect 298818 299058 298852 299086
rect 298880 299058 298914 299086
rect 298942 299058 298990 299086
rect -958 299024 298990 299058
rect -958 298996 -910 299024
rect -882 298996 -848 299024
rect -820 298996 -786 299024
rect -758 298996 -724 299024
rect -696 298996 4617 299024
rect 4645 298996 4679 299024
rect 4707 298996 4741 299024
rect 4769 298996 4803 299024
rect 4831 298996 19977 299024
rect 20005 298996 20039 299024
rect 20067 298996 20101 299024
rect 20129 298996 20163 299024
rect 20191 298996 35337 299024
rect 35365 298996 35399 299024
rect 35427 298996 35461 299024
rect 35489 298996 35523 299024
rect 35551 298996 50697 299024
rect 50725 298996 50759 299024
rect 50787 298996 50821 299024
rect 50849 298996 50883 299024
rect 50911 298996 66057 299024
rect 66085 298996 66119 299024
rect 66147 298996 66181 299024
rect 66209 298996 66243 299024
rect 66271 298996 81417 299024
rect 81445 298996 81479 299024
rect 81507 298996 81541 299024
rect 81569 298996 81603 299024
rect 81631 298996 96777 299024
rect 96805 298996 96839 299024
rect 96867 298996 96901 299024
rect 96929 298996 96963 299024
rect 96991 298996 112137 299024
rect 112165 298996 112199 299024
rect 112227 298996 112261 299024
rect 112289 298996 112323 299024
rect 112351 298996 127497 299024
rect 127525 298996 127559 299024
rect 127587 298996 127621 299024
rect 127649 298996 127683 299024
rect 127711 298996 142857 299024
rect 142885 298996 142919 299024
rect 142947 298996 142981 299024
rect 143009 298996 143043 299024
rect 143071 298996 158217 299024
rect 158245 298996 158279 299024
rect 158307 298996 158341 299024
rect 158369 298996 158403 299024
rect 158431 298996 173577 299024
rect 173605 298996 173639 299024
rect 173667 298996 173701 299024
rect 173729 298996 173763 299024
rect 173791 298996 188937 299024
rect 188965 298996 188999 299024
rect 189027 298996 189061 299024
rect 189089 298996 189123 299024
rect 189151 298996 204297 299024
rect 204325 298996 204359 299024
rect 204387 298996 204421 299024
rect 204449 298996 204483 299024
rect 204511 298996 219657 299024
rect 219685 298996 219719 299024
rect 219747 298996 219781 299024
rect 219809 298996 219843 299024
rect 219871 298996 235017 299024
rect 235045 298996 235079 299024
rect 235107 298996 235141 299024
rect 235169 298996 235203 299024
rect 235231 298996 250377 299024
rect 250405 298996 250439 299024
rect 250467 298996 250501 299024
rect 250529 298996 250563 299024
rect 250591 298996 265737 299024
rect 265765 298996 265799 299024
rect 265827 298996 265861 299024
rect 265889 298996 265923 299024
rect 265951 298996 281097 299024
rect 281125 298996 281159 299024
rect 281187 298996 281221 299024
rect 281249 298996 281283 299024
rect 281311 298996 296457 299024
rect 296485 298996 296519 299024
rect 296547 298996 296581 299024
rect 296609 298996 296643 299024
rect 296671 298996 298728 299024
rect 298756 298996 298790 299024
rect 298818 298996 298852 299024
rect 298880 298996 298914 299024
rect 298942 298996 298990 299024
rect -958 298962 298990 298996
rect -958 298934 -910 298962
rect -882 298934 -848 298962
rect -820 298934 -786 298962
rect -758 298934 -724 298962
rect -696 298934 4617 298962
rect 4645 298934 4679 298962
rect 4707 298934 4741 298962
rect 4769 298934 4803 298962
rect 4831 298934 19977 298962
rect 20005 298934 20039 298962
rect 20067 298934 20101 298962
rect 20129 298934 20163 298962
rect 20191 298934 35337 298962
rect 35365 298934 35399 298962
rect 35427 298934 35461 298962
rect 35489 298934 35523 298962
rect 35551 298934 50697 298962
rect 50725 298934 50759 298962
rect 50787 298934 50821 298962
rect 50849 298934 50883 298962
rect 50911 298934 66057 298962
rect 66085 298934 66119 298962
rect 66147 298934 66181 298962
rect 66209 298934 66243 298962
rect 66271 298934 81417 298962
rect 81445 298934 81479 298962
rect 81507 298934 81541 298962
rect 81569 298934 81603 298962
rect 81631 298934 96777 298962
rect 96805 298934 96839 298962
rect 96867 298934 96901 298962
rect 96929 298934 96963 298962
rect 96991 298934 112137 298962
rect 112165 298934 112199 298962
rect 112227 298934 112261 298962
rect 112289 298934 112323 298962
rect 112351 298934 127497 298962
rect 127525 298934 127559 298962
rect 127587 298934 127621 298962
rect 127649 298934 127683 298962
rect 127711 298934 142857 298962
rect 142885 298934 142919 298962
rect 142947 298934 142981 298962
rect 143009 298934 143043 298962
rect 143071 298934 158217 298962
rect 158245 298934 158279 298962
rect 158307 298934 158341 298962
rect 158369 298934 158403 298962
rect 158431 298934 173577 298962
rect 173605 298934 173639 298962
rect 173667 298934 173701 298962
rect 173729 298934 173763 298962
rect 173791 298934 188937 298962
rect 188965 298934 188999 298962
rect 189027 298934 189061 298962
rect 189089 298934 189123 298962
rect 189151 298934 204297 298962
rect 204325 298934 204359 298962
rect 204387 298934 204421 298962
rect 204449 298934 204483 298962
rect 204511 298934 219657 298962
rect 219685 298934 219719 298962
rect 219747 298934 219781 298962
rect 219809 298934 219843 298962
rect 219871 298934 235017 298962
rect 235045 298934 235079 298962
rect 235107 298934 235141 298962
rect 235169 298934 235203 298962
rect 235231 298934 250377 298962
rect 250405 298934 250439 298962
rect 250467 298934 250501 298962
rect 250529 298934 250563 298962
rect 250591 298934 265737 298962
rect 265765 298934 265799 298962
rect 265827 298934 265861 298962
rect 265889 298934 265923 298962
rect 265951 298934 281097 298962
rect 281125 298934 281159 298962
rect 281187 298934 281221 298962
rect 281249 298934 281283 298962
rect 281311 298934 296457 298962
rect 296485 298934 296519 298962
rect 296547 298934 296581 298962
rect 296609 298934 296643 298962
rect 296671 298934 298728 298962
rect 298756 298934 298790 298962
rect 298818 298934 298852 298962
rect 298880 298934 298914 298962
rect 298942 298934 298990 298962
rect -958 298900 298990 298934
rect -958 298872 -910 298900
rect -882 298872 -848 298900
rect -820 298872 -786 298900
rect -758 298872 -724 298900
rect -696 298872 4617 298900
rect 4645 298872 4679 298900
rect 4707 298872 4741 298900
rect 4769 298872 4803 298900
rect 4831 298872 19977 298900
rect 20005 298872 20039 298900
rect 20067 298872 20101 298900
rect 20129 298872 20163 298900
rect 20191 298872 35337 298900
rect 35365 298872 35399 298900
rect 35427 298872 35461 298900
rect 35489 298872 35523 298900
rect 35551 298872 50697 298900
rect 50725 298872 50759 298900
rect 50787 298872 50821 298900
rect 50849 298872 50883 298900
rect 50911 298872 66057 298900
rect 66085 298872 66119 298900
rect 66147 298872 66181 298900
rect 66209 298872 66243 298900
rect 66271 298872 81417 298900
rect 81445 298872 81479 298900
rect 81507 298872 81541 298900
rect 81569 298872 81603 298900
rect 81631 298872 96777 298900
rect 96805 298872 96839 298900
rect 96867 298872 96901 298900
rect 96929 298872 96963 298900
rect 96991 298872 112137 298900
rect 112165 298872 112199 298900
rect 112227 298872 112261 298900
rect 112289 298872 112323 298900
rect 112351 298872 127497 298900
rect 127525 298872 127559 298900
rect 127587 298872 127621 298900
rect 127649 298872 127683 298900
rect 127711 298872 142857 298900
rect 142885 298872 142919 298900
rect 142947 298872 142981 298900
rect 143009 298872 143043 298900
rect 143071 298872 158217 298900
rect 158245 298872 158279 298900
rect 158307 298872 158341 298900
rect 158369 298872 158403 298900
rect 158431 298872 173577 298900
rect 173605 298872 173639 298900
rect 173667 298872 173701 298900
rect 173729 298872 173763 298900
rect 173791 298872 188937 298900
rect 188965 298872 188999 298900
rect 189027 298872 189061 298900
rect 189089 298872 189123 298900
rect 189151 298872 204297 298900
rect 204325 298872 204359 298900
rect 204387 298872 204421 298900
rect 204449 298872 204483 298900
rect 204511 298872 219657 298900
rect 219685 298872 219719 298900
rect 219747 298872 219781 298900
rect 219809 298872 219843 298900
rect 219871 298872 235017 298900
rect 235045 298872 235079 298900
rect 235107 298872 235141 298900
rect 235169 298872 235203 298900
rect 235231 298872 250377 298900
rect 250405 298872 250439 298900
rect 250467 298872 250501 298900
rect 250529 298872 250563 298900
rect 250591 298872 265737 298900
rect 265765 298872 265799 298900
rect 265827 298872 265861 298900
rect 265889 298872 265923 298900
rect 265951 298872 281097 298900
rect 281125 298872 281159 298900
rect 281187 298872 281221 298900
rect 281249 298872 281283 298900
rect 281311 298872 296457 298900
rect 296485 298872 296519 298900
rect 296547 298872 296581 298900
rect 296609 298872 296643 298900
rect 296671 298872 298728 298900
rect 298756 298872 298790 298900
rect 298818 298872 298852 298900
rect 298880 298872 298914 298900
rect 298942 298872 298990 298900
rect -958 298824 298990 298872
rect -478 298606 298510 298654
rect -478 298578 -430 298606
rect -402 298578 -368 298606
rect -340 298578 -306 298606
rect -278 298578 -244 298606
rect -216 298578 2757 298606
rect 2785 298578 2819 298606
rect 2847 298578 2881 298606
rect 2909 298578 2943 298606
rect 2971 298578 18117 298606
rect 18145 298578 18179 298606
rect 18207 298578 18241 298606
rect 18269 298578 18303 298606
rect 18331 298578 33477 298606
rect 33505 298578 33539 298606
rect 33567 298578 33601 298606
rect 33629 298578 33663 298606
rect 33691 298578 48837 298606
rect 48865 298578 48899 298606
rect 48927 298578 48961 298606
rect 48989 298578 49023 298606
rect 49051 298578 64197 298606
rect 64225 298578 64259 298606
rect 64287 298578 64321 298606
rect 64349 298578 64383 298606
rect 64411 298578 79557 298606
rect 79585 298578 79619 298606
rect 79647 298578 79681 298606
rect 79709 298578 79743 298606
rect 79771 298578 94917 298606
rect 94945 298578 94979 298606
rect 95007 298578 95041 298606
rect 95069 298578 95103 298606
rect 95131 298578 110277 298606
rect 110305 298578 110339 298606
rect 110367 298578 110401 298606
rect 110429 298578 110463 298606
rect 110491 298578 125637 298606
rect 125665 298578 125699 298606
rect 125727 298578 125761 298606
rect 125789 298578 125823 298606
rect 125851 298578 140997 298606
rect 141025 298578 141059 298606
rect 141087 298578 141121 298606
rect 141149 298578 141183 298606
rect 141211 298578 156357 298606
rect 156385 298578 156419 298606
rect 156447 298578 156481 298606
rect 156509 298578 156543 298606
rect 156571 298578 171717 298606
rect 171745 298578 171779 298606
rect 171807 298578 171841 298606
rect 171869 298578 171903 298606
rect 171931 298578 187077 298606
rect 187105 298578 187139 298606
rect 187167 298578 187201 298606
rect 187229 298578 187263 298606
rect 187291 298578 202437 298606
rect 202465 298578 202499 298606
rect 202527 298578 202561 298606
rect 202589 298578 202623 298606
rect 202651 298578 217797 298606
rect 217825 298578 217859 298606
rect 217887 298578 217921 298606
rect 217949 298578 217983 298606
rect 218011 298578 233157 298606
rect 233185 298578 233219 298606
rect 233247 298578 233281 298606
rect 233309 298578 233343 298606
rect 233371 298578 248517 298606
rect 248545 298578 248579 298606
rect 248607 298578 248641 298606
rect 248669 298578 248703 298606
rect 248731 298578 263877 298606
rect 263905 298578 263939 298606
rect 263967 298578 264001 298606
rect 264029 298578 264063 298606
rect 264091 298578 279237 298606
rect 279265 298578 279299 298606
rect 279327 298578 279361 298606
rect 279389 298578 279423 298606
rect 279451 298578 294597 298606
rect 294625 298578 294659 298606
rect 294687 298578 294721 298606
rect 294749 298578 294783 298606
rect 294811 298578 298248 298606
rect 298276 298578 298310 298606
rect 298338 298578 298372 298606
rect 298400 298578 298434 298606
rect 298462 298578 298510 298606
rect -478 298544 298510 298578
rect -478 298516 -430 298544
rect -402 298516 -368 298544
rect -340 298516 -306 298544
rect -278 298516 -244 298544
rect -216 298516 2757 298544
rect 2785 298516 2819 298544
rect 2847 298516 2881 298544
rect 2909 298516 2943 298544
rect 2971 298516 18117 298544
rect 18145 298516 18179 298544
rect 18207 298516 18241 298544
rect 18269 298516 18303 298544
rect 18331 298516 33477 298544
rect 33505 298516 33539 298544
rect 33567 298516 33601 298544
rect 33629 298516 33663 298544
rect 33691 298516 48837 298544
rect 48865 298516 48899 298544
rect 48927 298516 48961 298544
rect 48989 298516 49023 298544
rect 49051 298516 64197 298544
rect 64225 298516 64259 298544
rect 64287 298516 64321 298544
rect 64349 298516 64383 298544
rect 64411 298516 79557 298544
rect 79585 298516 79619 298544
rect 79647 298516 79681 298544
rect 79709 298516 79743 298544
rect 79771 298516 94917 298544
rect 94945 298516 94979 298544
rect 95007 298516 95041 298544
rect 95069 298516 95103 298544
rect 95131 298516 110277 298544
rect 110305 298516 110339 298544
rect 110367 298516 110401 298544
rect 110429 298516 110463 298544
rect 110491 298516 125637 298544
rect 125665 298516 125699 298544
rect 125727 298516 125761 298544
rect 125789 298516 125823 298544
rect 125851 298516 140997 298544
rect 141025 298516 141059 298544
rect 141087 298516 141121 298544
rect 141149 298516 141183 298544
rect 141211 298516 156357 298544
rect 156385 298516 156419 298544
rect 156447 298516 156481 298544
rect 156509 298516 156543 298544
rect 156571 298516 171717 298544
rect 171745 298516 171779 298544
rect 171807 298516 171841 298544
rect 171869 298516 171903 298544
rect 171931 298516 187077 298544
rect 187105 298516 187139 298544
rect 187167 298516 187201 298544
rect 187229 298516 187263 298544
rect 187291 298516 202437 298544
rect 202465 298516 202499 298544
rect 202527 298516 202561 298544
rect 202589 298516 202623 298544
rect 202651 298516 217797 298544
rect 217825 298516 217859 298544
rect 217887 298516 217921 298544
rect 217949 298516 217983 298544
rect 218011 298516 233157 298544
rect 233185 298516 233219 298544
rect 233247 298516 233281 298544
rect 233309 298516 233343 298544
rect 233371 298516 248517 298544
rect 248545 298516 248579 298544
rect 248607 298516 248641 298544
rect 248669 298516 248703 298544
rect 248731 298516 263877 298544
rect 263905 298516 263939 298544
rect 263967 298516 264001 298544
rect 264029 298516 264063 298544
rect 264091 298516 279237 298544
rect 279265 298516 279299 298544
rect 279327 298516 279361 298544
rect 279389 298516 279423 298544
rect 279451 298516 294597 298544
rect 294625 298516 294659 298544
rect 294687 298516 294721 298544
rect 294749 298516 294783 298544
rect 294811 298516 298248 298544
rect 298276 298516 298310 298544
rect 298338 298516 298372 298544
rect 298400 298516 298434 298544
rect 298462 298516 298510 298544
rect -478 298482 298510 298516
rect -478 298454 -430 298482
rect -402 298454 -368 298482
rect -340 298454 -306 298482
rect -278 298454 -244 298482
rect -216 298454 2757 298482
rect 2785 298454 2819 298482
rect 2847 298454 2881 298482
rect 2909 298454 2943 298482
rect 2971 298454 18117 298482
rect 18145 298454 18179 298482
rect 18207 298454 18241 298482
rect 18269 298454 18303 298482
rect 18331 298454 33477 298482
rect 33505 298454 33539 298482
rect 33567 298454 33601 298482
rect 33629 298454 33663 298482
rect 33691 298454 48837 298482
rect 48865 298454 48899 298482
rect 48927 298454 48961 298482
rect 48989 298454 49023 298482
rect 49051 298454 64197 298482
rect 64225 298454 64259 298482
rect 64287 298454 64321 298482
rect 64349 298454 64383 298482
rect 64411 298454 79557 298482
rect 79585 298454 79619 298482
rect 79647 298454 79681 298482
rect 79709 298454 79743 298482
rect 79771 298454 94917 298482
rect 94945 298454 94979 298482
rect 95007 298454 95041 298482
rect 95069 298454 95103 298482
rect 95131 298454 110277 298482
rect 110305 298454 110339 298482
rect 110367 298454 110401 298482
rect 110429 298454 110463 298482
rect 110491 298454 125637 298482
rect 125665 298454 125699 298482
rect 125727 298454 125761 298482
rect 125789 298454 125823 298482
rect 125851 298454 140997 298482
rect 141025 298454 141059 298482
rect 141087 298454 141121 298482
rect 141149 298454 141183 298482
rect 141211 298454 156357 298482
rect 156385 298454 156419 298482
rect 156447 298454 156481 298482
rect 156509 298454 156543 298482
rect 156571 298454 171717 298482
rect 171745 298454 171779 298482
rect 171807 298454 171841 298482
rect 171869 298454 171903 298482
rect 171931 298454 187077 298482
rect 187105 298454 187139 298482
rect 187167 298454 187201 298482
rect 187229 298454 187263 298482
rect 187291 298454 202437 298482
rect 202465 298454 202499 298482
rect 202527 298454 202561 298482
rect 202589 298454 202623 298482
rect 202651 298454 217797 298482
rect 217825 298454 217859 298482
rect 217887 298454 217921 298482
rect 217949 298454 217983 298482
rect 218011 298454 233157 298482
rect 233185 298454 233219 298482
rect 233247 298454 233281 298482
rect 233309 298454 233343 298482
rect 233371 298454 248517 298482
rect 248545 298454 248579 298482
rect 248607 298454 248641 298482
rect 248669 298454 248703 298482
rect 248731 298454 263877 298482
rect 263905 298454 263939 298482
rect 263967 298454 264001 298482
rect 264029 298454 264063 298482
rect 264091 298454 279237 298482
rect 279265 298454 279299 298482
rect 279327 298454 279361 298482
rect 279389 298454 279423 298482
rect 279451 298454 294597 298482
rect 294625 298454 294659 298482
rect 294687 298454 294721 298482
rect 294749 298454 294783 298482
rect 294811 298454 298248 298482
rect 298276 298454 298310 298482
rect 298338 298454 298372 298482
rect 298400 298454 298434 298482
rect 298462 298454 298510 298482
rect -478 298420 298510 298454
rect -478 298392 -430 298420
rect -402 298392 -368 298420
rect -340 298392 -306 298420
rect -278 298392 -244 298420
rect -216 298392 2757 298420
rect 2785 298392 2819 298420
rect 2847 298392 2881 298420
rect 2909 298392 2943 298420
rect 2971 298392 18117 298420
rect 18145 298392 18179 298420
rect 18207 298392 18241 298420
rect 18269 298392 18303 298420
rect 18331 298392 33477 298420
rect 33505 298392 33539 298420
rect 33567 298392 33601 298420
rect 33629 298392 33663 298420
rect 33691 298392 48837 298420
rect 48865 298392 48899 298420
rect 48927 298392 48961 298420
rect 48989 298392 49023 298420
rect 49051 298392 64197 298420
rect 64225 298392 64259 298420
rect 64287 298392 64321 298420
rect 64349 298392 64383 298420
rect 64411 298392 79557 298420
rect 79585 298392 79619 298420
rect 79647 298392 79681 298420
rect 79709 298392 79743 298420
rect 79771 298392 94917 298420
rect 94945 298392 94979 298420
rect 95007 298392 95041 298420
rect 95069 298392 95103 298420
rect 95131 298392 110277 298420
rect 110305 298392 110339 298420
rect 110367 298392 110401 298420
rect 110429 298392 110463 298420
rect 110491 298392 125637 298420
rect 125665 298392 125699 298420
rect 125727 298392 125761 298420
rect 125789 298392 125823 298420
rect 125851 298392 140997 298420
rect 141025 298392 141059 298420
rect 141087 298392 141121 298420
rect 141149 298392 141183 298420
rect 141211 298392 156357 298420
rect 156385 298392 156419 298420
rect 156447 298392 156481 298420
rect 156509 298392 156543 298420
rect 156571 298392 171717 298420
rect 171745 298392 171779 298420
rect 171807 298392 171841 298420
rect 171869 298392 171903 298420
rect 171931 298392 187077 298420
rect 187105 298392 187139 298420
rect 187167 298392 187201 298420
rect 187229 298392 187263 298420
rect 187291 298392 202437 298420
rect 202465 298392 202499 298420
rect 202527 298392 202561 298420
rect 202589 298392 202623 298420
rect 202651 298392 217797 298420
rect 217825 298392 217859 298420
rect 217887 298392 217921 298420
rect 217949 298392 217983 298420
rect 218011 298392 233157 298420
rect 233185 298392 233219 298420
rect 233247 298392 233281 298420
rect 233309 298392 233343 298420
rect 233371 298392 248517 298420
rect 248545 298392 248579 298420
rect 248607 298392 248641 298420
rect 248669 298392 248703 298420
rect 248731 298392 263877 298420
rect 263905 298392 263939 298420
rect 263967 298392 264001 298420
rect 264029 298392 264063 298420
rect 264091 298392 279237 298420
rect 279265 298392 279299 298420
rect 279327 298392 279361 298420
rect 279389 298392 279423 298420
rect 279451 298392 294597 298420
rect 294625 298392 294659 298420
rect 294687 298392 294721 298420
rect 294749 298392 294783 298420
rect 294811 298392 298248 298420
rect 298276 298392 298310 298420
rect 298338 298392 298372 298420
rect 298400 298392 298434 298420
rect 298462 298392 298510 298420
rect -478 298344 298510 298392
rect -958 293175 298990 293223
rect -958 293147 -910 293175
rect -882 293147 -848 293175
rect -820 293147 -786 293175
rect -758 293147 -724 293175
rect -696 293147 4617 293175
rect 4645 293147 4679 293175
rect 4707 293147 4741 293175
rect 4769 293147 4803 293175
rect 4831 293147 19977 293175
rect 20005 293147 20039 293175
rect 20067 293147 20101 293175
rect 20129 293147 20163 293175
rect 20191 293147 35337 293175
rect 35365 293147 35399 293175
rect 35427 293147 35461 293175
rect 35489 293147 35523 293175
rect 35551 293147 50697 293175
rect 50725 293147 50759 293175
rect 50787 293147 50821 293175
rect 50849 293147 50883 293175
rect 50911 293147 66057 293175
rect 66085 293147 66119 293175
rect 66147 293147 66181 293175
rect 66209 293147 66243 293175
rect 66271 293147 81417 293175
rect 81445 293147 81479 293175
rect 81507 293147 81541 293175
rect 81569 293147 81603 293175
rect 81631 293147 96777 293175
rect 96805 293147 96839 293175
rect 96867 293147 96901 293175
rect 96929 293147 96963 293175
rect 96991 293147 112137 293175
rect 112165 293147 112199 293175
rect 112227 293147 112261 293175
rect 112289 293147 112323 293175
rect 112351 293147 127497 293175
rect 127525 293147 127559 293175
rect 127587 293147 127621 293175
rect 127649 293147 127683 293175
rect 127711 293147 142857 293175
rect 142885 293147 142919 293175
rect 142947 293147 142981 293175
rect 143009 293147 143043 293175
rect 143071 293147 158217 293175
rect 158245 293147 158279 293175
rect 158307 293147 158341 293175
rect 158369 293147 158403 293175
rect 158431 293147 173577 293175
rect 173605 293147 173639 293175
rect 173667 293147 173701 293175
rect 173729 293147 173763 293175
rect 173791 293147 188937 293175
rect 188965 293147 188999 293175
rect 189027 293147 189061 293175
rect 189089 293147 189123 293175
rect 189151 293147 204297 293175
rect 204325 293147 204359 293175
rect 204387 293147 204421 293175
rect 204449 293147 204483 293175
rect 204511 293147 219657 293175
rect 219685 293147 219719 293175
rect 219747 293147 219781 293175
rect 219809 293147 219843 293175
rect 219871 293147 235017 293175
rect 235045 293147 235079 293175
rect 235107 293147 235141 293175
rect 235169 293147 235203 293175
rect 235231 293147 250377 293175
rect 250405 293147 250439 293175
rect 250467 293147 250501 293175
rect 250529 293147 250563 293175
rect 250591 293147 265737 293175
rect 265765 293147 265799 293175
rect 265827 293147 265861 293175
rect 265889 293147 265923 293175
rect 265951 293147 281097 293175
rect 281125 293147 281159 293175
rect 281187 293147 281221 293175
rect 281249 293147 281283 293175
rect 281311 293147 296457 293175
rect 296485 293147 296519 293175
rect 296547 293147 296581 293175
rect 296609 293147 296643 293175
rect 296671 293147 298728 293175
rect 298756 293147 298790 293175
rect 298818 293147 298852 293175
rect 298880 293147 298914 293175
rect 298942 293147 298990 293175
rect -958 293113 298990 293147
rect -958 293085 -910 293113
rect -882 293085 -848 293113
rect -820 293085 -786 293113
rect -758 293085 -724 293113
rect -696 293085 4617 293113
rect 4645 293085 4679 293113
rect 4707 293085 4741 293113
rect 4769 293085 4803 293113
rect 4831 293085 19977 293113
rect 20005 293085 20039 293113
rect 20067 293085 20101 293113
rect 20129 293085 20163 293113
rect 20191 293085 35337 293113
rect 35365 293085 35399 293113
rect 35427 293085 35461 293113
rect 35489 293085 35523 293113
rect 35551 293085 50697 293113
rect 50725 293085 50759 293113
rect 50787 293085 50821 293113
rect 50849 293085 50883 293113
rect 50911 293085 66057 293113
rect 66085 293085 66119 293113
rect 66147 293085 66181 293113
rect 66209 293085 66243 293113
rect 66271 293085 81417 293113
rect 81445 293085 81479 293113
rect 81507 293085 81541 293113
rect 81569 293085 81603 293113
rect 81631 293085 96777 293113
rect 96805 293085 96839 293113
rect 96867 293085 96901 293113
rect 96929 293085 96963 293113
rect 96991 293085 112137 293113
rect 112165 293085 112199 293113
rect 112227 293085 112261 293113
rect 112289 293085 112323 293113
rect 112351 293085 127497 293113
rect 127525 293085 127559 293113
rect 127587 293085 127621 293113
rect 127649 293085 127683 293113
rect 127711 293085 142857 293113
rect 142885 293085 142919 293113
rect 142947 293085 142981 293113
rect 143009 293085 143043 293113
rect 143071 293085 158217 293113
rect 158245 293085 158279 293113
rect 158307 293085 158341 293113
rect 158369 293085 158403 293113
rect 158431 293085 173577 293113
rect 173605 293085 173639 293113
rect 173667 293085 173701 293113
rect 173729 293085 173763 293113
rect 173791 293085 188937 293113
rect 188965 293085 188999 293113
rect 189027 293085 189061 293113
rect 189089 293085 189123 293113
rect 189151 293085 204297 293113
rect 204325 293085 204359 293113
rect 204387 293085 204421 293113
rect 204449 293085 204483 293113
rect 204511 293085 219657 293113
rect 219685 293085 219719 293113
rect 219747 293085 219781 293113
rect 219809 293085 219843 293113
rect 219871 293085 235017 293113
rect 235045 293085 235079 293113
rect 235107 293085 235141 293113
rect 235169 293085 235203 293113
rect 235231 293085 250377 293113
rect 250405 293085 250439 293113
rect 250467 293085 250501 293113
rect 250529 293085 250563 293113
rect 250591 293085 265737 293113
rect 265765 293085 265799 293113
rect 265827 293085 265861 293113
rect 265889 293085 265923 293113
rect 265951 293085 281097 293113
rect 281125 293085 281159 293113
rect 281187 293085 281221 293113
rect 281249 293085 281283 293113
rect 281311 293085 296457 293113
rect 296485 293085 296519 293113
rect 296547 293085 296581 293113
rect 296609 293085 296643 293113
rect 296671 293085 298728 293113
rect 298756 293085 298790 293113
rect 298818 293085 298852 293113
rect 298880 293085 298914 293113
rect 298942 293085 298990 293113
rect -958 293051 298990 293085
rect -958 293023 -910 293051
rect -882 293023 -848 293051
rect -820 293023 -786 293051
rect -758 293023 -724 293051
rect -696 293023 4617 293051
rect 4645 293023 4679 293051
rect 4707 293023 4741 293051
rect 4769 293023 4803 293051
rect 4831 293023 19977 293051
rect 20005 293023 20039 293051
rect 20067 293023 20101 293051
rect 20129 293023 20163 293051
rect 20191 293023 35337 293051
rect 35365 293023 35399 293051
rect 35427 293023 35461 293051
rect 35489 293023 35523 293051
rect 35551 293023 50697 293051
rect 50725 293023 50759 293051
rect 50787 293023 50821 293051
rect 50849 293023 50883 293051
rect 50911 293023 66057 293051
rect 66085 293023 66119 293051
rect 66147 293023 66181 293051
rect 66209 293023 66243 293051
rect 66271 293023 81417 293051
rect 81445 293023 81479 293051
rect 81507 293023 81541 293051
rect 81569 293023 81603 293051
rect 81631 293023 96777 293051
rect 96805 293023 96839 293051
rect 96867 293023 96901 293051
rect 96929 293023 96963 293051
rect 96991 293023 112137 293051
rect 112165 293023 112199 293051
rect 112227 293023 112261 293051
rect 112289 293023 112323 293051
rect 112351 293023 127497 293051
rect 127525 293023 127559 293051
rect 127587 293023 127621 293051
rect 127649 293023 127683 293051
rect 127711 293023 142857 293051
rect 142885 293023 142919 293051
rect 142947 293023 142981 293051
rect 143009 293023 143043 293051
rect 143071 293023 158217 293051
rect 158245 293023 158279 293051
rect 158307 293023 158341 293051
rect 158369 293023 158403 293051
rect 158431 293023 173577 293051
rect 173605 293023 173639 293051
rect 173667 293023 173701 293051
rect 173729 293023 173763 293051
rect 173791 293023 188937 293051
rect 188965 293023 188999 293051
rect 189027 293023 189061 293051
rect 189089 293023 189123 293051
rect 189151 293023 204297 293051
rect 204325 293023 204359 293051
rect 204387 293023 204421 293051
rect 204449 293023 204483 293051
rect 204511 293023 219657 293051
rect 219685 293023 219719 293051
rect 219747 293023 219781 293051
rect 219809 293023 219843 293051
rect 219871 293023 235017 293051
rect 235045 293023 235079 293051
rect 235107 293023 235141 293051
rect 235169 293023 235203 293051
rect 235231 293023 250377 293051
rect 250405 293023 250439 293051
rect 250467 293023 250501 293051
rect 250529 293023 250563 293051
rect 250591 293023 265737 293051
rect 265765 293023 265799 293051
rect 265827 293023 265861 293051
rect 265889 293023 265923 293051
rect 265951 293023 281097 293051
rect 281125 293023 281159 293051
rect 281187 293023 281221 293051
rect 281249 293023 281283 293051
rect 281311 293023 296457 293051
rect 296485 293023 296519 293051
rect 296547 293023 296581 293051
rect 296609 293023 296643 293051
rect 296671 293023 298728 293051
rect 298756 293023 298790 293051
rect 298818 293023 298852 293051
rect 298880 293023 298914 293051
rect 298942 293023 298990 293051
rect -958 292989 298990 293023
rect -958 292961 -910 292989
rect -882 292961 -848 292989
rect -820 292961 -786 292989
rect -758 292961 -724 292989
rect -696 292961 4617 292989
rect 4645 292961 4679 292989
rect 4707 292961 4741 292989
rect 4769 292961 4803 292989
rect 4831 292961 19977 292989
rect 20005 292961 20039 292989
rect 20067 292961 20101 292989
rect 20129 292961 20163 292989
rect 20191 292961 35337 292989
rect 35365 292961 35399 292989
rect 35427 292961 35461 292989
rect 35489 292961 35523 292989
rect 35551 292961 50697 292989
rect 50725 292961 50759 292989
rect 50787 292961 50821 292989
rect 50849 292961 50883 292989
rect 50911 292961 66057 292989
rect 66085 292961 66119 292989
rect 66147 292961 66181 292989
rect 66209 292961 66243 292989
rect 66271 292961 81417 292989
rect 81445 292961 81479 292989
rect 81507 292961 81541 292989
rect 81569 292961 81603 292989
rect 81631 292961 96777 292989
rect 96805 292961 96839 292989
rect 96867 292961 96901 292989
rect 96929 292961 96963 292989
rect 96991 292961 112137 292989
rect 112165 292961 112199 292989
rect 112227 292961 112261 292989
rect 112289 292961 112323 292989
rect 112351 292961 127497 292989
rect 127525 292961 127559 292989
rect 127587 292961 127621 292989
rect 127649 292961 127683 292989
rect 127711 292961 142857 292989
rect 142885 292961 142919 292989
rect 142947 292961 142981 292989
rect 143009 292961 143043 292989
rect 143071 292961 158217 292989
rect 158245 292961 158279 292989
rect 158307 292961 158341 292989
rect 158369 292961 158403 292989
rect 158431 292961 173577 292989
rect 173605 292961 173639 292989
rect 173667 292961 173701 292989
rect 173729 292961 173763 292989
rect 173791 292961 188937 292989
rect 188965 292961 188999 292989
rect 189027 292961 189061 292989
rect 189089 292961 189123 292989
rect 189151 292961 204297 292989
rect 204325 292961 204359 292989
rect 204387 292961 204421 292989
rect 204449 292961 204483 292989
rect 204511 292961 219657 292989
rect 219685 292961 219719 292989
rect 219747 292961 219781 292989
rect 219809 292961 219843 292989
rect 219871 292961 235017 292989
rect 235045 292961 235079 292989
rect 235107 292961 235141 292989
rect 235169 292961 235203 292989
rect 235231 292961 250377 292989
rect 250405 292961 250439 292989
rect 250467 292961 250501 292989
rect 250529 292961 250563 292989
rect 250591 292961 265737 292989
rect 265765 292961 265799 292989
rect 265827 292961 265861 292989
rect 265889 292961 265923 292989
rect 265951 292961 281097 292989
rect 281125 292961 281159 292989
rect 281187 292961 281221 292989
rect 281249 292961 281283 292989
rect 281311 292961 296457 292989
rect 296485 292961 296519 292989
rect 296547 292961 296581 292989
rect 296609 292961 296643 292989
rect 296671 292961 298728 292989
rect 298756 292961 298790 292989
rect 298818 292961 298852 292989
rect 298880 292961 298914 292989
rect 298942 292961 298990 292989
rect -958 292913 298990 292961
rect -958 290175 298990 290223
rect -958 290147 -430 290175
rect -402 290147 -368 290175
rect -340 290147 -306 290175
rect -278 290147 -244 290175
rect -216 290147 2757 290175
rect 2785 290147 2819 290175
rect 2847 290147 2881 290175
rect 2909 290147 2943 290175
rect 2971 290147 18117 290175
rect 18145 290147 18179 290175
rect 18207 290147 18241 290175
rect 18269 290147 18303 290175
rect 18331 290147 33477 290175
rect 33505 290147 33539 290175
rect 33567 290147 33601 290175
rect 33629 290147 33663 290175
rect 33691 290147 48837 290175
rect 48865 290147 48899 290175
rect 48927 290147 48961 290175
rect 48989 290147 49023 290175
rect 49051 290147 64197 290175
rect 64225 290147 64259 290175
rect 64287 290147 64321 290175
rect 64349 290147 64383 290175
rect 64411 290147 79557 290175
rect 79585 290147 79619 290175
rect 79647 290147 79681 290175
rect 79709 290147 79743 290175
rect 79771 290147 94917 290175
rect 94945 290147 94979 290175
rect 95007 290147 95041 290175
rect 95069 290147 95103 290175
rect 95131 290147 110277 290175
rect 110305 290147 110339 290175
rect 110367 290147 110401 290175
rect 110429 290147 110463 290175
rect 110491 290147 125637 290175
rect 125665 290147 125699 290175
rect 125727 290147 125761 290175
rect 125789 290147 125823 290175
rect 125851 290147 140997 290175
rect 141025 290147 141059 290175
rect 141087 290147 141121 290175
rect 141149 290147 141183 290175
rect 141211 290147 156357 290175
rect 156385 290147 156419 290175
rect 156447 290147 156481 290175
rect 156509 290147 156543 290175
rect 156571 290147 171717 290175
rect 171745 290147 171779 290175
rect 171807 290147 171841 290175
rect 171869 290147 171903 290175
rect 171931 290147 187077 290175
rect 187105 290147 187139 290175
rect 187167 290147 187201 290175
rect 187229 290147 187263 290175
rect 187291 290147 202437 290175
rect 202465 290147 202499 290175
rect 202527 290147 202561 290175
rect 202589 290147 202623 290175
rect 202651 290147 217797 290175
rect 217825 290147 217859 290175
rect 217887 290147 217921 290175
rect 217949 290147 217983 290175
rect 218011 290147 233157 290175
rect 233185 290147 233219 290175
rect 233247 290147 233281 290175
rect 233309 290147 233343 290175
rect 233371 290147 248517 290175
rect 248545 290147 248579 290175
rect 248607 290147 248641 290175
rect 248669 290147 248703 290175
rect 248731 290147 263877 290175
rect 263905 290147 263939 290175
rect 263967 290147 264001 290175
rect 264029 290147 264063 290175
rect 264091 290147 279237 290175
rect 279265 290147 279299 290175
rect 279327 290147 279361 290175
rect 279389 290147 279423 290175
rect 279451 290147 294597 290175
rect 294625 290147 294659 290175
rect 294687 290147 294721 290175
rect 294749 290147 294783 290175
rect 294811 290147 298248 290175
rect 298276 290147 298310 290175
rect 298338 290147 298372 290175
rect 298400 290147 298434 290175
rect 298462 290147 298990 290175
rect -958 290113 298990 290147
rect -958 290085 -430 290113
rect -402 290085 -368 290113
rect -340 290085 -306 290113
rect -278 290085 -244 290113
rect -216 290085 2757 290113
rect 2785 290085 2819 290113
rect 2847 290085 2881 290113
rect 2909 290085 2943 290113
rect 2971 290085 18117 290113
rect 18145 290085 18179 290113
rect 18207 290085 18241 290113
rect 18269 290085 18303 290113
rect 18331 290085 33477 290113
rect 33505 290085 33539 290113
rect 33567 290085 33601 290113
rect 33629 290085 33663 290113
rect 33691 290085 48837 290113
rect 48865 290085 48899 290113
rect 48927 290085 48961 290113
rect 48989 290085 49023 290113
rect 49051 290085 64197 290113
rect 64225 290085 64259 290113
rect 64287 290085 64321 290113
rect 64349 290085 64383 290113
rect 64411 290085 79557 290113
rect 79585 290085 79619 290113
rect 79647 290085 79681 290113
rect 79709 290085 79743 290113
rect 79771 290085 94917 290113
rect 94945 290085 94979 290113
rect 95007 290085 95041 290113
rect 95069 290085 95103 290113
rect 95131 290085 110277 290113
rect 110305 290085 110339 290113
rect 110367 290085 110401 290113
rect 110429 290085 110463 290113
rect 110491 290085 125637 290113
rect 125665 290085 125699 290113
rect 125727 290085 125761 290113
rect 125789 290085 125823 290113
rect 125851 290085 140997 290113
rect 141025 290085 141059 290113
rect 141087 290085 141121 290113
rect 141149 290085 141183 290113
rect 141211 290085 156357 290113
rect 156385 290085 156419 290113
rect 156447 290085 156481 290113
rect 156509 290085 156543 290113
rect 156571 290085 171717 290113
rect 171745 290085 171779 290113
rect 171807 290085 171841 290113
rect 171869 290085 171903 290113
rect 171931 290085 187077 290113
rect 187105 290085 187139 290113
rect 187167 290085 187201 290113
rect 187229 290085 187263 290113
rect 187291 290085 202437 290113
rect 202465 290085 202499 290113
rect 202527 290085 202561 290113
rect 202589 290085 202623 290113
rect 202651 290085 217797 290113
rect 217825 290085 217859 290113
rect 217887 290085 217921 290113
rect 217949 290085 217983 290113
rect 218011 290085 233157 290113
rect 233185 290085 233219 290113
rect 233247 290085 233281 290113
rect 233309 290085 233343 290113
rect 233371 290085 248517 290113
rect 248545 290085 248579 290113
rect 248607 290085 248641 290113
rect 248669 290085 248703 290113
rect 248731 290085 263877 290113
rect 263905 290085 263939 290113
rect 263967 290085 264001 290113
rect 264029 290085 264063 290113
rect 264091 290085 279237 290113
rect 279265 290085 279299 290113
rect 279327 290085 279361 290113
rect 279389 290085 279423 290113
rect 279451 290085 294597 290113
rect 294625 290085 294659 290113
rect 294687 290085 294721 290113
rect 294749 290085 294783 290113
rect 294811 290085 298248 290113
rect 298276 290085 298310 290113
rect 298338 290085 298372 290113
rect 298400 290085 298434 290113
rect 298462 290085 298990 290113
rect -958 290051 298990 290085
rect -958 290023 -430 290051
rect -402 290023 -368 290051
rect -340 290023 -306 290051
rect -278 290023 -244 290051
rect -216 290023 2757 290051
rect 2785 290023 2819 290051
rect 2847 290023 2881 290051
rect 2909 290023 2943 290051
rect 2971 290023 18117 290051
rect 18145 290023 18179 290051
rect 18207 290023 18241 290051
rect 18269 290023 18303 290051
rect 18331 290023 33477 290051
rect 33505 290023 33539 290051
rect 33567 290023 33601 290051
rect 33629 290023 33663 290051
rect 33691 290023 48837 290051
rect 48865 290023 48899 290051
rect 48927 290023 48961 290051
rect 48989 290023 49023 290051
rect 49051 290023 64197 290051
rect 64225 290023 64259 290051
rect 64287 290023 64321 290051
rect 64349 290023 64383 290051
rect 64411 290023 79557 290051
rect 79585 290023 79619 290051
rect 79647 290023 79681 290051
rect 79709 290023 79743 290051
rect 79771 290023 94917 290051
rect 94945 290023 94979 290051
rect 95007 290023 95041 290051
rect 95069 290023 95103 290051
rect 95131 290023 110277 290051
rect 110305 290023 110339 290051
rect 110367 290023 110401 290051
rect 110429 290023 110463 290051
rect 110491 290023 125637 290051
rect 125665 290023 125699 290051
rect 125727 290023 125761 290051
rect 125789 290023 125823 290051
rect 125851 290023 140997 290051
rect 141025 290023 141059 290051
rect 141087 290023 141121 290051
rect 141149 290023 141183 290051
rect 141211 290023 156357 290051
rect 156385 290023 156419 290051
rect 156447 290023 156481 290051
rect 156509 290023 156543 290051
rect 156571 290023 171717 290051
rect 171745 290023 171779 290051
rect 171807 290023 171841 290051
rect 171869 290023 171903 290051
rect 171931 290023 187077 290051
rect 187105 290023 187139 290051
rect 187167 290023 187201 290051
rect 187229 290023 187263 290051
rect 187291 290023 202437 290051
rect 202465 290023 202499 290051
rect 202527 290023 202561 290051
rect 202589 290023 202623 290051
rect 202651 290023 217797 290051
rect 217825 290023 217859 290051
rect 217887 290023 217921 290051
rect 217949 290023 217983 290051
rect 218011 290023 233157 290051
rect 233185 290023 233219 290051
rect 233247 290023 233281 290051
rect 233309 290023 233343 290051
rect 233371 290023 248517 290051
rect 248545 290023 248579 290051
rect 248607 290023 248641 290051
rect 248669 290023 248703 290051
rect 248731 290023 263877 290051
rect 263905 290023 263939 290051
rect 263967 290023 264001 290051
rect 264029 290023 264063 290051
rect 264091 290023 279237 290051
rect 279265 290023 279299 290051
rect 279327 290023 279361 290051
rect 279389 290023 279423 290051
rect 279451 290023 294597 290051
rect 294625 290023 294659 290051
rect 294687 290023 294721 290051
rect 294749 290023 294783 290051
rect 294811 290023 298248 290051
rect 298276 290023 298310 290051
rect 298338 290023 298372 290051
rect 298400 290023 298434 290051
rect 298462 290023 298990 290051
rect -958 289989 298990 290023
rect -958 289961 -430 289989
rect -402 289961 -368 289989
rect -340 289961 -306 289989
rect -278 289961 -244 289989
rect -216 289961 2757 289989
rect 2785 289961 2819 289989
rect 2847 289961 2881 289989
rect 2909 289961 2943 289989
rect 2971 289961 18117 289989
rect 18145 289961 18179 289989
rect 18207 289961 18241 289989
rect 18269 289961 18303 289989
rect 18331 289961 33477 289989
rect 33505 289961 33539 289989
rect 33567 289961 33601 289989
rect 33629 289961 33663 289989
rect 33691 289961 48837 289989
rect 48865 289961 48899 289989
rect 48927 289961 48961 289989
rect 48989 289961 49023 289989
rect 49051 289961 64197 289989
rect 64225 289961 64259 289989
rect 64287 289961 64321 289989
rect 64349 289961 64383 289989
rect 64411 289961 79557 289989
rect 79585 289961 79619 289989
rect 79647 289961 79681 289989
rect 79709 289961 79743 289989
rect 79771 289961 94917 289989
rect 94945 289961 94979 289989
rect 95007 289961 95041 289989
rect 95069 289961 95103 289989
rect 95131 289961 110277 289989
rect 110305 289961 110339 289989
rect 110367 289961 110401 289989
rect 110429 289961 110463 289989
rect 110491 289961 125637 289989
rect 125665 289961 125699 289989
rect 125727 289961 125761 289989
rect 125789 289961 125823 289989
rect 125851 289961 140997 289989
rect 141025 289961 141059 289989
rect 141087 289961 141121 289989
rect 141149 289961 141183 289989
rect 141211 289961 156357 289989
rect 156385 289961 156419 289989
rect 156447 289961 156481 289989
rect 156509 289961 156543 289989
rect 156571 289961 171717 289989
rect 171745 289961 171779 289989
rect 171807 289961 171841 289989
rect 171869 289961 171903 289989
rect 171931 289961 187077 289989
rect 187105 289961 187139 289989
rect 187167 289961 187201 289989
rect 187229 289961 187263 289989
rect 187291 289961 202437 289989
rect 202465 289961 202499 289989
rect 202527 289961 202561 289989
rect 202589 289961 202623 289989
rect 202651 289961 217797 289989
rect 217825 289961 217859 289989
rect 217887 289961 217921 289989
rect 217949 289961 217983 289989
rect 218011 289961 233157 289989
rect 233185 289961 233219 289989
rect 233247 289961 233281 289989
rect 233309 289961 233343 289989
rect 233371 289961 248517 289989
rect 248545 289961 248579 289989
rect 248607 289961 248641 289989
rect 248669 289961 248703 289989
rect 248731 289961 263877 289989
rect 263905 289961 263939 289989
rect 263967 289961 264001 289989
rect 264029 289961 264063 289989
rect 264091 289961 279237 289989
rect 279265 289961 279299 289989
rect 279327 289961 279361 289989
rect 279389 289961 279423 289989
rect 279451 289961 294597 289989
rect 294625 289961 294659 289989
rect 294687 289961 294721 289989
rect 294749 289961 294783 289989
rect 294811 289961 298248 289989
rect 298276 289961 298310 289989
rect 298338 289961 298372 289989
rect 298400 289961 298434 289989
rect 298462 289961 298990 289989
rect -958 289913 298990 289961
rect -958 284175 298990 284223
rect -958 284147 -910 284175
rect -882 284147 -848 284175
rect -820 284147 -786 284175
rect -758 284147 -724 284175
rect -696 284147 4617 284175
rect 4645 284147 4679 284175
rect 4707 284147 4741 284175
rect 4769 284147 4803 284175
rect 4831 284147 19977 284175
rect 20005 284147 20039 284175
rect 20067 284147 20101 284175
rect 20129 284147 20163 284175
rect 20191 284147 35337 284175
rect 35365 284147 35399 284175
rect 35427 284147 35461 284175
rect 35489 284147 35523 284175
rect 35551 284147 50697 284175
rect 50725 284147 50759 284175
rect 50787 284147 50821 284175
rect 50849 284147 50883 284175
rect 50911 284147 66057 284175
rect 66085 284147 66119 284175
rect 66147 284147 66181 284175
rect 66209 284147 66243 284175
rect 66271 284147 81417 284175
rect 81445 284147 81479 284175
rect 81507 284147 81541 284175
rect 81569 284147 81603 284175
rect 81631 284147 96777 284175
rect 96805 284147 96839 284175
rect 96867 284147 96901 284175
rect 96929 284147 96963 284175
rect 96991 284147 112137 284175
rect 112165 284147 112199 284175
rect 112227 284147 112261 284175
rect 112289 284147 112323 284175
rect 112351 284147 127497 284175
rect 127525 284147 127559 284175
rect 127587 284147 127621 284175
rect 127649 284147 127683 284175
rect 127711 284147 142857 284175
rect 142885 284147 142919 284175
rect 142947 284147 142981 284175
rect 143009 284147 143043 284175
rect 143071 284147 158217 284175
rect 158245 284147 158279 284175
rect 158307 284147 158341 284175
rect 158369 284147 158403 284175
rect 158431 284147 173577 284175
rect 173605 284147 173639 284175
rect 173667 284147 173701 284175
rect 173729 284147 173763 284175
rect 173791 284147 188937 284175
rect 188965 284147 188999 284175
rect 189027 284147 189061 284175
rect 189089 284147 189123 284175
rect 189151 284147 204297 284175
rect 204325 284147 204359 284175
rect 204387 284147 204421 284175
rect 204449 284147 204483 284175
rect 204511 284147 219657 284175
rect 219685 284147 219719 284175
rect 219747 284147 219781 284175
rect 219809 284147 219843 284175
rect 219871 284147 235017 284175
rect 235045 284147 235079 284175
rect 235107 284147 235141 284175
rect 235169 284147 235203 284175
rect 235231 284147 250377 284175
rect 250405 284147 250439 284175
rect 250467 284147 250501 284175
rect 250529 284147 250563 284175
rect 250591 284147 265737 284175
rect 265765 284147 265799 284175
rect 265827 284147 265861 284175
rect 265889 284147 265923 284175
rect 265951 284147 281097 284175
rect 281125 284147 281159 284175
rect 281187 284147 281221 284175
rect 281249 284147 281283 284175
rect 281311 284147 296457 284175
rect 296485 284147 296519 284175
rect 296547 284147 296581 284175
rect 296609 284147 296643 284175
rect 296671 284147 298728 284175
rect 298756 284147 298790 284175
rect 298818 284147 298852 284175
rect 298880 284147 298914 284175
rect 298942 284147 298990 284175
rect -958 284113 298990 284147
rect -958 284085 -910 284113
rect -882 284085 -848 284113
rect -820 284085 -786 284113
rect -758 284085 -724 284113
rect -696 284085 4617 284113
rect 4645 284085 4679 284113
rect 4707 284085 4741 284113
rect 4769 284085 4803 284113
rect 4831 284085 19977 284113
rect 20005 284085 20039 284113
rect 20067 284085 20101 284113
rect 20129 284085 20163 284113
rect 20191 284085 35337 284113
rect 35365 284085 35399 284113
rect 35427 284085 35461 284113
rect 35489 284085 35523 284113
rect 35551 284085 50697 284113
rect 50725 284085 50759 284113
rect 50787 284085 50821 284113
rect 50849 284085 50883 284113
rect 50911 284085 66057 284113
rect 66085 284085 66119 284113
rect 66147 284085 66181 284113
rect 66209 284085 66243 284113
rect 66271 284085 81417 284113
rect 81445 284085 81479 284113
rect 81507 284085 81541 284113
rect 81569 284085 81603 284113
rect 81631 284085 96777 284113
rect 96805 284085 96839 284113
rect 96867 284085 96901 284113
rect 96929 284085 96963 284113
rect 96991 284085 112137 284113
rect 112165 284085 112199 284113
rect 112227 284085 112261 284113
rect 112289 284085 112323 284113
rect 112351 284085 127497 284113
rect 127525 284085 127559 284113
rect 127587 284085 127621 284113
rect 127649 284085 127683 284113
rect 127711 284085 142857 284113
rect 142885 284085 142919 284113
rect 142947 284085 142981 284113
rect 143009 284085 143043 284113
rect 143071 284085 158217 284113
rect 158245 284085 158279 284113
rect 158307 284085 158341 284113
rect 158369 284085 158403 284113
rect 158431 284085 173577 284113
rect 173605 284085 173639 284113
rect 173667 284085 173701 284113
rect 173729 284085 173763 284113
rect 173791 284085 188937 284113
rect 188965 284085 188999 284113
rect 189027 284085 189061 284113
rect 189089 284085 189123 284113
rect 189151 284085 204297 284113
rect 204325 284085 204359 284113
rect 204387 284085 204421 284113
rect 204449 284085 204483 284113
rect 204511 284085 219657 284113
rect 219685 284085 219719 284113
rect 219747 284085 219781 284113
rect 219809 284085 219843 284113
rect 219871 284085 235017 284113
rect 235045 284085 235079 284113
rect 235107 284085 235141 284113
rect 235169 284085 235203 284113
rect 235231 284085 250377 284113
rect 250405 284085 250439 284113
rect 250467 284085 250501 284113
rect 250529 284085 250563 284113
rect 250591 284085 265737 284113
rect 265765 284085 265799 284113
rect 265827 284085 265861 284113
rect 265889 284085 265923 284113
rect 265951 284085 281097 284113
rect 281125 284085 281159 284113
rect 281187 284085 281221 284113
rect 281249 284085 281283 284113
rect 281311 284085 296457 284113
rect 296485 284085 296519 284113
rect 296547 284085 296581 284113
rect 296609 284085 296643 284113
rect 296671 284085 298728 284113
rect 298756 284085 298790 284113
rect 298818 284085 298852 284113
rect 298880 284085 298914 284113
rect 298942 284085 298990 284113
rect -958 284051 298990 284085
rect -958 284023 -910 284051
rect -882 284023 -848 284051
rect -820 284023 -786 284051
rect -758 284023 -724 284051
rect -696 284023 4617 284051
rect 4645 284023 4679 284051
rect 4707 284023 4741 284051
rect 4769 284023 4803 284051
rect 4831 284023 19977 284051
rect 20005 284023 20039 284051
rect 20067 284023 20101 284051
rect 20129 284023 20163 284051
rect 20191 284023 35337 284051
rect 35365 284023 35399 284051
rect 35427 284023 35461 284051
rect 35489 284023 35523 284051
rect 35551 284023 50697 284051
rect 50725 284023 50759 284051
rect 50787 284023 50821 284051
rect 50849 284023 50883 284051
rect 50911 284023 66057 284051
rect 66085 284023 66119 284051
rect 66147 284023 66181 284051
rect 66209 284023 66243 284051
rect 66271 284023 81417 284051
rect 81445 284023 81479 284051
rect 81507 284023 81541 284051
rect 81569 284023 81603 284051
rect 81631 284023 96777 284051
rect 96805 284023 96839 284051
rect 96867 284023 96901 284051
rect 96929 284023 96963 284051
rect 96991 284023 112137 284051
rect 112165 284023 112199 284051
rect 112227 284023 112261 284051
rect 112289 284023 112323 284051
rect 112351 284023 127497 284051
rect 127525 284023 127559 284051
rect 127587 284023 127621 284051
rect 127649 284023 127683 284051
rect 127711 284023 142857 284051
rect 142885 284023 142919 284051
rect 142947 284023 142981 284051
rect 143009 284023 143043 284051
rect 143071 284023 158217 284051
rect 158245 284023 158279 284051
rect 158307 284023 158341 284051
rect 158369 284023 158403 284051
rect 158431 284023 173577 284051
rect 173605 284023 173639 284051
rect 173667 284023 173701 284051
rect 173729 284023 173763 284051
rect 173791 284023 188937 284051
rect 188965 284023 188999 284051
rect 189027 284023 189061 284051
rect 189089 284023 189123 284051
rect 189151 284023 204297 284051
rect 204325 284023 204359 284051
rect 204387 284023 204421 284051
rect 204449 284023 204483 284051
rect 204511 284023 219657 284051
rect 219685 284023 219719 284051
rect 219747 284023 219781 284051
rect 219809 284023 219843 284051
rect 219871 284023 235017 284051
rect 235045 284023 235079 284051
rect 235107 284023 235141 284051
rect 235169 284023 235203 284051
rect 235231 284023 250377 284051
rect 250405 284023 250439 284051
rect 250467 284023 250501 284051
rect 250529 284023 250563 284051
rect 250591 284023 265737 284051
rect 265765 284023 265799 284051
rect 265827 284023 265861 284051
rect 265889 284023 265923 284051
rect 265951 284023 281097 284051
rect 281125 284023 281159 284051
rect 281187 284023 281221 284051
rect 281249 284023 281283 284051
rect 281311 284023 296457 284051
rect 296485 284023 296519 284051
rect 296547 284023 296581 284051
rect 296609 284023 296643 284051
rect 296671 284023 298728 284051
rect 298756 284023 298790 284051
rect 298818 284023 298852 284051
rect 298880 284023 298914 284051
rect 298942 284023 298990 284051
rect -958 283989 298990 284023
rect -958 283961 -910 283989
rect -882 283961 -848 283989
rect -820 283961 -786 283989
rect -758 283961 -724 283989
rect -696 283961 4617 283989
rect 4645 283961 4679 283989
rect 4707 283961 4741 283989
rect 4769 283961 4803 283989
rect 4831 283961 19977 283989
rect 20005 283961 20039 283989
rect 20067 283961 20101 283989
rect 20129 283961 20163 283989
rect 20191 283961 35337 283989
rect 35365 283961 35399 283989
rect 35427 283961 35461 283989
rect 35489 283961 35523 283989
rect 35551 283961 50697 283989
rect 50725 283961 50759 283989
rect 50787 283961 50821 283989
rect 50849 283961 50883 283989
rect 50911 283961 66057 283989
rect 66085 283961 66119 283989
rect 66147 283961 66181 283989
rect 66209 283961 66243 283989
rect 66271 283961 81417 283989
rect 81445 283961 81479 283989
rect 81507 283961 81541 283989
rect 81569 283961 81603 283989
rect 81631 283961 96777 283989
rect 96805 283961 96839 283989
rect 96867 283961 96901 283989
rect 96929 283961 96963 283989
rect 96991 283961 112137 283989
rect 112165 283961 112199 283989
rect 112227 283961 112261 283989
rect 112289 283961 112323 283989
rect 112351 283961 127497 283989
rect 127525 283961 127559 283989
rect 127587 283961 127621 283989
rect 127649 283961 127683 283989
rect 127711 283961 142857 283989
rect 142885 283961 142919 283989
rect 142947 283961 142981 283989
rect 143009 283961 143043 283989
rect 143071 283961 158217 283989
rect 158245 283961 158279 283989
rect 158307 283961 158341 283989
rect 158369 283961 158403 283989
rect 158431 283961 173577 283989
rect 173605 283961 173639 283989
rect 173667 283961 173701 283989
rect 173729 283961 173763 283989
rect 173791 283961 188937 283989
rect 188965 283961 188999 283989
rect 189027 283961 189061 283989
rect 189089 283961 189123 283989
rect 189151 283961 204297 283989
rect 204325 283961 204359 283989
rect 204387 283961 204421 283989
rect 204449 283961 204483 283989
rect 204511 283961 219657 283989
rect 219685 283961 219719 283989
rect 219747 283961 219781 283989
rect 219809 283961 219843 283989
rect 219871 283961 235017 283989
rect 235045 283961 235079 283989
rect 235107 283961 235141 283989
rect 235169 283961 235203 283989
rect 235231 283961 250377 283989
rect 250405 283961 250439 283989
rect 250467 283961 250501 283989
rect 250529 283961 250563 283989
rect 250591 283961 265737 283989
rect 265765 283961 265799 283989
rect 265827 283961 265861 283989
rect 265889 283961 265923 283989
rect 265951 283961 281097 283989
rect 281125 283961 281159 283989
rect 281187 283961 281221 283989
rect 281249 283961 281283 283989
rect 281311 283961 296457 283989
rect 296485 283961 296519 283989
rect 296547 283961 296581 283989
rect 296609 283961 296643 283989
rect 296671 283961 298728 283989
rect 298756 283961 298790 283989
rect 298818 283961 298852 283989
rect 298880 283961 298914 283989
rect 298942 283961 298990 283989
rect -958 283913 298990 283961
rect -958 281175 298990 281223
rect -958 281147 -430 281175
rect -402 281147 -368 281175
rect -340 281147 -306 281175
rect -278 281147 -244 281175
rect -216 281147 2757 281175
rect 2785 281147 2819 281175
rect 2847 281147 2881 281175
rect 2909 281147 2943 281175
rect 2971 281147 18117 281175
rect 18145 281147 18179 281175
rect 18207 281147 18241 281175
rect 18269 281147 18303 281175
rect 18331 281147 33477 281175
rect 33505 281147 33539 281175
rect 33567 281147 33601 281175
rect 33629 281147 33663 281175
rect 33691 281147 48837 281175
rect 48865 281147 48899 281175
rect 48927 281147 48961 281175
rect 48989 281147 49023 281175
rect 49051 281147 64197 281175
rect 64225 281147 64259 281175
rect 64287 281147 64321 281175
rect 64349 281147 64383 281175
rect 64411 281147 79557 281175
rect 79585 281147 79619 281175
rect 79647 281147 79681 281175
rect 79709 281147 79743 281175
rect 79771 281147 94917 281175
rect 94945 281147 94979 281175
rect 95007 281147 95041 281175
rect 95069 281147 95103 281175
rect 95131 281147 110277 281175
rect 110305 281147 110339 281175
rect 110367 281147 110401 281175
rect 110429 281147 110463 281175
rect 110491 281147 125637 281175
rect 125665 281147 125699 281175
rect 125727 281147 125761 281175
rect 125789 281147 125823 281175
rect 125851 281147 140997 281175
rect 141025 281147 141059 281175
rect 141087 281147 141121 281175
rect 141149 281147 141183 281175
rect 141211 281147 156357 281175
rect 156385 281147 156419 281175
rect 156447 281147 156481 281175
rect 156509 281147 156543 281175
rect 156571 281147 171717 281175
rect 171745 281147 171779 281175
rect 171807 281147 171841 281175
rect 171869 281147 171903 281175
rect 171931 281147 187077 281175
rect 187105 281147 187139 281175
rect 187167 281147 187201 281175
rect 187229 281147 187263 281175
rect 187291 281147 202437 281175
rect 202465 281147 202499 281175
rect 202527 281147 202561 281175
rect 202589 281147 202623 281175
rect 202651 281147 217797 281175
rect 217825 281147 217859 281175
rect 217887 281147 217921 281175
rect 217949 281147 217983 281175
rect 218011 281147 233157 281175
rect 233185 281147 233219 281175
rect 233247 281147 233281 281175
rect 233309 281147 233343 281175
rect 233371 281147 248517 281175
rect 248545 281147 248579 281175
rect 248607 281147 248641 281175
rect 248669 281147 248703 281175
rect 248731 281147 263877 281175
rect 263905 281147 263939 281175
rect 263967 281147 264001 281175
rect 264029 281147 264063 281175
rect 264091 281147 279237 281175
rect 279265 281147 279299 281175
rect 279327 281147 279361 281175
rect 279389 281147 279423 281175
rect 279451 281147 294597 281175
rect 294625 281147 294659 281175
rect 294687 281147 294721 281175
rect 294749 281147 294783 281175
rect 294811 281147 298248 281175
rect 298276 281147 298310 281175
rect 298338 281147 298372 281175
rect 298400 281147 298434 281175
rect 298462 281147 298990 281175
rect -958 281113 298990 281147
rect -958 281085 -430 281113
rect -402 281085 -368 281113
rect -340 281085 -306 281113
rect -278 281085 -244 281113
rect -216 281085 2757 281113
rect 2785 281085 2819 281113
rect 2847 281085 2881 281113
rect 2909 281085 2943 281113
rect 2971 281085 18117 281113
rect 18145 281085 18179 281113
rect 18207 281085 18241 281113
rect 18269 281085 18303 281113
rect 18331 281085 33477 281113
rect 33505 281085 33539 281113
rect 33567 281085 33601 281113
rect 33629 281085 33663 281113
rect 33691 281085 48837 281113
rect 48865 281085 48899 281113
rect 48927 281085 48961 281113
rect 48989 281085 49023 281113
rect 49051 281085 64197 281113
rect 64225 281085 64259 281113
rect 64287 281085 64321 281113
rect 64349 281085 64383 281113
rect 64411 281085 79557 281113
rect 79585 281085 79619 281113
rect 79647 281085 79681 281113
rect 79709 281085 79743 281113
rect 79771 281085 94917 281113
rect 94945 281085 94979 281113
rect 95007 281085 95041 281113
rect 95069 281085 95103 281113
rect 95131 281085 110277 281113
rect 110305 281085 110339 281113
rect 110367 281085 110401 281113
rect 110429 281085 110463 281113
rect 110491 281085 125637 281113
rect 125665 281085 125699 281113
rect 125727 281085 125761 281113
rect 125789 281085 125823 281113
rect 125851 281085 140997 281113
rect 141025 281085 141059 281113
rect 141087 281085 141121 281113
rect 141149 281085 141183 281113
rect 141211 281085 156357 281113
rect 156385 281085 156419 281113
rect 156447 281085 156481 281113
rect 156509 281085 156543 281113
rect 156571 281085 171717 281113
rect 171745 281085 171779 281113
rect 171807 281085 171841 281113
rect 171869 281085 171903 281113
rect 171931 281085 187077 281113
rect 187105 281085 187139 281113
rect 187167 281085 187201 281113
rect 187229 281085 187263 281113
rect 187291 281085 202437 281113
rect 202465 281085 202499 281113
rect 202527 281085 202561 281113
rect 202589 281085 202623 281113
rect 202651 281085 217797 281113
rect 217825 281085 217859 281113
rect 217887 281085 217921 281113
rect 217949 281085 217983 281113
rect 218011 281085 233157 281113
rect 233185 281085 233219 281113
rect 233247 281085 233281 281113
rect 233309 281085 233343 281113
rect 233371 281085 248517 281113
rect 248545 281085 248579 281113
rect 248607 281085 248641 281113
rect 248669 281085 248703 281113
rect 248731 281085 263877 281113
rect 263905 281085 263939 281113
rect 263967 281085 264001 281113
rect 264029 281085 264063 281113
rect 264091 281085 279237 281113
rect 279265 281085 279299 281113
rect 279327 281085 279361 281113
rect 279389 281085 279423 281113
rect 279451 281085 294597 281113
rect 294625 281085 294659 281113
rect 294687 281085 294721 281113
rect 294749 281085 294783 281113
rect 294811 281085 298248 281113
rect 298276 281085 298310 281113
rect 298338 281085 298372 281113
rect 298400 281085 298434 281113
rect 298462 281085 298990 281113
rect -958 281051 298990 281085
rect -958 281023 -430 281051
rect -402 281023 -368 281051
rect -340 281023 -306 281051
rect -278 281023 -244 281051
rect -216 281023 2757 281051
rect 2785 281023 2819 281051
rect 2847 281023 2881 281051
rect 2909 281023 2943 281051
rect 2971 281023 18117 281051
rect 18145 281023 18179 281051
rect 18207 281023 18241 281051
rect 18269 281023 18303 281051
rect 18331 281023 33477 281051
rect 33505 281023 33539 281051
rect 33567 281023 33601 281051
rect 33629 281023 33663 281051
rect 33691 281023 48837 281051
rect 48865 281023 48899 281051
rect 48927 281023 48961 281051
rect 48989 281023 49023 281051
rect 49051 281023 64197 281051
rect 64225 281023 64259 281051
rect 64287 281023 64321 281051
rect 64349 281023 64383 281051
rect 64411 281023 79557 281051
rect 79585 281023 79619 281051
rect 79647 281023 79681 281051
rect 79709 281023 79743 281051
rect 79771 281023 94917 281051
rect 94945 281023 94979 281051
rect 95007 281023 95041 281051
rect 95069 281023 95103 281051
rect 95131 281023 110277 281051
rect 110305 281023 110339 281051
rect 110367 281023 110401 281051
rect 110429 281023 110463 281051
rect 110491 281023 125637 281051
rect 125665 281023 125699 281051
rect 125727 281023 125761 281051
rect 125789 281023 125823 281051
rect 125851 281023 140997 281051
rect 141025 281023 141059 281051
rect 141087 281023 141121 281051
rect 141149 281023 141183 281051
rect 141211 281023 156357 281051
rect 156385 281023 156419 281051
rect 156447 281023 156481 281051
rect 156509 281023 156543 281051
rect 156571 281023 171717 281051
rect 171745 281023 171779 281051
rect 171807 281023 171841 281051
rect 171869 281023 171903 281051
rect 171931 281023 187077 281051
rect 187105 281023 187139 281051
rect 187167 281023 187201 281051
rect 187229 281023 187263 281051
rect 187291 281023 202437 281051
rect 202465 281023 202499 281051
rect 202527 281023 202561 281051
rect 202589 281023 202623 281051
rect 202651 281023 217797 281051
rect 217825 281023 217859 281051
rect 217887 281023 217921 281051
rect 217949 281023 217983 281051
rect 218011 281023 233157 281051
rect 233185 281023 233219 281051
rect 233247 281023 233281 281051
rect 233309 281023 233343 281051
rect 233371 281023 248517 281051
rect 248545 281023 248579 281051
rect 248607 281023 248641 281051
rect 248669 281023 248703 281051
rect 248731 281023 263877 281051
rect 263905 281023 263939 281051
rect 263967 281023 264001 281051
rect 264029 281023 264063 281051
rect 264091 281023 279237 281051
rect 279265 281023 279299 281051
rect 279327 281023 279361 281051
rect 279389 281023 279423 281051
rect 279451 281023 294597 281051
rect 294625 281023 294659 281051
rect 294687 281023 294721 281051
rect 294749 281023 294783 281051
rect 294811 281023 298248 281051
rect 298276 281023 298310 281051
rect 298338 281023 298372 281051
rect 298400 281023 298434 281051
rect 298462 281023 298990 281051
rect -958 280989 298990 281023
rect -958 280961 -430 280989
rect -402 280961 -368 280989
rect -340 280961 -306 280989
rect -278 280961 -244 280989
rect -216 280961 2757 280989
rect 2785 280961 2819 280989
rect 2847 280961 2881 280989
rect 2909 280961 2943 280989
rect 2971 280961 18117 280989
rect 18145 280961 18179 280989
rect 18207 280961 18241 280989
rect 18269 280961 18303 280989
rect 18331 280961 33477 280989
rect 33505 280961 33539 280989
rect 33567 280961 33601 280989
rect 33629 280961 33663 280989
rect 33691 280961 48837 280989
rect 48865 280961 48899 280989
rect 48927 280961 48961 280989
rect 48989 280961 49023 280989
rect 49051 280961 64197 280989
rect 64225 280961 64259 280989
rect 64287 280961 64321 280989
rect 64349 280961 64383 280989
rect 64411 280961 79557 280989
rect 79585 280961 79619 280989
rect 79647 280961 79681 280989
rect 79709 280961 79743 280989
rect 79771 280961 94917 280989
rect 94945 280961 94979 280989
rect 95007 280961 95041 280989
rect 95069 280961 95103 280989
rect 95131 280961 110277 280989
rect 110305 280961 110339 280989
rect 110367 280961 110401 280989
rect 110429 280961 110463 280989
rect 110491 280961 125637 280989
rect 125665 280961 125699 280989
rect 125727 280961 125761 280989
rect 125789 280961 125823 280989
rect 125851 280961 140997 280989
rect 141025 280961 141059 280989
rect 141087 280961 141121 280989
rect 141149 280961 141183 280989
rect 141211 280961 156357 280989
rect 156385 280961 156419 280989
rect 156447 280961 156481 280989
rect 156509 280961 156543 280989
rect 156571 280961 171717 280989
rect 171745 280961 171779 280989
rect 171807 280961 171841 280989
rect 171869 280961 171903 280989
rect 171931 280961 187077 280989
rect 187105 280961 187139 280989
rect 187167 280961 187201 280989
rect 187229 280961 187263 280989
rect 187291 280961 202437 280989
rect 202465 280961 202499 280989
rect 202527 280961 202561 280989
rect 202589 280961 202623 280989
rect 202651 280961 217797 280989
rect 217825 280961 217859 280989
rect 217887 280961 217921 280989
rect 217949 280961 217983 280989
rect 218011 280961 233157 280989
rect 233185 280961 233219 280989
rect 233247 280961 233281 280989
rect 233309 280961 233343 280989
rect 233371 280961 248517 280989
rect 248545 280961 248579 280989
rect 248607 280961 248641 280989
rect 248669 280961 248703 280989
rect 248731 280961 263877 280989
rect 263905 280961 263939 280989
rect 263967 280961 264001 280989
rect 264029 280961 264063 280989
rect 264091 280961 279237 280989
rect 279265 280961 279299 280989
rect 279327 280961 279361 280989
rect 279389 280961 279423 280989
rect 279451 280961 294597 280989
rect 294625 280961 294659 280989
rect 294687 280961 294721 280989
rect 294749 280961 294783 280989
rect 294811 280961 298248 280989
rect 298276 280961 298310 280989
rect 298338 280961 298372 280989
rect 298400 280961 298434 280989
rect 298462 280961 298990 280989
rect -958 280913 298990 280961
rect -958 275175 298990 275223
rect -958 275147 -910 275175
rect -882 275147 -848 275175
rect -820 275147 -786 275175
rect -758 275147 -724 275175
rect -696 275147 4617 275175
rect 4645 275147 4679 275175
rect 4707 275147 4741 275175
rect 4769 275147 4803 275175
rect 4831 275147 19977 275175
rect 20005 275147 20039 275175
rect 20067 275147 20101 275175
rect 20129 275147 20163 275175
rect 20191 275147 35337 275175
rect 35365 275147 35399 275175
rect 35427 275147 35461 275175
rect 35489 275147 35523 275175
rect 35551 275147 50697 275175
rect 50725 275147 50759 275175
rect 50787 275147 50821 275175
rect 50849 275147 50883 275175
rect 50911 275147 66057 275175
rect 66085 275147 66119 275175
rect 66147 275147 66181 275175
rect 66209 275147 66243 275175
rect 66271 275147 81417 275175
rect 81445 275147 81479 275175
rect 81507 275147 81541 275175
rect 81569 275147 81603 275175
rect 81631 275147 96777 275175
rect 96805 275147 96839 275175
rect 96867 275147 96901 275175
rect 96929 275147 96963 275175
rect 96991 275147 112137 275175
rect 112165 275147 112199 275175
rect 112227 275147 112261 275175
rect 112289 275147 112323 275175
rect 112351 275147 127497 275175
rect 127525 275147 127559 275175
rect 127587 275147 127621 275175
rect 127649 275147 127683 275175
rect 127711 275147 142857 275175
rect 142885 275147 142919 275175
rect 142947 275147 142981 275175
rect 143009 275147 143043 275175
rect 143071 275147 158217 275175
rect 158245 275147 158279 275175
rect 158307 275147 158341 275175
rect 158369 275147 158403 275175
rect 158431 275147 173577 275175
rect 173605 275147 173639 275175
rect 173667 275147 173701 275175
rect 173729 275147 173763 275175
rect 173791 275147 188937 275175
rect 188965 275147 188999 275175
rect 189027 275147 189061 275175
rect 189089 275147 189123 275175
rect 189151 275147 204297 275175
rect 204325 275147 204359 275175
rect 204387 275147 204421 275175
rect 204449 275147 204483 275175
rect 204511 275147 219657 275175
rect 219685 275147 219719 275175
rect 219747 275147 219781 275175
rect 219809 275147 219843 275175
rect 219871 275147 235017 275175
rect 235045 275147 235079 275175
rect 235107 275147 235141 275175
rect 235169 275147 235203 275175
rect 235231 275147 250377 275175
rect 250405 275147 250439 275175
rect 250467 275147 250501 275175
rect 250529 275147 250563 275175
rect 250591 275147 265737 275175
rect 265765 275147 265799 275175
rect 265827 275147 265861 275175
rect 265889 275147 265923 275175
rect 265951 275147 281097 275175
rect 281125 275147 281159 275175
rect 281187 275147 281221 275175
rect 281249 275147 281283 275175
rect 281311 275147 296457 275175
rect 296485 275147 296519 275175
rect 296547 275147 296581 275175
rect 296609 275147 296643 275175
rect 296671 275147 298728 275175
rect 298756 275147 298790 275175
rect 298818 275147 298852 275175
rect 298880 275147 298914 275175
rect 298942 275147 298990 275175
rect -958 275113 298990 275147
rect -958 275085 -910 275113
rect -882 275085 -848 275113
rect -820 275085 -786 275113
rect -758 275085 -724 275113
rect -696 275085 4617 275113
rect 4645 275085 4679 275113
rect 4707 275085 4741 275113
rect 4769 275085 4803 275113
rect 4831 275085 19977 275113
rect 20005 275085 20039 275113
rect 20067 275085 20101 275113
rect 20129 275085 20163 275113
rect 20191 275085 35337 275113
rect 35365 275085 35399 275113
rect 35427 275085 35461 275113
rect 35489 275085 35523 275113
rect 35551 275085 50697 275113
rect 50725 275085 50759 275113
rect 50787 275085 50821 275113
rect 50849 275085 50883 275113
rect 50911 275085 66057 275113
rect 66085 275085 66119 275113
rect 66147 275085 66181 275113
rect 66209 275085 66243 275113
rect 66271 275085 81417 275113
rect 81445 275085 81479 275113
rect 81507 275085 81541 275113
rect 81569 275085 81603 275113
rect 81631 275085 96777 275113
rect 96805 275085 96839 275113
rect 96867 275085 96901 275113
rect 96929 275085 96963 275113
rect 96991 275085 112137 275113
rect 112165 275085 112199 275113
rect 112227 275085 112261 275113
rect 112289 275085 112323 275113
rect 112351 275085 127497 275113
rect 127525 275085 127559 275113
rect 127587 275085 127621 275113
rect 127649 275085 127683 275113
rect 127711 275085 142857 275113
rect 142885 275085 142919 275113
rect 142947 275085 142981 275113
rect 143009 275085 143043 275113
rect 143071 275085 158217 275113
rect 158245 275085 158279 275113
rect 158307 275085 158341 275113
rect 158369 275085 158403 275113
rect 158431 275085 173577 275113
rect 173605 275085 173639 275113
rect 173667 275085 173701 275113
rect 173729 275085 173763 275113
rect 173791 275085 188937 275113
rect 188965 275085 188999 275113
rect 189027 275085 189061 275113
rect 189089 275085 189123 275113
rect 189151 275085 204297 275113
rect 204325 275085 204359 275113
rect 204387 275085 204421 275113
rect 204449 275085 204483 275113
rect 204511 275085 219657 275113
rect 219685 275085 219719 275113
rect 219747 275085 219781 275113
rect 219809 275085 219843 275113
rect 219871 275085 235017 275113
rect 235045 275085 235079 275113
rect 235107 275085 235141 275113
rect 235169 275085 235203 275113
rect 235231 275085 250377 275113
rect 250405 275085 250439 275113
rect 250467 275085 250501 275113
rect 250529 275085 250563 275113
rect 250591 275085 265737 275113
rect 265765 275085 265799 275113
rect 265827 275085 265861 275113
rect 265889 275085 265923 275113
rect 265951 275085 281097 275113
rect 281125 275085 281159 275113
rect 281187 275085 281221 275113
rect 281249 275085 281283 275113
rect 281311 275085 296457 275113
rect 296485 275085 296519 275113
rect 296547 275085 296581 275113
rect 296609 275085 296643 275113
rect 296671 275085 298728 275113
rect 298756 275085 298790 275113
rect 298818 275085 298852 275113
rect 298880 275085 298914 275113
rect 298942 275085 298990 275113
rect -958 275051 298990 275085
rect -958 275023 -910 275051
rect -882 275023 -848 275051
rect -820 275023 -786 275051
rect -758 275023 -724 275051
rect -696 275023 4617 275051
rect 4645 275023 4679 275051
rect 4707 275023 4741 275051
rect 4769 275023 4803 275051
rect 4831 275023 19977 275051
rect 20005 275023 20039 275051
rect 20067 275023 20101 275051
rect 20129 275023 20163 275051
rect 20191 275023 35337 275051
rect 35365 275023 35399 275051
rect 35427 275023 35461 275051
rect 35489 275023 35523 275051
rect 35551 275023 50697 275051
rect 50725 275023 50759 275051
rect 50787 275023 50821 275051
rect 50849 275023 50883 275051
rect 50911 275023 66057 275051
rect 66085 275023 66119 275051
rect 66147 275023 66181 275051
rect 66209 275023 66243 275051
rect 66271 275023 81417 275051
rect 81445 275023 81479 275051
rect 81507 275023 81541 275051
rect 81569 275023 81603 275051
rect 81631 275023 96777 275051
rect 96805 275023 96839 275051
rect 96867 275023 96901 275051
rect 96929 275023 96963 275051
rect 96991 275023 112137 275051
rect 112165 275023 112199 275051
rect 112227 275023 112261 275051
rect 112289 275023 112323 275051
rect 112351 275023 127497 275051
rect 127525 275023 127559 275051
rect 127587 275023 127621 275051
rect 127649 275023 127683 275051
rect 127711 275023 142857 275051
rect 142885 275023 142919 275051
rect 142947 275023 142981 275051
rect 143009 275023 143043 275051
rect 143071 275023 158217 275051
rect 158245 275023 158279 275051
rect 158307 275023 158341 275051
rect 158369 275023 158403 275051
rect 158431 275023 173577 275051
rect 173605 275023 173639 275051
rect 173667 275023 173701 275051
rect 173729 275023 173763 275051
rect 173791 275023 188937 275051
rect 188965 275023 188999 275051
rect 189027 275023 189061 275051
rect 189089 275023 189123 275051
rect 189151 275023 204297 275051
rect 204325 275023 204359 275051
rect 204387 275023 204421 275051
rect 204449 275023 204483 275051
rect 204511 275023 219657 275051
rect 219685 275023 219719 275051
rect 219747 275023 219781 275051
rect 219809 275023 219843 275051
rect 219871 275023 235017 275051
rect 235045 275023 235079 275051
rect 235107 275023 235141 275051
rect 235169 275023 235203 275051
rect 235231 275023 250377 275051
rect 250405 275023 250439 275051
rect 250467 275023 250501 275051
rect 250529 275023 250563 275051
rect 250591 275023 265737 275051
rect 265765 275023 265799 275051
rect 265827 275023 265861 275051
rect 265889 275023 265923 275051
rect 265951 275023 281097 275051
rect 281125 275023 281159 275051
rect 281187 275023 281221 275051
rect 281249 275023 281283 275051
rect 281311 275023 296457 275051
rect 296485 275023 296519 275051
rect 296547 275023 296581 275051
rect 296609 275023 296643 275051
rect 296671 275023 298728 275051
rect 298756 275023 298790 275051
rect 298818 275023 298852 275051
rect 298880 275023 298914 275051
rect 298942 275023 298990 275051
rect -958 274989 298990 275023
rect -958 274961 -910 274989
rect -882 274961 -848 274989
rect -820 274961 -786 274989
rect -758 274961 -724 274989
rect -696 274961 4617 274989
rect 4645 274961 4679 274989
rect 4707 274961 4741 274989
rect 4769 274961 4803 274989
rect 4831 274961 19977 274989
rect 20005 274961 20039 274989
rect 20067 274961 20101 274989
rect 20129 274961 20163 274989
rect 20191 274961 35337 274989
rect 35365 274961 35399 274989
rect 35427 274961 35461 274989
rect 35489 274961 35523 274989
rect 35551 274961 50697 274989
rect 50725 274961 50759 274989
rect 50787 274961 50821 274989
rect 50849 274961 50883 274989
rect 50911 274961 66057 274989
rect 66085 274961 66119 274989
rect 66147 274961 66181 274989
rect 66209 274961 66243 274989
rect 66271 274961 81417 274989
rect 81445 274961 81479 274989
rect 81507 274961 81541 274989
rect 81569 274961 81603 274989
rect 81631 274961 96777 274989
rect 96805 274961 96839 274989
rect 96867 274961 96901 274989
rect 96929 274961 96963 274989
rect 96991 274961 112137 274989
rect 112165 274961 112199 274989
rect 112227 274961 112261 274989
rect 112289 274961 112323 274989
rect 112351 274961 127497 274989
rect 127525 274961 127559 274989
rect 127587 274961 127621 274989
rect 127649 274961 127683 274989
rect 127711 274961 142857 274989
rect 142885 274961 142919 274989
rect 142947 274961 142981 274989
rect 143009 274961 143043 274989
rect 143071 274961 158217 274989
rect 158245 274961 158279 274989
rect 158307 274961 158341 274989
rect 158369 274961 158403 274989
rect 158431 274961 173577 274989
rect 173605 274961 173639 274989
rect 173667 274961 173701 274989
rect 173729 274961 173763 274989
rect 173791 274961 188937 274989
rect 188965 274961 188999 274989
rect 189027 274961 189061 274989
rect 189089 274961 189123 274989
rect 189151 274961 204297 274989
rect 204325 274961 204359 274989
rect 204387 274961 204421 274989
rect 204449 274961 204483 274989
rect 204511 274961 219657 274989
rect 219685 274961 219719 274989
rect 219747 274961 219781 274989
rect 219809 274961 219843 274989
rect 219871 274961 235017 274989
rect 235045 274961 235079 274989
rect 235107 274961 235141 274989
rect 235169 274961 235203 274989
rect 235231 274961 250377 274989
rect 250405 274961 250439 274989
rect 250467 274961 250501 274989
rect 250529 274961 250563 274989
rect 250591 274961 265737 274989
rect 265765 274961 265799 274989
rect 265827 274961 265861 274989
rect 265889 274961 265923 274989
rect 265951 274961 281097 274989
rect 281125 274961 281159 274989
rect 281187 274961 281221 274989
rect 281249 274961 281283 274989
rect 281311 274961 296457 274989
rect 296485 274961 296519 274989
rect 296547 274961 296581 274989
rect 296609 274961 296643 274989
rect 296671 274961 298728 274989
rect 298756 274961 298790 274989
rect 298818 274961 298852 274989
rect 298880 274961 298914 274989
rect 298942 274961 298990 274989
rect -958 274913 298990 274961
rect -958 272175 298990 272223
rect -958 272147 -430 272175
rect -402 272147 -368 272175
rect -340 272147 -306 272175
rect -278 272147 -244 272175
rect -216 272147 2757 272175
rect 2785 272147 2819 272175
rect 2847 272147 2881 272175
rect 2909 272147 2943 272175
rect 2971 272147 18117 272175
rect 18145 272147 18179 272175
rect 18207 272147 18241 272175
rect 18269 272147 18303 272175
rect 18331 272147 33477 272175
rect 33505 272147 33539 272175
rect 33567 272147 33601 272175
rect 33629 272147 33663 272175
rect 33691 272147 48837 272175
rect 48865 272147 48899 272175
rect 48927 272147 48961 272175
rect 48989 272147 49023 272175
rect 49051 272147 64197 272175
rect 64225 272147 64259 272175
rect 64287 272147 64321 272175
rect 64349 272147 64383 272175
rect 64411 272147 79557 272175
rect 79585 272147 79619 272175
rect 79647 272147 79681 272175
rect 79709 272147 79743 272175
rect 79771 272147 94917 272175
rect 94945 272147 94979 272175
rect 95007 272147 95041 272175
rect 95069 272147 95103 272175
rect 95131 272147 110277 272175
rect 110305 272147 110339 272175
rect 110367 272147 110401 272175
rect 110429 272147 110463 272175
rect 110491 272147 125637 272175
rect 125665 272147 125699 272175
rect 125727 272147 125761 272175
rect 125789 272147 125823 272175
rect 125851 272147 140997 272175
rect 141025 272147 141059 272175
rect 141087 272147 141121 272175
rect 141149 272147 141183 272175
rect 141211 272147 156357 272175
rect 156385 272147 156419 272175
rect 156447 272147 156481 272175
rect 156509 272147 156543 272175
rect 156571 272147 171717 272175
rect 171745 272147 171779 272175
rect 171807 272147 171841 272175
rect 171869 272147 171903 272175
rect 171931 272147 187077 272175
rect 187105 272147 187139 272175
rect 187167 272147 187201 272175
rect 187229 272147 187263 272175
rect 187291 272147 202437 272175
rect 202465 272147 202499 272175
rect 202527 272147 202561 272175
rect 202589 272147 202623 272175
rect 202651 272147 217797 272175
rect 217825 272147 217859 272175
rect 217887 272147 217921 272175
rect 217949 272147 217983 272175
rect 218011 272147 233157 272175
rect 233185 272147 233219 272175
rect 233247 272147 233281 272175
rect 233309 272147 233343 272175
rect 233371 272147 248517 272175
rect 248545 272147 248579 272175
rect 248607 272147 248641 272175
rect 248669 272147 248703 272175
rect 248731 272147 263877 272175
rect 263905 272147 263939 272175
rect 263967 272147 264001 272175
rect 264029 272147 264063 272175
rect 264091 272147 279237 272175
rect 279265 272147 279299 272175
rect 279327 272147 279361 272175
rect 279389 272147 279423 272175
rect 279451 272147 294597 272175
rect 294625 272147 294659 272175
rect 294687 272147 294721 272175
rect 294749 272147 294783 272175
rect 294811 272147 298248 272175
rect 298276 272147 298310 272175
rect 298338 272147 298372 272175
rect 298400 272147 298434 272175
rect 298462 272147 298990 272175
rect -958 272113 298990 272147
rect -958 272085 -430 272113
rect -402 272085 -368 272113
rect -340 272085 -306 272113
rect -278 272085 -244 272113
rect -216 272085 2757 272113
rect 2785 272085 2819 272113
rect 2847 272085 2881 272113
rect 2909 272085 2943 272113
rect 2971 272085 18117 272113
rect 18145 272085 18179 272113
rect 18207 272085 18241 272113
rect 18269 272085 18303 272113
rect 18331 272085 33477 272113
rect 33505 272085 33539 272113
rect 33567 272085 33601 272113
rect 33629 272085 33663 272113
rect 33691 272085 48837 272113
rect 48865 272085 48899 272113
rect 48927 272085 48961 272113
rect 48989 272085 49023 272113
rect 49051 272085 64197 272113
rect 64225 272085 64259 272113
rect 64287 272085 64321 272113
rect 64349 272085 64383 272113
rect 64411 272085 79557 272113
rect 79585 272085 79619 272113
rect 79647 272085 79681 272113
rect 79709 272085 79743 272113
rect 79771 272085 94917 272113
rect 94945 272085 94979 272113
rect 95007 272085 95041 272113
rect 95069 272085 95103 272113
rect 95131 272085 110277 272113
rect 110305 272085 110339 272113
rect 110367 272085 110401 272113
rect 110429 272085 110463 272113
rect 110491 272085 125637 272113
rect 125665 272085 125699 272113
rect 125727 272085 125761 272113
rect 125789 272085 125823 272113
rect 125851 272085 140997 272113
rect 141025 272085 141059 272113
rect 141087 272085 141121 272113
rect 141149 272085 141183 272113
rect 141211 272085 156357 272113
rect 156385 272085 156419 272113
rect 156447 272085 156481 272113
rect 156509 272085 156543 272113
rect 156571 272085 171717 272113
rect 171745 272085 171779 272113
rect 171807 272085 171841 272113
rect 171869 272085 171903 272113
rect 171931 272085 187077 272113
rect 187105 272085 187139 272113
rect 187167 272085 187201 272113
rect 187229 272085 187263 272113
rect 187291 272085 202437 272113
rect 202465 272085 202499 272113
rect 202527 272085 202561 272113
rect 202589 272085 202623 272113
rect 202651 272085 217797 272113
rect 217825 272085 217859 272113
rect 217887 272085 217921 272113
rect 217949 272085 217983 272113
rect 218011 272085 233157 272113
rect 233185 272085 233219 272113
rect 233247 272085 233281 272113
rect 233309 272085 233343 272113
rect 233371 272085 248517 272113
rect 248545 272085 248579 272113
rect 248607 272085 248641 272113
rect 248669 272085 248703 272113
rect 248731 272085 263877 272113
rect 263905 272085 263939 272113
rect 263967 272085 264001 272113
rect 264029 272085 264063 272113
rect 264091 272085 279237 272113
rect 279265 272085 279299 272113
rect 279327 272085 279361 272113
rect 279389 272085 279423 272113
rect 279451 272085 294597 272113
rect 294625 272085 294659 272113
rect 294687 272085 294721 272113
rect 294749 272085 294783 272113
rect 294811 272085 298248 272113
rect 298276 272085 298310 272113
rect 298338 272085 298372 272113
rect 298400 272085 298434 272113
rect 298462 272085 298990 272113
rect -958 272051 298990 272085
rect -958 272023 -430 272051
rect -402 272023 -368 272051
rect -340 272023 -306 272051
rect -278 272023 -244 272051
rect -216 272023 2757 272051
rect 2785 272023 2819 272051
rect 2847 272023 2881 272051
rect 2909 272023 2943 272051
rect 2971 272023 18117 272051
rect 18145 272023 18179 272051
rect 18207 272023 18241 272051
rect 18269 272023 18303 272051
rect 18331 272023 33477 272051
rect 33505 272023 33539 272051
rect 33567 272023 33601 272051
rect 33629 272023 33663 272051
rect 33691 272023 48837 272051
rect 48865 272023 48899 272051
rect 48927 272023 48961 272051
rect 48989 272023 49023 272051
rect 49051 272023 64197 272051
rect 64225 272023 64259 272051
rect 64287 272023 64321 272051
rect 64349 272023 64383 272051
rect 64411 272023 79557 272051
rect 79585 272023 79619 272051
rect 79647 272023 79681 272051
rect 79709 272023 79743 272051
rect 79771 272023 94917 272051
rect 94945 272023 94979 272051
rect 95007 272023 95041 272051
rect 95069 272023 95103 272051
rect 95131 272023 110277 272051
rect 110305 272023 110339 272051
rect 110367 272023 110401 272051
rect 110429 272023 110463 272051
rect 110491 272023 125637 272051
rect 125665 272023 125699 272051
rect 125727 272023 125761 272051
rect 125789 272023 125823 272051
rect 125851 272023 140997 272051
rect 141025 272023 141059 272051
rect 141087 272023 141121 272051
rect 141149 272023 141183 272051
rect 141211 272023 156357 272051
rect 156385 272023 156419 272051
rect 156447 272023 156481 272051
rect 156509 272023 156543 272051
rect 156571 272023 171717 272051
rect 171745 272023 171779 272051
rect 171807 272023 171841 272051
rect 171869 272023 171903 272051
rect 171931 272023 187077 272051
rect 187105 272023 187139 272051
rect 187167 272023 187201 272051
rect 187229 272023 187263 272051
rect 187291 272023 202437 272051
rect 202465 272023 202499 272051
rect 202527 272023 202561 272051
rect 202589 272023 202623 272051
rect 202651 272023 217797 272051
rect 217825 272023 217859 272051
rect 217887 272023 217921 272051
rect 217949 272023 217983 272051
rect 218011 272023 233157 272051
rect 233185 272023 233219 272051
rect 233247 272023 233281 272051
rect 233309 272023 233343 272051
rect 233371 272023 248517 272051
rect 248545 272023 248579 272051
rect 248607 272023 248641 272051
rect 248669 272023 248703 272051
rect 248731 272023 263877 272051
rect 263905 272023 263939 272051
rect 263967 272023 264001 272051
rect 264029 272023 264063 272051
rect 264091 272023 279237 272051
rect 279265 272023 279299 272051
rect 279327 272023 279361 272051
rect 279389 272023 279423 272051
rect 279451 272023 294597 272051
rect 294625 272023 294659 272051
rect 294687 272023 294721 272051
rect 294749 272023 294783 272051
rect 294811 272023 298248 272051
rect 298276 272023 298310 272051
rect 298338 272023 298372 272051
rect 298400 272023 298434 272051
rect 298462 272023 298990 272051
rect -958 271989 298990 272023
rect -958 271961 -430 271989
rect -402 271961 -368 271989
rect -340 271961 -306 271989
rect -278 271961 -244 271989
rect -216 271961 2757 271989
rect 2785 271961 2819 271989
rect 2847 271961 2881 271989
rect 2909 271961 2943 271989
rect 2971 271961 18117 271989
rect 18145 271961 18179 271989
rect 18207 271961 18241 271989
rect 18269 271961 18303 271989
rect 18331 271961 33477 271989
rect 33505 271961 33539 271989
rect 33567 271961 33601 271989
rect 33629 271961 33663 271989
rect 33691 271961 48837 271989
rect 48865 271961 48899 271989
rect 48927 271961 48961 271989
rect 48989 271961 49023 271989
rect 49051 271961 64197 271989
rect 64225 271961 64259 271989
rect 64287 271961 64321 271989
rect 64349 271961 64383 271989
rect 64411 271961 79557 271989
rect 79585 271961 79619 271989
rect 79647 271961 79681 271989
rect 79709 271961 79743 271989
rect 79771 271961 94917 271989
rect 94945 271961 94979 271989
rect 95007 271961 95041 271989
rect 95069 271961 95103 271989
rect 95131 271961 110277 271989
rect 110305 271961 110339 271989
rect 110367 271961 110401 271989
rect 110429 271961 110463 271989
rect 110491 271961 125637 271989
rect 125665 271961 125699 271989
rect 125727 271961 125761 271989
rect 125789 271961 125823 271989
rect 125851 271961 140997 271989
rect 141025 271961 141059 271989
rect 141087 271961 141121 271989
rect 141149 271961 141183 271989
rect 141211 271961 156357 271989
rect 156385 271961 156419 271989
rect 156447 271961 156481 271989
rect 156509 271961 156543 271989
rect 156571 271961 171717 271989
rect 171745 271961 171779 271989
rect 171807 271961 171841 271989
rect 171869 271961 171903 271989
rect 171931 271961 187077 271989
rect 187105 271961 187139 271989
rect 187167 271961 187201 271989
rect 187229 271961 187263 271989
rect 187291 271961 202437 271989
rect 202465 271961 202499 271989
rect 202527 271961 202561 271989
rect 202589 271961 202623 271989
rect 202651 271961 217797 271989
rect 217825 271961 217859 271989
rect 217887 271961 217921 271989
rect 217949 271961 217983 271989
rect 218011 271961 233157 271989
rect 233185 271961 233219 271989
rect 233247 271961 233281 271989
rect 233309 271961 233343 271989
rect 233371 271961 248517 271989
rect 248545 271961 248579 271989
rect 248607 271961 248641 271989
rect 248669 271961 248703 271989
rect 248731 271961 263877 271989
rect 263905 271961 263939 271989
rect 263967 271961 264001 271989
rect 264029 271961 264063 271989
rect 264091 271961 279237 271989
rect 279265 271961 279299 271989
rect 279327 271961 279361 271989
rect 279389 271961 279423 271989
rect 279451 271961 294597 271989
rect 294625 271961 294659 271989
rect 294687 271961 294721 271989
rect 294749 271961 294783 271989
rect 294811 271961 298248 271989
rect 298276 271961 298310 271989
rect 298338 271961 298372 271989
rect 298400 271961 298434 271989
rect 298462 271961 298990 271989
rect -958 271913 298990 271961
rect -958 266175 298990 266223
rect -958 266147 -910 266175
rect -882 266147 -848 266175
rect -820 266147 -786 266175
rect -758 266147 -724 266175
rect -696 266147 4617 266175
rect 4645 266147 4679 266175
rect 4707 266147 4741 266175
rect 4769 266147 4803 266175
rect 4831 266147 19977 266175
rect 20005 266147 20039 266175
rect 20067 266147 20101 266175
rect 20129 266147 20163 266175
rect 20191 266147 35337 266175
rect 35365 266147 35399 266175
rect 35427 266147 35461 266175
rect 35489 266147 35523 266175
rect 35551 266147 50697 266175
rect 50725 266147 50759 266175
rect 50787 266147 50821 266175
rect 50849 266147 50883 266175
rect 50911 266147 66057 266175
rect 66085 266147 66119 266175
rect 66147 266147 66181 266175
rect 66209 266147 66243 266175
rect 66271 266147 81417 266175
rect 81445 266147 81479 266175
rect 81507 266147 81541 266175
rect 81569 266147 81603 266175
rect 81631 266147 96777 266175
rect 96805 266147 96839 266175
rect 96867 266147 96901 266175
rect 96929 266147 96963 266175
rect 96991 266147 112137 266175
rect 112165 266147 112199 266175
rect 112227 266147 112261 266175
rect 112289 266147 112323 266175
rect 112351 266147 127497 266175
rect 127525 266147 127559 266175
rect 127587 266147 127621 266175
rect 127649 266147 127683 266175
rect 127711 266147 142857 266175
rect 142885 266147 142919 266175
rect 142947 266147 142981 266175
rect 143009 266147 143043 266175
rect 143071 266147 158217 266175
rect 158245 266147 158279 266175
rect 158307 266147 158341 266175
rect 158369 266147 158403 266175
rect 158431 266147 173577 266175
rect 173605 266147 173639 266175
rect 173667 266147 173701 266175
rect 173729 266147 173763 266175
rect 173791 266147 188937 266175
rect 188965 266147 188999 266175
rect 189027 266147 189061 266175
rect 189089 266147 189123 266175
rect 189151 266147 204297 266175
rect 204325 266147 204359 266175
rect 204387 266147 204421 266175
rect 204449 266147 204483 266175
rect 204511 266147 219657 266175
rect 219685 266147 219719 266175
rect 219747 266147 219781 266175
rect 219809 266147 219843 266175
rect 219871 266147 235017 266175
rect 235045 266147 235079 266175
rect 235107 266147 235141 266175
rect 235169 266147 235203 266175
rect 235231 266147 250377 266175
rect 250405 266147 250439 266175
rect 250467 266147 250501 266175
rect 250529 266147 250563 266175
rect 250591 266147 265737 266175
rect 265765 266147 265799 266175
rect 265827 266147 265861 266175
rect 265889 266147 265923 266175
rect 265951 266147 281097 266175
rect 281125 266147 281159 266175
rect 281187 266147 281221 266175
rect 281249 266147 281283 266175
rect 281311 266147 296457 266175
rect 296485 266147 296519 266175
rect 296547 266147 296581 266175
rect 296609 266147 296643 266175
rect 296671 266147 298728 266175
rect 298756 266147 298790 266175
rect 298818 266147 298852 266175
rect 298880 266147 298914 266175
rect 298942 266147 298990 266175
rect -958 266113 298990 266147
rect -958 266085 -910 266113
rect -882 266085 -848 266113
rect -820 266085 -786 266113
rect -758 266085 -724 266113
rect -696 266085 4617 266113
rect 4645 266085 4679 266113
rect 4707 266085 4741 266113
rect 4769 266085 4803 266113
rect 4831 266085 19977 266113
rect 20005 266085 20039 266113
rect 20067 266085 20101 266113
rect 20129 266085 20163 266113
rect 20191 266085 35337 266113
rect 35365 266085 35399 266113
rect 35427 266085 35461 266113
rect 35489 266085 35523 266113
rect 35551 266085 50697 266113
rect 50725 266085 50759 266113
rect 50787 266085 50821 266113
rect 50849 266085 50883 266113
rect 50911 266085 66057 266113
rect 66085 266085 66119 266113
rect 66147 266085 66181 266113
rect 66209 266085 66243 266113
rect 66271 266085 81417 266113
rect 81445 266085 81479 266113
rect 81507 266085 81541 266113
rect 81569 266085 81603 266113
rect 81631 266085 96777 266113
rect 96805 266085 96839 266113
rect 96867 266085 96901 266113
rect 96929 266085 96963 266113
rect 96991 266085 112137 266113
rect 112165 266085 112199 266113
rect 112227 266085 112261 266113
rect 112289 266085 112323 266113
rect 112351 266085 127497 266113
rect 127525 266085 127559 266113
rect 127587 266085 127621 266113
rect 127649 266085 127683 266113
rect 127711 266085 142857 266113
rect 142885 266085 142919 266113
rect 142947 266085 142981 266113
rect 143009 266085 143043 266113
rect 143071 266085 158217 266113
rect 158245 266085 158279 266113
rect 158307 266085 158341 266113
rect 158369 266085 158403 266113
rect 158431 266085 173577 266113
rect 173605 266085 173639 266113
rect 173667 266085 173701 266113
rect 173729 266085 173763 266113
rect 173791 266085 188937 266113
rect 188965 266085 188999 266113
rect 189027 266085 189061 266113
rect 189089 266085 189123 266113
rect 189151 266085 204297 266113
rect 204325 266085 204359 266113
rect 204387 266085 204421 266113
rect 204449 266085 204483 266113
rect 204511 266085 219657 266113
rect 219685 266085 219719 266113
rect 219747 266085 219781 266113
rect 219809 266085 219843 266113
rect 219871 266085 235017 266113
rect 235045 266085 235079 266113
rect 235107 266085 235141 266113
rect 235169 266085 235203 266113
rect 235231 266085 250377 266113
rect 250405 266085 250439 266113
rect 250467 266085 250501 266113
rect 250529 266085 250563 266113
rect 250591 266085 265737 266113
rect 265765 266085 265799 266113
rect 265827 266085 265861 266113
rect 265889 266085 265923 266113
rect 265951 266085 281097 266113
rect 281125 266085 281159 266113
rect 281187 266085 281221 266113
rect 281249 266085 281283 266113
rect 281311 266085 296457 266113
rect 296485 266085 296519 266113
rect 296547 266085 296581 266113
rect 296609 266085 296643 266113
rect 296671 266085 298728 266113
rect 298756 266085 298790 266113
rect 298818 266085 298852 266113
rect 298880 266085 298914 266113
rect 298942 266085 298990 266113
rect -958 266051 298990 266085
rect -958 266023 -910 266051
rect -882 266023 -848 266051
rect -820 266023 -786 266051
rect -758 266023 -724 266051
rect -696 266023 4617 266051
rect 4645 266023 4679 266051
rect 4707 266023 4741 266051
rect 4769 266023 4803 266051
rect 4831 266023 19977 266051
rect 20005 266023 20039 266051
rect 20067 266023 20101 266051
rect 20129 266023 20163 266051
rect 20191 266023 35337 266051
rect 35365 266023 35399 266051
rect 35427 266023 35461 266051
rect 35489 266023 35523 266051
rect 35551 266023 50697 266051
rect 50725 266023 50759 266051
rect 50787 266023 50821 266051
rect 50849 266023 50883 266051
rect 50911 266023 66057 266051
rect 66085 266023 66119 266051
rect 66147 266023 66181 266051
rect 66209 266023 66243 266051
rect 66271 266023 81417 266051
rect 81445 266023 81479 266051
rect 81507 266023 81541 266051
rect 81569 266023 81603 266051
rect 81631 266023 96777 266051
rect 96805 266023 96839 266051
rect 96867 266023 96901 266051
rect 96929 266023 96963 266051
rect 96991 266023 112137 266051
rect 112165 266023 112199 266051
rect 112227 266023 112261 266051
rect 112289 266023 112323 266051
rect 112351 266023 127497 266051
rect 127525 266023 127559 266051
rect 127587 266023 127621 266051
rect 127649 266023 127683 266051
rect 127711 266023 142857 266051
rect 142885 266023 142919 266051
rect 142947 266023 142981 266051
rect 143009 266023 143043 266051
rect 143071 266023 158217 266051
rect 158245 266023 158279 266051
rect 158307 266023 158341 266051
rect 158369 266023 158403 266051
rect 158431 266023 173577 266051
rect 173605 266023 173639 266051
rect 173667 266023 173701 266051
rect 173729 266023 173763 266051
rect 173791 266023 188937 266051
rect 188965 266023 188999 266051
rect 189027 266023 189061 266051
rect 189089 266023 189123 266051
rect 189151 266023 204297 266051
rect 204325 266023 204359 266051
rect 204387 266023 204421 266051
rect 204449 266023 204483 266051
rect 204511 266023 219657 266051
rect 219685 266023 219719 266051
rect 219747 266023 219781 266051
rect 219809 266023 219843 266051
rect 219871 266023 235017 266051
rect 235045 266023 235079 266051
rect 235107 266023 235141 266051
rect 235169 266023 235203 266051
rect 235231 266023 250377 266051
rect 250405 266023 250439 266051
rect 250467 266023 250501 266051
rect 250529 266023 250563 266051
rect 250591 266023 265737 266051
rect 265765 266023 265799 266051
rect 265827 266023 265861 266051
rect 265889 266023 265923 266051
rect 265951 266023 281097 266051
rect 281125 266023 281159 266051
rect 281187 266023 281221 266051
rect 281249 266023 281283 266051
rect 281311 266023 296457 266051
rect 296485 266023 296519 266051
rect 296547 266023 296581 266051
rect 296609 266023 296643 266051
rect 296671 266023 298728 266051
rect 298756 266023 298790 266051
rect 298818 266023 298852 266051
rect 298880 266023 298914 266051
rect 298942 266023 298990 266051
rect -958 265989 298990 266023
rect -958 265961 -910 265989
rect -882 265961 -848 265989
rect -820 265961 -786 265989
rect -758 265961 -724 265989
rect -696 265961 4617 265989
rect 4645 265961 4679 265989
rect 4707 265961 4741 265989
rect 4769 265961 4803 265989
rect 4831 265961 19977 265989
rect 20005 265961 20039 265989
rect 20067 265961 20101 265989
rect 20129 265961 20163 265989
rect 20191 265961 35337 265989
rect 35365 265961 35399 265989
rect 35427 265961 35461 265989
rect 35489 265961 35523 265989
rect 35551 265961 50697 265989
rect 50725 265961 50759 265989
rect 50787 265961 50821 265989
rect 50849 265961 50883 265989
rect 50911 265961 66057 265989
rect 66085 265961 66119 265989
rect 66147 265961 66181 265989
rect 66209 265961 66243 265989
rect 66271 265961 81417 265989
rect 81445 265961 81479 265989
rect 81507 265961 81541 265989
rect 81569 265961 81603 265989
rect 81631 265961 96777 265989
rect 96805 265961 96839 265989
rect 96867 265961 96901 265989
rect 96929 265961 96963 265989
rect 96991 265961 112137 265989
rect 112165 265961 112199 265989
rect 112227 265961 112261 265989
rect 112289 265961 112323 265989
rect 112351 265961 127497 265989
rect 127525 265961 127559 265989
rect 127587 265961 127621 265989
rect 127649 265961 127683 265989
rect 127711 265961 142857 265989
rect 142885 265961 142919 265989
rect 142947 265961 142981 265989
rect 143009 265961 143043 265989
rect 143071 265961 158217 265989
rect 158245 265961 158279 265989
rect 158307 265961 158341 265989
rect 158369 265961 158403 265989
rect 158431 265961 173577 265989
rect 173605 265961 173639 265989
rect 173667 265961 173701 265989
rect 173729 265961 173763 265989
rect 173791 265961 188937 265989
rect 188965 265961 188999 265989
rect 189027 265961 189061 265989
rect 189089 265961 189123 265989
rect 189151 265961 204297 265989
rect 204325 265961 204359 265989
rect 204387 265961 204421 265989
rect 204449 265961 204483 265989
rect 204511 265961 219657 265989
rect 219685 265961 219719 265989
rect 219747 265961 219781 265989
rect 219809 265961 219843 265989
rect 219871 265961 235017 265989
rect 235045 265961 235079 265989
rect 235107 265961 235141 265989
rect 235169 265961 235203 265989
rect 235231 265961 250377 265989
rect 250405 265961 250439 265989
rect 250467 265961 250501 265989
rect 250529 265961 250563 265989
rect 250591 265961 265737 265989
rect 265765 265961 265799 265989
rect 265827 265961 265861 265989
rect 265889 265961 265923 265989
rect 265951 265961 281097 265989
rect 281125 265961 281159 265989
rect 281187 265961 281221 265989
rect 281249 265961 281283 265989
rect 281311 265961 296457 265989
rect 296485 265961 296519 265989
rect 296547 265961 296581 265989
rect 296609 265961 296643 265989
rect 296671 265961 298728 265989
rect 298756 265961 298790 265989
rect 298818 265961 298852 265989
rect 298880 265961 298914 265989
rect 298942 265961 298990 265989
rect -958 265913 298990 265961
rect -958 263175 298990 263223
rect -958 263147 -430 263175
rect -402 263147 -368 263175
rect -340 263147 -306 263175
rect -278 263147 -244 263175
rect -216 263147 2757 263175
rect 2785 263147 2819 263175
rect 2847 263147 2881 263175
rect 2909 263147 2943 263175
rect 2971 263147 18117 263175
rect 18145 263147 18179 263175
rect 18207 263147 18241 263175
rect 18269 263147 18303 263175
rect 18331 263147 33477 263175
rect 33505 263147 33539 263175
rect 33567 263147 33601 263175
rect 33629 263147 33663 263175
rect 33691 263147 48837 263175
rect 48865 263147 48899 263175
rect 48927 263147 48961 263175
rect 48989 263147 49023 263175
rect 49051 263147 64197 263175
rect 64225 263147 64259 263175
rect 64287 263147 64321 263175
rect 64349 263147 64383 263175
rect 64411 263147 79557 263175
rect 79585 263147 79619 263175
rect 79647 263147 79681 263175
rect 79709 263147 79743 263175
rect 79771 263147 94917 263175
rect 94945 263147 94979 263175
rect 95007 263147 95041 263175
rect 95069 263147 95103 263175
rect 95131 263147 110277 263175
rect 110305 263147 110339 263175
rect 110367 263147 110401 263175
rect 110429 263147 110463 263175
rect 110491 263147 125637 263175
rect 125665 263147 125699 263175
rect 125727 263147 125761 263175
rect 125789 263147 125823 263175
rect 125851 263147 140997 263175
rect 141025 263147 141059 263175
rect 141087 263147 141121 263175
rect 141149 263147 141183 263175
rect 141211 263147 156357 263175
rect 156385 263147 156419 263175
rect 156447 263147 156481 263175
rect 156509 263147 156543 263175
rect 156571 263147 171717 263175
rect 171745 263147 171779 263175
rect 171807 263147 171841 263175
rect 171869 263147 171903 263175
rect 171931 263147 187077 263175
rect 187105 263147 187139 263175
rect 187167 263147 187201 263175
rect 187229 263147 187263 263175
rect 187291 263147 202437 263175
rect 202465 263147 202499 263175
rect 202527 263147 202561 263175
rect 202589 263147 202623 263175
rect 202651 263147 217797 263175
rect 217825 263147 217859 263175
rect 217887 263147 217921 263175
rect 217949 263147 217983 263175
rect 218011 263147 233157 263175
rect 233185 263147 233219 263175
rect 233247 263147 233281 263175
rect 233309 263147 233343 263175
rect 233371 263147 248517 263175
rect 248545 263147 248579 263175
rect 248607 263147 248641 263175
rect 248669 263147 248703 263175
rect 248731 263147 263877 263175
rect 263905 263147 263939 263175
rect 263967 263147 264001 263175
rect 264029 263147 264063 263175
rect 264091 263147 279237 263175
rect 279265 263147 279299 263175
rect 279327 263147 279361 263175
rect 279389 263147 279423 263175
rect 279451 263147 294597 263175
rect 294625 263147 294659 263175
rect 294687 263147 294721 263175
rect 294749 263147 294783 263175
rect 294811 263147 298248 263175
rect 298276 263147 298310 263175
rect 298338 263147 298372 263175
rect 298400 263147 298434 263175
rect 298462 263147 298990 263175
rect -958 263113 298990 263147
rect -958 263085 -430 263113
rect -402 263085 -368 263113
rect -340 263085 -306 263113
rect -278 263085 -244 263113
rect -216 263085 2757 263113
rect 2785 263085 2819 263113
rect 2847 263085 2881 263113
rect 2909 263085 2943 263113
rect 2971 263085 18117 263113
rect 18145 263085 18179 263113
rect 18207 263085 18241 263113
rect 18269 263085 18303 263113
rect 18331 263085 33477 263113
rect 33505 263085 33539 263113
rect 33567 263085 33601 263113
rect 33629 263085 33663 263113
rect 33691 263085 48837 263113
rect 48865 263085 48899 263113
rect 48927 263085 48961 263113
rect 48989 263085 49023 263113
rect 49051 263085 64197 263113
rect 64225 263085 64259 263113
rect 64287 263085 64321 263113
rect 64349 263085 64383 263113
rect 64411 263085 79557 263113
rect 79585 263085 79619 263113
rect 79647 263085 79681 263113
rect 79709 263085 79743 263113
rect 79771 263085 94917 263113
rect 94945 263085 94979 263113
rect 95007 263085 95041 263113
rect 95069 263085 95103 263113
rect 95131 263085 110277 263113
rect 110305 263085 110339 263113
rect 110367 263085 110401 263113
rect 110429 263085 110463 263113
rect 110491 263085 125637 263113
rect 125665 263085 125699 263113
rect 125727 263085 125761 263113
rect 125789 263085 125823 263113
rect 125851 263085 140997 263113
rect 141025 263085 141059 263113
rect 141087 263085 141121 263113
rect 141149 263085 141183 263113
rect 141211 263085 156357 263113
rect 156385 263085 156419 263113
rect 156447 263085 156481 263113
rect 156509 263085 156543 263113
rect 156571 263085 171717 263113
rect 171745 263085 171779 263113
rect 171807 263085 171841 263113
rect 171869 263085 171903 263113
rect 171931 263085 187077 263113
rect 187105 263085 187139 263113
rect 187167 263085 187201 263113
rect 187229 263085 187263 263113
rect 187291 263085 202437 263113
rect 202465 263085 202499 263113
rect 202527 263085 202561 263113
rect 202589 263085 202623 263113
rect 202651 263085 217797 263113
rect 217825 263085 217859 263113
rect 217887 263085 217921 263113
rect 217949 263085 217983 263113
rect 218011 263085 233157 263113
rect 233185 263085 233219 263113
rect 233247 263085 233281 263113
rect 233309 263085 233343 263113
rect 233371 263085 248517 263113
rect 248545 263085 248579 263113
rect 248607 263085 248641 263113
rect 248669 263085 248703 263113
rect 248731 263085 263877 263113
rect 263905 263085 263939 263113
rect 263967 263085 264001 263113
rect 264029 263085 264063 263113
rect 264091 263085 279237 263113
rect 279265 263085 279299 263113
rect 279327 263085 279361 263113
rect 279389 263085 279423 263113
rect 279451 263085 294597 263113
rect 294625 263085 294659 263113
rect 294687 263085 294721 263113
rect 294749 263085 294783 263113
rect 294811 263085 298248 263113
rect 298276 263085 298310 263113
rect 298338 263085 298372 263113
rect 298400 263085 298434 263113
rect 298462 263085 298990 263113
rect -958 263051 298990 263085
rect -958 263023 -430 263051
rect -402 263023 -368 263051
rect -340 263023 -306 263051
rect -278 263023 -244 263051
rect -216 263023 2757 263051
rect 2785 263023 2819 263051
rect 2847 263023 2881 263051
rect 2909 263023 2943 263051
rect 2971 263023 18117 263051
rect 18145 263023 18179 263051
rect 18207 263023 18241 263051
rect 18269 263023 18303 263051
rect 18331 263023 33477 263051
rect 33505 263023 33539 263051
rect 33567 263023 33601 263051
rect 33629 263023 33663 263051
rect 33691 263023 48837 263051
rect 48865 263023 48899 263051
rect 48927 263023 48961 263051
rect 48989 263023 49023 263051
rect 49051 263023 64197 263051
rect 64225 263023 64259 263051
rect 64287 263023 64321 263051
rect 64349 263023 64383 263051
rect 64411 263023 79557 263051
rect 79585 263023 79619 263051
rect 79647 263023 79681 263051
rect 79709 263023 79743 263051
rect 79771 263023 94917 263051
rect 94945 263023 94979 263051
rect 95007 263023 95041 263051
rect 95069 263023 95103 263051
rect 95131 263023 110277 263051
rect 110305 263023 110339 263051
rect 110367 263023 110401 263051
rect 110429 263023 110463 263051
rect 110491 263023 125637 263051
rect 125665 263023 125699 263051
rect 125727 263023 125761 263051
rect 125789 263023 125823 263051
rect 125851 263023 140997 263051
rect 141025 263023 141059 263051
rect 141087 263023 141121 263051
rect 141149 263023 141183 263051
rect 141211 263023 156357 263051
rect 156385 263023 156419 263051
rect 156447 263023 156481 263051
rect 156509 263023 156543 263051
rect 156571 263023 171717 263051
rect 171745 263023 171779 263051
rect 171807 263023 171841 263051
rect 171869 263023 171903 263051
rect 171931 263023 187077 263051
rect 187105 263023 187139 263051
rect 187167 263023 187201 263051
rect 187229 263023 187263 263051
rect 187291 263023 202437 263051
rect 202465 263023 202499 263051
rect 202527 263023 202561 263051
rect 202589 263023 202623 263051
rect 202651 263023 217797 263051
rect 217825 263023 217859 263051
rect 217887 263023 217921 263051
rect 217949 263023 217983 263051
rect 218011 263023 233157 263051
rect 233185 263023 233219 263051
rect 233247 263023 233281 263051
rect 233309 263023 233343 263051
rect 233371 263023 248517 263051
rect 248545 263023 248579 263051
rect 248607 263023 248641 263051
rect 248669 263023 248703 263051
rect 248731 263023 263877 263051
rect 263905 263023 263939 263051
rect 263967 263023 264001 263051
rect 264029 263023 264063 263051
rect 264091 263023 279237 263051
rect 279265 263023 279299 263051
rect 279327 263023 279361 263051
rect 279389 263023 279423 263051
rect 279451 263023 294597 263051
rect 294625 263023 294659 263051
rect 294687 263023 294721 263051
rect 294749 263023 294783 263051
rect 294811 263023 298248 263051
rect 298276 263023 298310 263051
rect 298338 263023 298372 263051
rect 298400 263023 298434 263051
rect 298462 263023 298990 263051
rect -958 262989 298990 263023
rect -958 262961 -430 262989
rect -402 262961 -368 262989
rect -340 262961 -306 262989
rect -278 262961 -244 262989
rect -216 262961 2757 262989
rect 2785 262961 2819 262989
rect 2847 262961 2881 262989
rect 2909 262961 2943 262989
rect 2971 262961 18117 262989
rect 18145 262961 18179 262989
rect 18207 262961 18241 262989
rect 18269 262961 18303 262989
rect 18331 262961 33477 262989
rect 33505 262961 33539 262989
rect 33567 262961 33601 262989
rect 33629 262961 33663 262989
rect 33691 262961 48837 262989
rect 48865 262961 48899 262989
rect 48927 262961 48961 262989
rect 48989 262961 49023 262989
rect 49051 262961 64197 262989
rect 64225 262961 64259 262989
rect 64287 262961 64321 262989
rect 64349 262961 64383 262989
rect 64411 262961 79557 262989
rect 79585 262961 79619 262989
rect 79647 262961 79681 262989
rect 79709 262961 79743 262989
rect 79771 262961 94917 262989
rect 94945 262961 94979 262989
rect 95007 262961 95041 262989
rect 95069 262961 95103 262989
rect 95131 262961 110277 262989
rect 110305 262961 110339 262989
rect 110367 262961 110401 262989
rect 110429 262961 110463 262989
rect 110491 262961 125637 262989
rect 125665 262961 125699 262989
rect 125727 262961 125761 262989
rect 125789 262961 125823 262989
rect 125851 262961 140997 262989
rect 141025 262961 141059 262989
rect 141087 262961 141121 262989
rect 141149 262961 141183 262989
rect 141211 262961 156357 262989
rect 156385 262961 156419 262989
rect 156447 262961 156481 262989
rect 156509 262961 156543 262989
rect 156571 262961 171717 262989
rect 171745 262961 171779 262989
rect 171807 262961 171841 262989
rect 171869 262961 171903 262989
rect 171931 262961 187077 262989
rect 187105 262961 187139 262989
rect 187167 262961 187201 262989
rect 187229 262961 187263 262989
rect 187291 262961 202437 262989
rect 202465 262961 202499 262989
rect 202527 262961 202561 262989
rect 202589 262961 202623 262989
rect 202651 262961 217797 262989
rect 217825 262961 217859 262989
rect 217887 262961 217921 262989
rect 217949 262961 217983 262989
rect 218011 262961 233157 262989
rect 233185 262961 233219 262989
rect 233247 262961 233281 262989
rect 233309 262961 233343 262989
rect 233371 262961 248517 262989
rect 248545 262961 248579 262989
rect 248607 262961 248641 262989
rect 248669 262961 248703 262989
rect 248731 262961 263877 262989
rect 263905 262961 263939 262989
rect 263967 262961 264001 262989
rect 264029 262961 264063 262989
rect 264091 262961 279237 262989
rect 279265 262961 279299 262989
rect 279327 262961 279361 262989
rect 279389 262961 279423 262989
rect 279451 262961 294597 262989
rect 294625 262961 294659 262989
rect 294687 262961 294721 262989
rect 294749 262961 294783 262989
rect 294811 262961 298248 262989
rect 298276 262961 298310 262989
rect 298338 262961 298372 262989
rect 298400 262961 298434 262989
rect 298462 262961 298990 262989
rect -958 262913 298990 262961
rect -958 257175 298990 257223
rect -958 257147 -910 257175
rect -882 257147 -848 257175
rect -820 257147 -786 257175
rect -758 257147 -724 257175
rect -696 257147 4617 257175
rect 4645 257147 4679 257175
rect 4707 257147 4741 257175
rect 4769 257147 4803 257175
rect 4831 257147 19977 257175
rect 20005 257147 20039 257175
rect 20067 257147 20101 257175
rect 20129 257147 20163 257175
rect 20191 257147 35337 257175
rect 35365 257147 35399 257175
rect 35427 257147 35461 257175
rect 35489 257147 35523 257175
rect 35551 257147 50697 257175
rect 50725 257147 50759 257175
rect 50787 257147 50821 257175
rect 50849 257147 50883 257175
rect 50911 257147 66057 257175
rect 66085 257147 66119 257175
rect 66147 257147 66181 257175
rect 66209 257147 66243 257175
rect 66271 257147 81417 257175
rect 81445 257147 81479 257175
rect 81507 257147 81541 257175
rect 81569 257147 81603 257175
rect 81631 257147 96777 257175
rect 96805 257147 96839 257175
rect 96867 257147 96901 257175
rect 96929 257147 96963 257175
rect 96991 257147 112137 257175
rect 112165 257147 112199 257175
rect 112227 257147 112261 257175
rect 112289 257147 112323 257175
rect 112351 257147 127497 257175
rect 127525 257147 127559 257175
rect 127587 257147 127621 257175
rect 127649 257147 127683 257175
rect 127711 257147 142857 257175
rect 142885 257147 142919 257175
rect 142947 257147 142981 257175
rect 143009 257147 143043 257175
rect 143071 257147 158217 257175
rect 158245 257147 158279 257175
rect 158307 257147 158341 257175
rect 158369 257147 158403 257175
rect 158431 257147 173577 257175
rect 173605 257147 173639 257175
rect 173667 257147 173701 257175
rect 173729 257147 173763 257175
rect 173791 257147 188937 257175
rect 188965 257147 188999 257175
rect 189027 257147 189061 257175
rect 189089 257147 189123 257175
rect 189151 257147 204297 257175
rect 204325 257147 204359 257175
rect 204387 257147 204421 257175
rect 204449 257147 204483 257175
rect 204511 257147 219657 257175
rect 219685 257147 219719 257175
rect 219747 257147 219781 257175
rect 219809 257147 219843 257175
rect 219871 257147 235017 257175
rect 235045 257147 235079 257175
rect 235107 257147 235141 257175
rect 235169 257147 235203 257175
rect 235231 257147 250377 257175
rect 250405 257147 250439 257175
rect 250467 257147 250501 257175
rect 250529 257147 250563 257175
rect 250591 257147 265737 257175
rect 265765 257147 265799 257175
rect 265827 257147 265861 257175
rect 265889 257147 265923 257175
rect 265951 257147 281097 257175
rect 281125 257147 281159 257175
rect 281187 257147 281221 257175
rect 281249 257147 281283 257175
rect 281311 257147 296457 257175
rect 296485 257147 296519 257175
rect 296547 257147 296581 257175
rect 296609 257147 296643 257175
rect 296671 257147 298728 257175
rect 298756 257147 298790 257175
rect 298818 257147 298852 257175
rect 298880 257147 298914 257175
rect 298942 257147 298990 257175
rect -958 257113 298990 257147
rect -958 257085 -910 257113
rect -882 257085 -848 257113
rect -820 257085 -786 257113
rect -758 257085 -724 257113
rect -696 257085 4617 257113
rect 4645 257085 4679 257113
rect 4707 257085 4741 257113
rect 4769 257085 4803 257113
rect 4831 257085 19977 257113
rect 20005 257085 20039 257113
rect 20067 257085 20101 257113
rect 20129 257085 20163 257113
rect 20191 257085 35337 257113
rect 35365 257085 35399 257113
rect 35427 257085 35461 257113
rect 35489 257085 35523 257113
rect 35551 257085 50697 257113
rect 50725 257085 50759 257113
rect 50787 257085 50821 257113
rect 50849 257085 50883 257113
rect 50911 257085 66057 257113
rect 66085 257085 66119 257113
rect 66147 257085 66181 257113
rect 66209 257085 66243 257113
rect 66271 257085 81417 257113
rect 81445 257085 81479 257113
rect 81507 257085 81541 257113
rect 81569 257085 81603 257113
rect 81631 257085 96777 257113
rect 96805 257085 96839 257113
rect 96867 257085 96901 257113
rect 96929 257085 96963 257113
rect 96991 257085 112137 257113
rect 112165 257085 112199 257113
rect 112227 257085 112261 257113
rect 112289 257085 112323 257113
rect 112351 257085 127497 257113
rect 127525 257085 127559 257113
rect 127587 257085 127621 257113
rect 127649 257085 127683 257113
rect 127711 257085 142857 257113
rect 142885 257085 142919 257113
rect 142947 257085 142981 257113
rect 143009 257085 143043 257113
rect 143071 257085 158217 257113
rect 158245 257085 158279 257113
rect 158307 257085 158341 257113
rect 158369 257085 158403 257113
rect 158431 257085 173577 257113
rect 173605 257085 173639 257113
rect 173667 257085 173701 257113
rect 173729 257085 173763 257113
rect 173791 257085 188937 257113
rect 188965 257085 188999 257113
rect 189027 257085 189061 257113
rect 189089 257085 189123 257113
rect 189151 257085 204297 257113
rect 204325 257085 204359 257113
rect 204387 257085 204421 257113
rect 204449 257085 204483 257113
rect 204511 257085 219657 257113
rect 219685 257085 219719 257113
rect 219747 257085 219781 257113
rect 219809 257085 219843 257113
rect 219871 257085 235017 257113
rect 235045 257085 235079 257113
rect 235107 257085 235141 257113
rect 235169 257085 235203 257113
rect 235231 257085 250377 257113
rect 250405 257085 250439 257113
rect 250467 257085 250501 257113
rect 250529 257085 250563 257113
rect 250591 257085 265737 257113
rect 265765 257085 265799 257113
rect 265827 257085 265861 257113
rect 265889 257085 265923 257113
rect 265951 257085 281097 257113
rect 281125 257085 281159 257113
rect 281187 257085 281221 257113
rect 281249 257085 281283 257113
rect 281311 257085 296457 257113
rect 296485 257085 296519 257113
rect 296547 257085 296581 257113
rect 296609 257085 296643 257113
rect 296671 257085 298728 257113
rect 298756 257085 298790 257113
rect 298818 257085 298852 257113
rect 298880 257085 298914 257113
rect 298942 257085 298990 257113
rect -958 257051 298990 257085
rect -958 257023 -910 257051
rect -882 257023 -848 257051
rect -820 257023 -786 257051
rect -758 257023 -724 257051
rect -696 257023 4617 257051
rect 4645 257023 4679 257051
rect 4707 257023 4741 257051
rect 4769 257023 4803 257051
rect 4831 257023 19977 257051
rect 20005 257023 20039 257051
rect 20067 257023 20101 257051
rect 20129 257023 20163 257051
rect 20191 257023 35337 257051
rect 35365 257023 35399 257051
rect 35427 257023 35461 257051
rect 35489 257023 35523 257051
rect 35551 257023 50697 257051
rect 50725 257023 50759 257051
rect 50787 257023 50821 257051
rect 50849 257023 50883 257051
rect 50911 257023 66057 257051
rect 66085 257023 66119 257051
rect 66147 257023 66181 257051
rect 66209 257023 66243 257051
rect 66271 257023 81417 257051
rect 81445 257023 81479 257051
rect 81507 257023 81541 257051
rect 81569 257023 81603 257051
rect 81631 257023 96777 257051
rect 96805 257023 96839 257051
rect 96867 257023 96901 257051
rect 96929 257023 96963 257051
rect 96991 257023 112137 257051
rect 112165 257023 112199 257051
rect 112227 257023 112261 257051
rect 112289 257023 112323 257051
rect 112351 257023 127497 257051
rect 127525 257023 127559 257051
rect 127587 257023 127621 257051
rect 127649 257023 127683 257051
rect 127711 257023 142857 257051
rect 142885 257023 142919 257051
rect 142947 257023 142981 257051
rect 143009 257023 143043 257051
rect 143071 257023 158217 257051
rect 158245 257023 158279 257051
rect 158307 257023 158341 257051
rect 158369 257023 158403 257051
rect 158431 257023 173577 257051
rect 173605 257023 173639 257051
rect 173667 257023 173701 257051
rect 173729 257023 173763 257051
rect 173791 257023 188937 257051
rect 188965 257023 188999 257051
rect 189027 257023 189061 257051
rect 189089 257023 189123 257051
rect 189151 257023 204297 257051
rect 204325 257023 204359 257051
rect 204387 257023 204421 257051
rect 204449 257023 204483 257051
rect 204511 257023 219657 257051
rect 219685 257023 219719 257051
rect 219747 257023 219781 257051
rect 219809 257023 219843 257051
rect 219871 257023 235017 257051
rect 235045 257023 235079 257051
rect 235107 257023 235141 257051
rect 235169 257023 235203 257051
rect 235231 257023 250377 257051
rect 250405 257023 250439 257051
rect 250467 257023 250501 257051
rect 250529 257023 250563 257051
rect 250591 257023 265737 257051
rect 265765 257023 265799 257051
rect 265827 257023 265861 257051
rect 265889 257023 265923 257051
rect 265951 257023 281097 257051
rect 281125 257023 281159 257051
rect 281187 257023 281221 257051
rect 281249 257023 281283 257051
rect 281311 257023 296457 257051
rect 296485 257023 296519 257051
rect 296547 257023 296581 257051
rect 296609 257023 296643 257051
rect 296671 257023 298728 257051
rect 298756 257023 298790 257051
rect 298818 257023 298852 257051
rect 298880 257023 298914 257051
rect 298942 257023 298990 257051
rect -958 256989 298990 257023
rect -958 256961 -910 256989
rect -882 256961 -848 256989
rect -820 256961 -786 256989
rect -758 256961 -724 256989
rect -696 256961 4617 256989
rect 4645 256961 4679 256989
rect 4707 256961 4741 256989
rect 4769 256961 4803 256989
rect 4831 256961 19977 256989
rect 20005 256961 20039 256989
rect 20067 256961 20101 256989
rect 20129 256961 20163 256989
rect 20191 256961 35337 256989
rect 35365 256961 35399 256989
rect 35427 256961 35461 256989
rect 35489 256961 35523 256989
rect 35551 256961 50697 256989
rect 50725 256961 50759 256989
rect 50787 256961 50821 256989
rect 50849 256961 50883 256989
rect 50911 256961 66057 256989
rect 66085 256961 66119 256989
rect 66147 256961 66181 256989
rect 66209 256961 66243 256989
rect 66271 256961 81417 256989
rect 81445 256961 81479 256989
rect 81507 256961 81541 256989
rect 81569 256961 81603 256989
rect 81631 256961 96777 256989
rect 96805 256961 96839 256989
rect 96867 256961 96901 256989
rect 96929 256961 96963 256989
rect 96991 256961 112137 256989
rect 112165 256961 112199 256989
rect 112227 256961 112261 256989
rect 112289 256961 112323 256989
rect 112351 256961 127497 256989
rect 127525 256961 127559 256989
rect 127587 256961 127621 256989
rect 127649 256961 127683 256989
rect 127711 256961 142857 256989
rect 142885 256961 142919 256989
rect 142947 256961 142981 256989
rect 143009 256961 143043 256989
rect 143071 256961 158217 256989
rect 158245 256961 158279 256989
rect 158307 256961 158341 256989
rect 158369 256961 158403 256989
rect 158431 256961 173577 256989
rect 173605 256961 173639 256989
rect 173667 256961 173701 256989
rect 173729 256961 173763 256989
rect 173791 256961 188937 256989
rect 188965 256961 188999 256989
rect 189027 256961 189061 256989
rect 189089 256961 189123 256989
rect 189151 256961 204297 256989
rect 204325 256961 204359 256989
rect 204387 256961 204421 256989
rect 204449 256961 204483 256989
rect 204511 256961 219657 256989
rect 219685 256961 219719 256989
rect 219747 256961 219781 256989
rect 219809 256961 219843 256989
rect 219871 256961 235017 256989
rect 235045 256961 235079 256989
rect 235107 256961 235141 256989
rect 235169 256961 235203 256989
rect 235231 256961 250377 256989
rect 250405 256961 250439 256989
rect 250467 256961 250501 256989
rect 250529 256961 250563 256989
rect 250591 256961 265737 256989
rect 265765 256961 265799 256989
rect 265827 256961 265861 256989
rect 265889 256961 265923 256989
rect 265951 256961 281097 256989
rect 281125 256961 281159 256989
rect 281187 256961 281221 256989
rect 281249 256961 281283 256989
rect 281311 256961 296457 256989
rect 296485 256961 296519 256989
rect 296547 256961 296581 256989
rect 296609 256961 296643 256989
rect 296671 256961 298728 256989
rect 298756 256961 298790 256989
rect 298818 256961 298852 256989
rect 298880 256961 298914 256989
rect 298942 256961 298990 256989
rect -958 256913 298990 256961
rect -958 254175 298990 254223
rect -958 254147 -430 254175
rect -402 254147 -368 254175
rect -340 254147 -306 254175
rect -278 254147 -244 254175
rect -216 254147 2757 254175
rect 2785 254147 2819 254175
rect 2847 254147 2881 254175
rect 2909 254147 2943 254175
rect 2971 254147 18117 254175
rect 18145 254147 18179 254175
rect 18207 254147 18241 254175
rect 18269 254147 18303 254175
rect 18331 254147 33477 254175
rect 33505 254147 33539 254175
rect 33567 254147 33601 254175
rect 33629 254147 33663 254175
rect 33691 254147 48837 254175
rect 48865 254147 48899 254175
rect 48927 254147 48961 254175
rect 48989 254147 49023 254175
rect 49051 254147 64197 254175
rect 64225 254147 64259 254175
rect 64287 254147 64321 254175
rect 64349 254147 64383 254175
rect 64411 254147 79557 254175
rect 79585 254147 79619 254175
rect 79647 254147 79681 254175
rect 79709 254147 79743 254175
rect 79771 254147 94917 254175
rect 94945 254147 94979 254175
rect 95007 254147 95041 254175
rect 95069 254147 95103 254175
rect 95131 254147 110277 254175
rect 110305 254147 110339 254175
rect 110367 254147 110401 254175
rect 110429 254147 110463 254175
rect 110491 254147 125637 254175
rect 125665 254147 125699 254175
rect 125727 254147 125761 254175
rect 125789 254147 125823 254175
rect 125851 254147 140997 254175
rect 141025 254147 141059 254175
rect 141087 254147 141121 254175
rect 141149 254147 141183 254175
rect 141211 254147 156357 254175
rect 156385 254147 156419 254175
rect 156447 254147 156481 254175
rect 156509 254147 156543 254175
rect 156571 254147 171717 254175
rect 171745 254147 171779 254175
rect 171807 254147 171841 254175
rect 171869 254147 171903 254175
rect 171931 254147 187077 254175
rect 187105 254147 187139 254175
rect 187167 254147 187201 254175
rect 187229 254147 187263 254175
rect 187291 254147 202437 254175
rect 202465 254147 202499 254175
rect 202527 254147 202561 254175
rect 202589 254147 202623 254175
rect 202651 254147 217797 254175
rect 217825 254147 217859 254175
rect 217887 254147 217921 254175
rect 217949 254147 217983 254175
rect 218011 254147 233157 254175
rect 233185 254147 233219 254175
rect 233247 254147 233281 254175
rect 233309 254147 233343 254175
rect 233371 254147 248517 254175
rect 248545 254147 248579 254175
rect 248607 254147 248641 254175
rect 248669 254147 248703 254175
rect 248731 254147 263877 254175
rect 263905 254147 263939 254175
rect 263967 254147 264001 254175
rect 264029 254147 264063 254175
rect 264091 254147 279237 254175
rect 279265 254147 279299 254175
rect 279327 254147 279361 254175
rect 279389 254147 279423 254175
rect 279451 254147 294597 254175
rect 294625 254147 294659 254175
rect 294687 254147 294721 254175
rect 294749 254147 294783 254175
rect 294811 254147 298248 254175
rect 298276 254147 298310 254175
rect 298338 254147 298372 254175
rect 298400 254147 298434 254175
rect 298462 254147 298990 254175
rect -958 254113 298990 254147
rect -958 254085 -430 254113
rect -402 254085 -368 254113
rect -340 254085 -306 254113
rect -278 254085 -244 254113
rect -216 254085 2757 254113
rect 2785 254085 2819 254113
rect 2847 254085 2881 254113
rect 2909 254085 2943 254113
rect 2971 254085 18117 254113
rect 18145 254085 18179 254113
rect 18207 254085 18241 254113
rect 18269 254085 18303 254113
rect 18331 254085 33477 254113
rect 33505 254085 33539 254113
rect 33567 254085 33601 254113
rect 33629 254085 33663 254113
rect 33691 254085 48837 254113
rect 48865 254085 48899 254113
rect 48927 254085 48961 254113
rect 48989 254085 49023 254113
rect 49051 254085 64197 254113
rect 64225 254085 64259 254113
rect 64287 254085 64321 254113
rect 64349 254085 64383 254113
rect 64411 254085 79557 254113
rect 79585 254085 79619 254113
rect 79647 254085 79681 254113
rect 79709 254085 79743 254113
rect 79771 254085 94917 254113
rect 94945 254085 94979 254113
rect 95007 254085 95041 254113
rect 95069 254085 95103 254113
rect 95131 254085 110277 254113
rect 110305 254085 110339 254113
rect 110367 254085 110401 254113
rect 110429 254085 110463 254113
rect 110491 254085 125637 254113
rect 125665 254085 125699 254113
rect 125727 254085 125761 254113
rect 125789 254085 125823 254113
rect 125851 254085 140997 254113
rect 141025 254085 141059 254113
rect 141087 254085 141121 254113
rect 141149 254085 141183 254113
rect 141211 254085 156357 254113
rect 156385 254085 156419 254113
rect 156447 254085 156481 254113
rect 156509 254085 156543 254113
rect 156571 254085 171717 254113
rect 171745 254085 171779 254113
rect 171807 254085 171841 254113
rect 171869 254085 171903 254113
rect 171931 254085 187077 254113
rect 187105 254085 187139 254113
rect 187167 254085 187201 254113
rect 187229 254085 187263 254113
rect 187291 254085 202437 254113
rect 202465 254085 202499 254113
rect 202527 254085 202561 254113
rect 202589 254085 202623 254113
rect 202651 254085 217797 254113
rect 217825 254085 217859 254113
rect 217887 254085 217921 254113
rect 217949 254085 217983 254113
rect 218011 254085 233157 254113
rect 233185 254085 233219 254113
rect 233247 254085 233281 254113
rect 233309 254085 233343 254113
rect 233371 254085 248517 254113
rect 248545 254085 248579 254113
rect 248607 254085 248641 254113
rect 248669 254085 248703 254113
rect 248731 254085 263877 254113
rect 263905 254085 263939 254113
rect 263967 254085 264001 254113
rect 264029 254085 264063 254113
rect 264091 254085 279237 254113
rect 279265 254085 279299 254113
rect 279327 254085 279361 254113
rect 279389 254085 279423 254113
rect 279451 254085 294597 254113
rect 294625 254085 294659 254113
rect 294687 254085 294721 254113
rect 294749 254085 294783 254113
rect 294811 254085 298248 254113
rect 298276 254085 298310 254113
rect 298338 254085 298372 254113
rect 298400 254085 298434 254113
rect 298462 254085 298990 254113
rect -958 254051 298990 254085
rect -958 254023 -430 254051
rect -402 254023 -368 254051
rect -340 254023 -306 254051
rect -278 254023 -244 254051
rect -216 254023 2757 254051
rect 2785 254023 2819 254051
rect 2847 254023 2881 254051
rect 2909 254023 2943 254051
rect 2971 254023 18117 254051
rect 18145 254023 18179 254051
rect 18207 254023 18241 254051
rect 18269 254023 18303 254051
rect 18331 254023 33477 254051
rect 33505 254023 33539 254051
rect 33567 254023 33601 254051
rect 33629 254023 33663 254051
rect 33691 254023 48837 254051
rect 48865 254023 48899 254051
rect 48927 254023 48961 254051
rect 48989 254023 49023 254051
rect 49051 254023 64197 254051
rect 64225 254023 64259 254051
rect 64287 254023 64321 254051
rect 64349 254023 64383 254051
rect 64411 254023 79557 254051
rect 79585 254023 79619 254051
rect 79647 254023 79681 254051
rect 79709 254023 79743 254051
rect 79771 254023 94917 254051
rect 94945 254023 94979 254051
rect 95007 254023 95041 254051
rect 95069 254023 95103 254051
rect 95131 254023 110277 254051
rect 110305 254023 110339 254051
rect 110367 254023 110401 254051
rect 110429 254023 110463 254051
rect 110491 254023 125637 254051
rect 125665 254023 125699 254051
rect 125727 254023 125761 254051
rect 125789 254023 125823 254051
rect 125851 254023 140997 254051
rect 141025 254023 141059 254051
rect 141087 254023 141121 254051
rect 141149 254023 141183 254051
rect 141211 254023 156357 254051
rect 156385 254023 156419 254051
rect 156447 254023 156481 254051
rect 156509 254023 156543 254051
rect 156571 254023 171717 254051
rect 171745 254023 171779 254051
rect 171807 254023 171841 254051
rect 171869 254023 171903 254051
rect 171931 254023 187077 254051
rect 187105 254023 187139 254051
rect 187167 254023 187201 254051
rect 187229 254023 187263 254051
rect 187291 254023 202437 254051
rect 202465 254023 202499 254051
rect 202527 254023 202561 254051
rect 202589 254023 202623 254051
rect 202651 254023 217797 254051
rect 217825 254023 217859 254051
rect 217887 254023 217921 254051
rect 217949 254023 217983 254051
rect 218011 254023 233157 254051
rect 233185 254023 233219 254051
rect 233247 254023 233281 254051
rect 233309 254023 233343 254051
rect 233371 254023 248517 254051
rect 248545 254023 248579 254051
rect 248607 254023 248641 254051
rect 248669 254023 248703 254051
rect 248731 254023 263877 254051
rect 263905 254023 263939 254051
rect 263967 254023 264001 254051
rect 264029 254023 264063 254051
rect 264091 254023 279237 254051
rect 279265 254023 279299 254051
rect 279327 254023 279361 254051
rect 279389 254023 279423 254051
rect 279451 254023 294597 254051
rect 294625 254023 294659 254051
rect 294687 254023 294721 254051
rect 294749 254023 294783 254051
rect 294811 254023 298248 254051
rect 298276 254023 298310 254051
rect 298338 254023 298372 254051
rect 298400 254023 298434 254051
rect 298462 254023 298990 254051
rect -958 253989 298990 254023
rect -958 253961 -430 253989
rect -402 253961 -368 253989
rect -340 253961 -306 253989
rect -278 253961 -244 253989
rect -216 253961 2757 253989
rect 2785 253961 2819 253989
rect 2847 253961 2881 253989
rect 2909 253961 2943 253989
rect 2971 253961 18117 253989
rect 18145 253961 18179 253989
rect 18207 253961 18241 253989
rect 18269 253961 18303 253989
rect 18331 253961 33477 253989
rect 33505 253961 33539 253989
rect 33567 253961 33601 253989
rect 33629 253961 33663 253989
rect 33691 253961 48837 253989
rect 48865 253961 48899 253989
rect 48927 253961 48961 253989
rect 48989 253961 49023 253989
rect 49051 253961 64197 253989
rect 64225 253961 64259 253989
rect 64287 253961 64321 253989
rect 64349 253961 64383 253989
rect 64411 253961 79557 253989
rect 79585 253961 79619 253989
rect 79647 253961 79681 253989
rect 79709 253961 79743 253989
rect 79771 253961 94917 253989
rect 94945 253961 94979 253989
rect 95007 253961 95041 253989
rect 95069 253961 95103 253989
rect 95131 253961 110277 253989
rect 110305 253961 110339 253989
rect 110367 253961 110401 253989
rect 110429 253961 110463 253989
rect 110491 253961 125637 253989
rect 125665 253961 125699 253989
rect 125727 253961 125761 253989
rect 125789 253961 125823 253989
rect 125851 253961 140997 253989
rect 141025 253961 141059 253989
rect 141087 253961 141121 253989
rect 141149 253961 141183 253989
rect 141211 253961 156357 253989
rect 156385 253961 156419 253989
rect 156447 253961 156481 253989
rect 156509 253961 156543 253989
rect 156571 253961 171717 253989
rect 171745 253961 171779 253989
rect 171807 253961 171841 253989
rect 171869 253961 171903 253989
rect 171931 253961 187077 253989
rect 187105 253961 187139 253989
rect 187167 253961 187201 253989
rect 187229 253961 187263 253989
rect 187291 253961 202437 253989
rect 202465 253961 202499 253989
rect 202527 253961 202561 253989
rect 202589 253961 202623 253989
rect 202651 253961 217797 253989
rect 217825 253961 217859 253989
rect 217887 253961 217921 253989
rect 217949 253961 217983 253989
rect 218011 253961 233157 253989
rect 233185 253961 233219 253989
rect 233247 253961 233281 253989
rect 233309 253961 233343 253989
rect 233371 253961 248517 253989
rect 248545 253961 248579 253989
rect 248607 253961 248641 253989
rect 248669 253961 248703 253989
rect 248731 253961 263877 253989
rect 263905 253961 263939 253989
rect 263967 253961 264001 253989
rect 264029 253961 264063 253989
rect 264091 253961 279237 253989
rect 279265 253961 279299 253989
rect 279327 253961 279361 253989
rect 279389 253961 279423 253989
rect 279451 253961 294597 253989
rect 294625 253961 294659 253989
rect 294687 253961 294721 253989
rect 294749 253961 294783 253989
rect 294811 253961 298248 253989
rect 298276 253961 298310 253989
rect 298338 253961 298372 253989
rect 298400 253961 298434 253989
rect 298462 253961 298990 253989
rect -958 253913 298990 253961
rect -958 248175 298990 248223
rect -958 248147 -910 248175
rect -882 248147 -848 248175
rect -820 248147 -786 248175
rect -758 248147 -724 248175
rect -696 248147 4617 248175
rect 4645 248147 4679 248175
rect 4707 248147 4741 248175
rect 4769 248147 4803 248175
rect 4831 248147 19977 248175
rect 20005 248147 20039 248175
rect 20067 248147 20101 248175
rect 20129 248147 20163 248175
rect 20191 248147 35337 248175
rect 35365 248147 35399 248175
rect 35427 248147 35461 248175
rect 35489 248147 35523 248175
rect 35551 248147 50697 248175
rect 50725 248147 50759 248175
rect 50787 248147 50821 248175
rect 50849 248147 50883 248175
rect 50911 248147 66057 248175
rect 66085 248147 66119 248175
rect 66147 248147 66181 248175
rect 66209 248147 66243 248175
rect 66271 248147 81417 248175
rect 81445 248147 81479 248175
rect 81507 248147 81541 248175
rect 81569 248147 81603 248175
rect 81631 248147 96777 248175
rect 96805 248147 96839 248175
rect 96867 248147 96901 248175
rect 96929 248147 96963 248175
rect 96991 248147 112137 248175
rect 112165 248147 112199 248175
rect 112227 248147 112261 248175
rect 112289 248147 112323 248175
rect 112351 248147 127497 248175
rect 127525 248147 127559 248175
rect 127587 248147 127621 248175
rect 127649 248147 127683 248175
rect 127711 248147 142857 248175
rect 142885 248147 142919 248175
rect 142947 248147 142981 248175
rect 143009 248147 143043 248175
rect 143071 248147 158217 248175
rect 158245 248147 158279 248175
rect 158307 248147 158341 248175
rect 158369 248147 158403 248175
rect 158431 248147 173577 248175
rect 173605 248147 173639 248175
rect 173667 248147 173701 248175
rect 173729 248147 173763 248175
rect 173791 248147 188937 248175
rect 188965 248147 188999 248175
rect 189027 248147 189061 248175
rect 189089 248147 189123 248175
rect 189151 248147 204297 248175
rect 204325 248147 204359 248175
rect 204387 248147 204421 248175
rect 204449 248147 204483 248175
rect 204511 248147 219657 248175
rect 219685 248147 219719 248175
rect 219747 248147 219781 248175
rect 219809 248147 219843 248175
rect 219871 248147 235017 248175
rect 235045 248147 235079 248175
rect 235107 248147 235141 248175
rect 235169 248147 235203 248175
rect 235231 248147 250377 248175
rect 250405 248147 250439 248175
rect 250467 248147 250501 248175
rect 250529 248147 250563 248175
rect 250591 248147 265737 248175
rect 265765 248147 265799 248175
rect 265827 248147 265861 248175
rect 265889 248147 265923 248175
rect 265951 248147 281097 248175
rect 281125 248147 281159 248175
rect 281187 248147 281221 248175
rect 281249 248147 281283 248175
rect 281311 248147 296457 248175
rect 296485 248147 296519 248175
rect 296547 248147 296581 248175
rect 296609 248147 296643 248175
rect 296671 248147 298728 248175
rect 298756 248147 298790 248175
rect 298818 248147 298852 248175
rect 298880 248147 298914 248175
rect 298942 248147 298990 248175
rect -958 248113 298990 248147
rect -958 248085 -910 248113
rect -882 248085 -848 248113
rect -820 248085 -786 248113
rect -758 248085 -724 248113
rect -696 248085 4617 248113
rect 4645 248085 4679 248113
rect 4707 248085 4741 248113
rect 4769 248085 4803 248113
rect 4831 248085 19977 248113
rect 20005 248085 20039 248113
rect 20067 248085 20101 248113
rect 20129 248085 20163 248113
rect 20191 248085 35337 248113
rect 35365 248085 35399 248113
rect 35427 248085 35461 248113
rect 35489 248085 35523 248113
rect 35551 248085 50697 248113
rect 50725 248085 50759 248113
rect 50787 248085 50821 248113
rect 50849 248085 50883 248113
rect 50911 248085 66057 248113
rect 66085 248085 66119 248113
rect 66147 248085 66181 248113
rect 66209 248085 66243 248113
rect 66271 248085 81417 248113
rect 81445 248085 81479 248113
rect 81507 248085 81541 248113
rect 81569 248085 81603 248113
rect 81631 248085 96777 248113
rect 96805 248085 96839 248113
rect 96867 248085 96901 248113
rect 96929 248085 96963 248113
rect 96991 248085 112137 248113
rect 112165 248085 112199 248113
rect 112227 248085 112261 248113
rect 112289 248085 112323 248113
rect 112351 248085 127497 248113
rect 127525 248085 127559 248113
rect 127587 248085 127621 248113
rect 127649 248085 127683 248113
rect 127711 248085 142857 248113
rect 142885 248085 142919 248113
rect 142947 248085 142981 248113
rect 143009 248085 143043 248113
rect 143071 248085 158217 248113
rect 158245 248085 158279 248113
rect 158307 248085 158341 248113
rect 158369 248085 158403 248113
rect 158431 248085 173577 248113
rect 173605 248085 173639 248113
rect 173667 248085 173701 248113
rect 173729 248085 173763 248113
rect 173791 248085 188937 248113
rect 188965 248085 188999 248113
rect 189027 248085 189061 248113
rect 189089 248085 189123 248113
rect 189151 248085 204297 248113
rect 204325 248085 204359 248113
rect 204387 248085 204421 248113
rect 204449 248085 204483 248113
rect 204511 248085 219657 248113
rect 219685 248085 219719 248113
rect 219747 248085 219781 248113
rect 219809 248085 219843 248113
rect 219871 248085 235017 248113
rect 235045 248085 235079 248113
rect 235107 248085 235141 248113
rect 235169 248085 235203 248113
rect 235231 248085 250377 248113
rect 250405 248085 250439 248113
rect 250467 248085 250501 248113
rect 250529 248085 250563 248113
rect 250591 248085 265737 248113
rect 265765 248085 265799 248113
rect 265827 248085 265861 248113
rect 265889 248085 265923 248113
rect 265951 248085 281097 248113
rect 281125 248085 281159 248113
rect 281187 248085 281221 248113
rect 281249 248085 281283 248113
rect 281311 248085 296457 248113
rect 296485 248085 296519 248113
rect 296547 248085 296581 248113
rect 296609 248085 296643 248113
rect 296671 248085 298728 248113
rect 298756 248085 298790 248113
rect 298818 248085 298852 248113
rect 298880 248085 298914 248113
rect 298942 248085 298990 248113
rect -958 248051 298990 248085
rect -958 248023 -910 248051
rect -882 248023 -848 248051
rect -820 248023 -786 248051
rect -758 248023 -724 248051
rect -696 248023 4617 248051
rect 4645 248023 4679 248051
rect 4707 248023 4741 248051
rect 4769 248023 4803 248051
rect 4831 248023 19977 248051
rect 20005 248023 20039 248051
rect 20067 248023 20101 248051
rect 20129 248023 20163 248051
rect 20191 248023 35337 248051
rect 35365 248023 35399 248051
rect 35427 248023 35461 248051
rect 35489 248023 35523 248051
rect 35551 248023 50697 248051
rect 50725 248023 50759 248051
rect 50787 248023 50821 248051
rect 50849 248023 50883 248051
rect 50911 248023 66057 248051
rect 66085 248023 66119 248051
rect 66147 248023 66181 248051
rect 66209 248023 66243 248051
rect 66271 248023 81417 248051
rect 81445 248023 81479 248051
rect 81507 248023 81541 248051
rect 81569 248023 81603 248051
rect 81631 248023 96777 248051
rect 96805 248023 96839 248051
rect 96867 248023 96901 248051
rect 96929 248023 96963 248051
rect 96991 248023 112137 248051
rect 112165 248023 112199 248051
rect 112227 248023 112261 248051
rect 112289 248023 112323 248051
rect 112351 248023 127497 248051
rect 127525 248023 127559 248051
rect 127587 248023 127621 248051
rect 127649 248023 127683 248051
rect 127711 248023 142857 248051
rect 142885 248023 142919 248051
rect 142947 248023 142981 248051
rect 143009 248023 143043 248051
rect 143071 248023 158217 248051
rect 158245 248023 158279 248051
rect 158307 248023 158341 248051
rect 158369 248023 158403 248051
rect 158431 248023 173577 248051
rect 173605 248023 173639 248051
rect 173667 248023 173701 248051
rect 173729 248023 173763 248051
rect 173791 248023 188937 248051
rect 188965 248023 188999 248051
rect 189027 248023 189061 248051
rect 189089 248023 189123 248051
rect 189151 248023 204297 248051
rect 204325 248023 204359 248051
rect 204387 248023 204421 248051
rect 204449 248023 204483 248051
rect 204511 248023 219657 248051
rect 219685 248023 219719 248051
rect 219747 248023 219781 248051
rect 219809 248023 219843 248051
rect 219871 248023 235017 248051
rect 235045 248023 235079 248051
rect 235107 248023 235141 248051
rect 235169 248023 235203 248051
rect 235231 248023 250377 248051
rect 250405 248023 250439 248051
rect 250467 248023 250501 248051
rect 250529 248023 250563 248051
rect 250591 248023 265737 248051
rect 265765 248023 265799 248051
rect 265827 248023 265861 248051
rect 265889 248023 265923 248051
rect 265951 248023 281097 248051
rect 281125 248023 281159 248051
rect 281187 248023 281221 248051
rect 281249 248023 281283 248051
rect 281311 248023 296457 248051
rect 296485 248023 296519 248051
rect 296547 248023 296581 248051
rect 296609 248023 296643 248051
rect 296671 248023 298728 248051
rect 298756 248023 298790 248051
rect 298818 248023 298852 248051
rect 298880 248023 298914 248051
rect 298942 248023 298990 248051
rect -958 247989 298990 248023
rect -958 247961 -910 247989
rect -882 247961 -848 247989
rect -820 247961 -786 247989
rect -758 247961 -724 247989
rect -696 247961 4617 247989
rect 4645 247961 4679 247989
rect 4707 247961 4741 247989
rect 4769 247961 4803 247989
rect 4831 247961 19977 247989
rect 20005 247961 20039 247989
rect 20067 247961 20101 247989
rect 20129 247961 20163 247989
rect 20191 247961 35337 247989
rect 35365 247961 35399 247989
rect 35427 247961 35461 247989
rect 35489 247961 35523 247989
rect 35551 247961 50697 247989
rect 50725 247961 50759 247989
rect 50787 247961 50821 247989
rect 50849 247961 50883 247989
rect 50911 247961 66057 247989
rect 66085 247961 66119 247989
rect 66147 247961 66181 247989
rect 66209 247961 66243 247989
rect 66271 247961 81417 247989
rect 81445 247961 81479 247989
rect 81507 247961 81541 247989
rect 81569 247961 81603 247989
rect 81631 247961 96777 247989
rect 96805 247961 96839 247989
rect 96867 247961 96901 247989
rect 96929 247961 96963 247989
rect 96991 247961 112137 247989
rect 112165 247961 112199 247989
rect 112227 247961 112261 247989
rect 112289 247961 112323 247989
rect 112351 247961 127497 247989
rect 127525 247961 127559 247989
rect 127587 247961 127621 247989
rect 127649 247961 127683 247989
rect 127711 247961 142857 247989
rect 142885 247961 142919 247989
rect 142947 247961 142981 247989
rect 143009 247961 143043 247989
rect 143071 247961 158217 247989
rect 158245 247961 158279 247989
rect 158307 247961 158341 247989
rect 158369 247961 158403 247989
rect 158431 247961 173577 247989
rect 173605 247961 173639 247989
rect 173667 247961 173701 247989
rect 173729 247961 173763 247989
rect 173791 247961 188937 247989
rect 188965 247961 188999 247989
rect 189027 247961 189061 247989
rect 189089 247961 189123 247989
rect 189151 247961 204297 247989
rect 204325 247961 204359 247989
rect 204387 247961 204421 247989
rect 204449 247961 204483 247989
rect 204511 247961 219657 247989
rect 219685 247961 219719 247989
rect 219747 247961 219781 247989
rect 219809 247961 219843 247989
rect 219871 247961 235017 247989
rect 235045 247961 235079 247989
rect 235107 247961 235141 247989
rect 235169 247961 235203 247989
rect 235231 247961 250377 247989
rect 250405 247961 250439 247989
rect 250467 247961 250501 247989
rect 250529 247961 250563 247989
rect 250591 247961 265737 247989
rect 265765 247961 265799 247989
rect 265827 247961 265861 247989
rect 265889 247961 265923 247989
rect 265951 247961 281097 247989
rect 281125 247961 281159 247989
rect 281187 247961 281221 247989
rect 281249 247961 281283 247989
rect 281311 247961 296457 247989
rect 296485 247961 296519 247989
rect 296547 247961 296581 247989
rect 296609 247961 296643 247989
rect 296671 247961 298728 247989
rect 298756 247961 298790 247989
rect 298818 247961 298852 247989
rect 298880 247961 298914 247989
rect 298942 247961 298990 247989
rect -958 247913 298990 247961
rect -958 245175 298990 245223
rect -958 245147 -430 245175
rect -402 245147 -368 245175
rect -340 245147 -306 245175
rect -278 245147 -244 245175
rect -216 245147 2757 245175
rect 2785 245147 2819 245175
rect 2847 245147 2881 245175
rect 2909 245147 2943 245175
rect 2971 245147 18117 245175
rect 18145 245147 18179 245175
rect 18207 245147 18241 245175
rect 18269 245147 18303 245175
rect 18331 245147 33477 245175
rect 33505 245147 33539 245175
rect 33567 245147 33601 245175
rect 33629 245147 33663 245175
rect 33691 245147 48837 245175
rect 48865 245147 48899 245175
rect 48927 245147 48961 245175
rect 48989 245147 49023 245175
rect 49051 245147 64197 245175
rect 64225 245147 64259 245175
rect 64287 245147 64321 245175
rect 64349 245147 64383 245175
rect 64411 245147 79557 245175
rect 79585 245147 79619 245175
rect 79647 245147 79681 245175
rect 79709 245147 79743 245175
rect 79771 245147 94917 245175
rect 94945 245147 94979 245175
rect 95007 245147 95041 245175
rect 95069 245147 95103 245175
rect 95131 245147 110277 245175
rect 110305 245147 110339 245175
rect 110367 245147 110401 245175
rect 110429 245147 110463 245175
rect 110491 245147 125637 245175
rect 125665 245147 125699 245175
rect 125727 245147 125761 245175
rect 125789 245147 125823 245175
rect 125851 245147 140997 245175
rect 141025 245147 141059 245175
rect 141087 245147 141121 245175
rect 141149 245147 141183 245175
rect 141211 245147 156357 245175
rect 156385 245147 156419 245175
rect 156447 245147 156481 245175
rect 156509 245147 156543 245175
rect 156571 245147 171717 245175
rect 171745 245147 171779 245175
rect 171807 245147 171841 245175
rect 171869 245147 171903 245175
rect 171931 245147 187077 245175
rect 187105 245147 187139 245175
rect 187167 245147 187201 245175
rect 187229 245147 187263 245175
rect 187291 245147 202437 245175
rect 202465 245147 202499 245175
rect 202527 245147 202561 245175
rect 202589 245147 202623 245175
rect 202651 245147 217797 245175
rect 217825 245147 217859 245175
rect 217887 245147 217921 245175
rect 217949 245147 217983 245175
rect 218011 245147 233157 245175
rect 233185 245147 233219 245175
rect 233247 245147 233281 245175
rect 233309 245147 233343 245175
rect 233371 245147 248517 245175
rect 248545 245147 248579 245175
rect 248607 245147 248641 245175
rect 248669 245147 248703 245175
rect 248731 245147 263877 245175
rect 263905 245147 263939 245175
rect 263967 245147 264001 245175
rect 264029 245147 264063 245175
rect 264091 245147 279237 245175
rect 279265 245147 279299 245175
rect 279327 245147 279361 245175
rect 279389 245147 279423 245175
rect 279451 245147 294597 245175
rect 294625 245147 294659 245175
rect 294687 245147 294721 245175
rect 294749 245147 294783 245175
rect 294811 245147 298248 245175
rect 298276 245147 298310 245175
rect 298338 245147 298372 245175
rect 298400 245147 298434 245175
rect 298462 245147 298990 245175
rect -958 245113 298990 245147
rect -958 245085 -430 245113
rect -402 245085 -368 245113
rect -340 245085 -306 245113
rect -278 245085 -244 245113
rect -216 245085 2757 245113
rect 2785 245085 2819 245113
rect 2847 245085 2881 245113
rect 2909 245085 2943 245113
rect 2971 245085 18117 245113
rect 18145 245085 18179 245113
rect 18207 245085 18241 245113
rect 18269 245085 18303 245113
rect 18331 245085 33477 245113
rect 33505 245085 33539 245113
rect 33567 245085 33601 245113
rect 33629 245085 33663 245113
rect 33691 245085 48837 245113
rect 48865 245085 48899 245113
rect 48927 245085 48961 245113
rect 48989 245085 49023 245113
rect 49051 245085 64197 245113
rect 64225 245085 64259 245113
rect 64287 245085 64321 245113
rect 64349 245085 64383 245113
rect 64411 245085 79557 245113
rect 79585 245085 79619 245113
rect 79647 245085 79681 245113
rect 79709 245085 79743 245113
rect 79771 245085 94917 245113
rect 94945 245085 94979 245113
rect 95007 245085 95041 245113
rect 95069 245085 95103 245113
rect 95131 245085 110277 245113
rect 110305 245085 110339 245113
rect 110367 245085 110401 245113
rect 110429 245085 110463 245113
rect 110491 245085 125637 245113
rect 125665 245085 125699 245113
rect 125727 245085 125761 245113
rect 125789 245085 125823 245113
rect 125851 245085 140997 245113
rect 141025 245085 141059 245113
rect 141087 245085 141121 245113
rect 141149 245085 141183 245113
rect 141211 245085 156357 245113
rect 156385 245085 156419 245113
rect 156447 245085 156481 245113
rect 156509 245085 156543 245113
rect 156571 245085 171717 245113
rect 171745 245085 171779 245113
rect 171807 245085 171841 245113
rect 171869 245085 171903 245113
rect 171931 245085 187077 245113
rect 187105 245085 187139 245113
rect 187167 245085 187201 245113
rect 187229 245085 187263 245113
rect 187291 245085 202437 245113
rect 202465 245085 202499 245113
rect 202527 245085 202561 245113
rect 202589 245085 202623 245113
rect 202651 245085 217797 245113
rect 217825 245085 217859 245113
rect 217887 245085 217921 245113
rect 217949 245085 217983 245113
rect 218011 245085 233157 245113
rect 233185 245085 233219 245113
rect 233247 245085 233281 245113
rect 233309 245085 233343 245113
rect 233371 245085 248517 245113
rect 248545 245085 248579 245113
rect 248607 245085 248641 245113
rect 248669 245085 248703 245113
rect 248731 245085 263877 245113
rect 263905 245085 263939 245113
rect 263967 245085 264001 245113
rect 264029 245085 264063 245113
rect 264091 245085 279237 245113
rect 279265 245085 279299 245113
rect 279327 245085 279361 245113
rect 279389 245085 279423 245113
rect 279451 245085 294597 245113
rect 294625 245085 294659 245113
rect 294687 245085 294721 245113
rect 294749 245085 294783 245113
rect 294811 245085 298248 245113
rect 298276 245085 298310 245113
rect 298338 245085 298372 245113
rect 298400 245085 298434 245113
rect 298462 245085 298990 245113
rect -958 245051 298990 245085
rect -958 245023 -430 245051
rect -402 245023 -368 245051
rect -340 245023 -306 245051
rect -278 245023 -244 245051
rect -216 245023 2757 245051
rect 2785 245023 2819 245051
rect 2847 245023 2881 245051
rect 2909 245023 2943 245051
rect 2971 245023 18117 245051
rect 18145 245023 18179 245051
rect 18207 245023 18241 245051
rect 18269 245023 18303 245051
rect 18331 245023 33477 245051
rect 33505 245023 33539 245051
rect 33567 245023 33601 245051
rect 33629 245023 33663 245051
rect 33691 245023 48837 245051
rect 48865 245023 48899 245051
rect 48927 245023 48961 245051
rect 48989 245023 49023 245051
rect 49051 245023 64197 245051
rect 64225 245023 64259 245051
rect 64287 245023 64321 245051
rect 64349 245023 64383 245051
rect 64411 245023 79557 245051
rect 79585 245023 79619 245051
rect 79647 245023 79681 245051
rect 79709 245023 79743 245051
rect 79771 245023 94917 245051
rect 94945 245023 94979 245051
rect 95007 245023 95041 245051
rect 95069 245023 95103 245051
rect 95131 245023 110277 245051
rect 110305 245023 110339 245051
rect 110367 245023 110401 245051
rect 110429 245023 110463 245051
rect 110491 245023 125637 245051
rect 125665 245023 125699 245051
rect 125727 245023 125761 245051
rect 125789 245023 125823 245051
rect 125851 245023 140997 245051
rect 141025 245023 141059 245051
rect 141087 245023 141121 245051
rect 141149 245023 141183 245051
rect 141211 245023 156357 245051
rect 156385 245023 156419 245051
rect 156447 245023 156481 245051
rect 156509 245023 156543 245051
rect 156571 245023 171717 245051
rect 171745 245023 171779 245051
rect 171807 245023 171841 245051
rect 171869 245023 171903 245051
rect 171931 245023 187077 245051
rect 187105 245023 187139 245051
rect 187167 245023 187201 245051
rect 187229 245023 187263 245051
rect 187291 245023 202437 245051
rect 202465 245023 202499 245051
rect 202527 245023 202561 245051
rect 202589 245023 202623 245051
rect 202651 245023 217797 245051
rect 217825 245023 217859 245051
rect 217887 245023 217921 245051
rect 217949 245023 217983 245051
rect 218011 245023 233157 245051
rect 233185 245023 233219 245051
rect 233247 245023 233281 245051
rect 233309 245023 233343 245051
rect 233371 245023 248517 245051
rect 248545 245023 248579 245051
rect 248607 245023 248641 245051
rect 248669 245023 248703 245051
rect 248731 245023 263877 245051
rect 263905 245023 263939 245051
rect 263967 245023 264001 245051
rect 264029 245023 264063 245051
rect 264091 245023 279237 245051
rect 279265 245023 279299 245051
rect 279327 245023 279361 245051
rect 279389 245023 279423 245051
rect 279451 245023 294597 245051
rect 294625 245023 294659 245051
rect 294687 245023 294721 245051
rect 294749 245023 294783 245051
rect 294811 245023 298248 245051
rect 298276 245023 298310 245051
rect 298338 245023 298372 245051
rect 298400 245023 298434 245051
rect 298462 245023 298990 245051
rect -958 244989 298990 245023
rect -958 244961 -430 244989
rect -402 244961 -368 244989
rect -340 244961 -306 244989
rect -278 244961 -244 244989
rect -216 244961 2757 244989
rect 2785 244961 2819 244989
rect 2847 244961 2881 244989
rect 2909 244961 2943 244989
rect 2971 244961 18117 244989
rect 18145 244961 18179 244989
rect 18207 244961 18241 244989
rect 18269 244961 18303 244989
rect 18331 244961 33477 244989
rect 33505 244961 33539 244989
rect 33567 244961 33601 244989
rect 33629 244961 33663 244989
rect 33691 244961 48837 244989
rect 48865 244961 48899 244989
rect 48927 244961 48961 244989
rect 48989 244961 49023 244989
rect 49051 244961 64197 244989
rect 64225 244961 64259 244989
rect 64287 244961 64321 244989
rect 64349 244961 64383 244989
rect 64411 244961 79557 244989
rect 79585 244961 79619 244989
rect 79647 244961 79681 244989
rect 79709 244961 79743 244989
rect 79771 244961 94917 244989
rect 94945 244961 94979 244989
rect 95007 244961 95041 244989
rect 95069 244961 95103 244989
rect 95131 244961 110277 244989
rect 110305 244961 110339 244989
rect 110367 244961 110401 244989
rect 110429 244961 110463 244989
rect 110491 244961 125637 244989
rect 125665 244961 125699 244989
rect 125727 244961 125761 244989
rect 125789 244961 125823 244989
rect 125851 244961 140997 244989
rect 141025 244961 141059 244989
rect 141087 244961 141121 244989
rect 141149 244961 141183 244989
rect 141211 244961 156357 244989
rect 156385 244961 156419 244989
rect 156447 244961 156481 244989
rect 156509 244961 156543 244989
rect 156571 244961 171717 244989
rect 171745 244961 171779 244989
rect 171807 244961 171841 244989
rect 171869 244961 171903 244989
rect 171931 244961 187077 244989
rect 187105 244961 187139 244989
rect 187167 244961 187201 244989
rect 187229 244961 187263 244989
rect 187291 244961 202437 244989
rect 202465 244961 202499 244989
rect 202527 244961 202561 244989
rect 202589 244961 202623 244989
rect 202651 244961 217797 244989
rect 217825 244961 217859 244989
rect 217887 244961 217921 244989
rect 217949 244961 217983 244989
rect 218011 244961 233157 244989
rect 233185 244961 233219 244989
rect 233247 244961 233281 244989
rect 233309 244961 233343 244989
rect 233371 244961 248517 244989
rect 248545 244961 248579 244989
rect 248607 244961 248641 244989
rect 248669 244961 248703 244989
rect 248731 244961 263877 244989
rect 263905 244961 263939 244989
rect 263967 244961 264001 244989
rect 264029 244961 264063 244989
rect 264091 244961 279237 244989
rect 279265 244961 279299 244989
rect 279327 244961 279361 244989
rect 279389 244961 279423 244989
rect 279451 244961 294597 244989
rect 294625 244961 294659 244989
rect 294687 244961 294721 244989
rect 294749 244961 294783 244989
rect 294811 244961 298248 244989
rect 298276 244961 298310 244989
rect 298338 244961 298372 244989
rect 298400 244961 298434 244989
rect 298462 244961 298990 244989
rect -958 244913 298990 244961
rect -958 239175 298990 239223
rect -958 239147 -910 239175
rect -882 239147 -848 239175
rect -820 239147 -786 239175
rect -758 239147 -724 239175
rect -696 239147 4617 239175
rect 4645 239147 4679 239175
rect 4707 239147 4741 239175
rect 4769 239147 4803 239175
rect 4831 239147 19977 239175
rect 20005 239147 20039 239175
rect 20067 239147 20101 239175
rect 20129 239147 20163 239175
rect 20191 239147 35337 239175
rect 35365 239147 35399 239175
rect 35427 239147 35461 239175
rect 35489 239147 35523 239175
rect 35551 239147 50697 239175
rect 50725 239147 50759 239175
rect 50787 239147 50821 239175
rect 50849 239147 50883 239175
rect 50911 239147 66057 239175
rect 66085 239147 66119 239175
rect 66147 239147 66181 239175
rect 66209 239147 66243 239175
rect 66271 239147 81417 239175
rect 81445 239147 81479 239175
rect 81507 239147 81541 239175
rect 81569 239147 81603 239175
rect 81631 239147 96777 239175
rect 96805 239147 96839 239175
rect 96867 239147 96901 239175
rect 96929 239147 96963 239175
rect 96991 239147 112137 239175
rect 112165 239147 112199 239175
rect 112227 239147 112261 239175
rect 112289 239147 112323 239175
rect 112351 239147 127497 239175
rect 127525 239147 127559 239175
rect 127587 239147 127621 239175
rect 127649 239147 127683 239175
rect 127711 239147 142857 239175
rect 142885 239147 142919 239175
rect 142947 239147 142981 239175
rect 143009 239147 143043 239175
rect 143071 239147 158217 239175
rect 158245 239147 158279 239175
rect 158307 239147 158341 239175
rect 158369 239147 158403 239175
rect 158431 239147 173577 239175
rect 173605 239147 173639 239175
rect 173667 239147 173701 239175
rect 173729 239147 173763 239175
rect 173791 239147 188937 239175
rect 188965 239147 188999 239175
rect 189027 239147 189061 239175
rect 189089 239147 189123 239175
rect 189151 239147 204297 239175
rect 204325 239147 204359 239175
rect 204387 239147 204421 239175
rect 204449 239147 204483 239175
rect 204511 239147 219657 239175
rect 219685 239147 219719 239175
rect 219747 239147 219781 239175
rect 219809 239147 219843 239175
rect 219871 239147 235017 239175
rect 235045 239147 235079 239175
rect 235107 239147 235141 239175
rect 235169 239147 235203 239175
rect 235231 239147 250377 239175
rect 250405 239147 250439 239175
rect 250467 239147 250501 239175
rect 250529 239147 250563 239175
rect 250591 239147 265737 239175
rect 265765 239147 265799 239175
rect 265827 239147 265861 239175
rect 265889 239147 265923 239175
rect 265951 239147 281097 239175
rect 281125 239147 281159 239175
rect 281187 239147 281221 239175
rect 281249 239147 281283 239175
rect 281311 239147 296457 239175
rect 296485 239147 296519 239175
rect 296547 239147 296581 239175
rect 296609 239147 296643 239175
rect 296671 239147 298728 239175
rect 298756 239147 298790 239175
rect 298818 239147 298852 239175
rect 298880 239147 298914 239175
rect 298942 239147 298990 239175
rect -958 239113 298990 239147
rect -958 239085 -910 239113
rect -882 239085 -848 239113
rect -820 239085 -786 239113
rect -758 239085 -724 239113
rect -696 239085 4617 239113
rect 4645 239085 4679 239113
rect 4707 239085 4741 239113
rect 4769 239085 4803 239113
rect 4831 239085 19977 239113
rect 20005 239085 20039 239113
rect 20067 239085 20101 239113
rect 20129 239085 20163 239113
rect 20191 239085 35337 239113
rect 35365 239085 35399 239113
rect 35427 239085 35461 239113
rect 35489 239085 35523 239113
rect 35551 239085 50697 239113
rect 50725 239085 50759 239113
rect 50787 239085 50821 239113
rect 50849 239085 50883 239113
rect 50911 239085 66057 239113
rect 66085 239085 66119 239113
rect 66147 239085 66181 239113
rect 66209 239085 66243 239113
rect 66271 239085 81417 239113
rect 81445 239085 81479 239113
rect 81507 239085 81541 239113
rect 81569 239085 81603 239113
rect 81631 239085 96777 239113
rect 96805 239085 96839 239113
rect 96867 239085 96901 239113
rect 96929 239085 96963 239113
rect 96991 239085 112137 239113
rect 112165 239085 112199 239113
rect 112227 239085 112261 239113
rect 112289 239085 112323 239113
rect 112351 239085 127497 239113
rect 127525 239085 127559 239113
rect 127587 239085 127621 239113
rect 127649 239085 127683 239113
rect 127711 239085 142857 239113
rect 142885 239085 142919 239113
rect 142947 239085 142981 239113
rect 143009 239085 143043 239113
rect 143071 239085 158217 239113
rect 158245 239085 158279 239113
rect 158307 239085 158341 239113
rect 158369 239085 158403 239113
rect 158431 239085 173577 239113
rect 173605 239085 173639 239113
rect 173667 239085 173701 239113
rect 173729 239085 173763 239113
rect 173791 239085 188937 239113
rect 188965 239085 188999 239113
rect 189027 239085 189061 239113
rect 189089 239085 189123 239113
rect 189151 239085 204297 239113
rect 204325 239085 204359 239113
rect 204387 239085 204421 239113
rect 204449 239085 204483 239113
rect 204511 239085 219657 239113
rect 219685 239085 219719 239113
rect 219747 239085 219781 239113
rect 219809 239085 219843 239113
rect 219871 239085 235017 239113
rect 235045 239085 235079 239113
rect 235107 239085 235141 239113
rect 235169 239085 235203 239113
rect 235231 239085 250377 239113
rect 250405 239085 250439 239113
rect 250467 239085 250501 239113
rect 250529 239085 250563 239113
rect 250591 239085 265737 239113
rect 265765 239085 265799 239113
rect 265827 239085 265861 239113
rect 265889 239085 265923 239113
rect 265951 239085 281097 239113
rect 281125 239085 281159 239113
rect 281187 239085 281221 239113
rect 281249 239085 281283 239113
rect 281311 239085 296457 239113
rect 296485 239085 296519 239113
rect 296547 239085 296581 239113
rect 296609 239085 296643 239113
rect 296671 239085 298728 239113
rect 298756 239085 298790 239113
rect 298818 239085 298852 239113
rect 298880 239085 298914 239113
rect 298942 239085 298990 239113
rect -958 239051 298990 239085
rect -958 239023 -910 239051
rect -882 239023 -848 239051
rect -820 239023 -786 239051
rect -758 239023 -724 239051
rect -696 239023 4617 239051
rect 4645 239023 4679 239051
rect 4707 239023 4741 239051
rect 4769 239023 4803 239051
rect 4831 239023 19977 239051
rect 20005 239023 20039 239051
rect 20067 239023 20101 239051
rect 20129 239023 20163 239051
rect 20191 239023 35337 239051
rect 35365 239023 35399 239051
rect 35427 239023 35461 239051
rect 35489 239023 35523 239051
rect 35551 239023 50697 239051
rect 50725 239023 50759 239051
rect 50787 239023 50821 239051
rect 50849 239023 50883 239051
rect 50911 239023 66057 239051
rect 66085 239023 66119 239051
rect 66147 239023 66181 239051
rect 66209 239023 66243 239051
rect 66271 239023 81417 239051
rect 81445 239023 81479 239051
rect 81507 239023 81541 239051
rect 81569 239023 81603 239051
rect 81631 239023 96777 239051
rect 96805 239023 96839 239051
rect 96867 239023 96901 239051
rect 96929 239023 96963 239051
rect 96991 239023 112137 239051
rect 112165 239023 112199 239051
rect 112227 239023 112261 239051
rect 112289 239023 112323 239051
rect 112351 239023 127497 239051
rect 127525 239023 127559 239051
rect 127587 239023 127621 239051
rect 127649 239023 127683 239051
rect 127711 239023 142857 239051
rect 142885 239023 142919 239051
rect 142947 239023 142981 239051
rect 143009 239023 143043 239051
rect 143071 239023 158217 239051
rect 158245 239023 158279 239051
rect 158307 239023 158341 239051
rect 158369 239023 158403 239051
rect 158431 239023 173577 239051
rect 173605 239023 173639 239051
rect 173667 239023 173701 239051
rect 173729 239023 173763 239051
rect 173791 239023 188937 239051
rect 188965 239023 188999 239051
rect 189027 239023 189061 239051
rect 189089 239023 189123 239051
rect 189151 239023 204297 239051
rect 204325 239023 204359 239051
rect 204387 239023 204421 239051
rect 204449 239023 204483 239051
rect 204511 239023 219657 239051
rect 219685 239023 219719 239051
rect 219747 239023 219781 239051
rect 219809 239023 219843 239051
rect 219871 239023 235017 239051
rect 235045 239023 235079 239051
rect 235107 239023 235141 239051
rect 235169 239023 235203 239051
rect 235231 239023 250377 239051
rect 250405 239023 250439 239051
rect 250467 239023 250501 239051
rect 250529 239023 250563 239051
rect 250591 239023 265737 239051
rect 265765 239023 265799 239051
rect 265827 239023 265861 239051
rect 265889 239023 265923 239051
rect 265951 239023 281097 239051
rect 281125 239023 281159 239051
rect 281187 239023 281221 239051
rect 281249 239023 281283 239051
rect 281311 239023 296457 239051
rect 296485 239023 296519 239051
rect 296547 239023 296581 239051
rect 296609 239023 296643 239051
rect 296671 239023 298728 239051
rect 298756 239023 298790 239051
rect 298818 239023 298852 239051
rect 298880 239023 298914 239051
rect 298942 239023 298990 239051
rect -958 238989 298990 239023
rect -958 238961 -910 238989
rect -882 238961 -848 238989
rect -820 238961 -786 238989
rect -758 238961 -724 238989
rect -696 238961 4617 238989
rect 4645 238961 4679 238989
rect 4707 238961 4741 238989
rect 4769 238961 4803 238989
rect 4831 238961 19977 238989
rect 20005 238961 20039 238989
rect 20067 238961 20101 238989
rect 20129 238961 20163 238989
rect 20191 238961 35337 238989
rect 35365 238961 35399 238989
rect 35427 238961 35461 238989
rect 35489 238961 35523 238989
rect 35551 238961 50697 238989
rect 50725 238961 50759 238989
rect 50787 238961 50821 238989
rect 50849 238961 50883 238989
rect 50911 238961 66057 238989
rect 66085 238961 66119 238989
rect 66147 238961 66181 238989
rect 66209 238961 66243 238989
rect 66271 238961 81417 238989
rect 81445 238961 81479 238989
rect 81507 238961 81541 238989
rect 81569 238961 81603 238989
rect 81631 238961 96777 238989
rect 96805 238961 96839 238989
rect 96867 238961 96901 238989
rect 96929 238961 96963 238989
rect 96991 238961 112137 238989
rect 112165 238961 112199 238989
rect 112227 238961 112261 238989
rect 112289 238961 112323 238989
rect 112351 238961 127497 238989
rect 127525 238961 127559 238989
rect 127587 238961 127621 238989
rect 127649 238961 127683 238989
rect 127711 238961 142857 238989
rect 142885 238961 142919 238989
rect 142947 238961 142981 238989
rect 143009 238961 143043 238989
rect 143071 238961 158217 238989
rect 158245 238961 158279 238989
rect 158307 238961 158341 238989
rect 158369 238961 158403 238989
rect 158431 238961 173577 238989
rect 173605 238961 173639 238989
rect 173667 238961 173701 238989
rect 173729 238961 173763 238989
rect 173791 238961 188937 238989
rect 188965 238961 188999 238989
rect 189027 238961 189061 238989
rect 189089 238961 189123 238989
rect 189151 238961 204297 238989
rect 204325 238961 204359 238989
rect 204387 238961 204421 238989
rect 204449 238961 204483 238989
rect 204511 238961 219657 238989
rect 219685 238961 219719 238989
rect 219747 238961 219781 238989
rect 219809 238961 219843 238989
rect 219871 238961 235017 238989
rect 235045 238961 235079 238989
rect 235107 238961 235141 238989
rect 235169 238961 235203 238989
rect 235231 238961 250377 238989
rect 250405 238961 250439 238989
rect 250467 238961 250501 238989
rect 250529 238961 250563 238989
rect 250591 238961 265737 238989
rect 265765 238961 265799 238989
rect 265827 238961 265861 238989
rect 265889 238961 265923 238989
rect 265951 238961 281097 238989
rect 281125 238961 281159 238989
rect 281187 238961 281221 238989
rect 281249 238961 281283 238989
rect 281311 238961 296457 238989
rect 296485 238961 296519 238989
rect 296547 238961 296581 238989
rect 296609 238961 296643 238989
rect 296671 238961 298728 238989
rect 298756 238961 298790 238989
rect 298818 238961 298852 238989
rect 298880 238961 298914 238989
rect 298942 238961 298990 238989
rect -958 238913 298990 238961
rect -958 236175 298990 236223
rect -958 236147 -430 236175
rect -402 236147 -368 236175
rect -340 236147 -306 236175
rect -278 236147 -244 236175
rect -216 236147 2757 236175
rect 2785 236147 2819 236175
rect 2847 236147 2881 236175
rect 2909 236147 2943 236175
rect 2971 236147 18117 236175
rect 18145 236147 18179 236175
rect 18207 236147 18241 236175
rect 18269 236147 18303 236175
rect 18331 236147 33477 236175
rect 33505 236147 33539 236175
rect 33567 236147 33601 236175
rect 33629 236147 33663 236175
rect 33691 236147 48837 236175
rect 48865 236147 48899 236175
rect 48927 236147 48961 236175
rect 48989 236147 49023 236175
rect 49051 236147 64197 236175
rect 64225 236147 64259 236175
rect 64287 236147 64321 236175
rect 64349 236147 64383 236175
rect 64411 236147 79557 236175
rect 79585 236147 79619 236175
rect 79647 236147 79681 236175
rect 79709 236147 79743 236175
rect 79771 236147 94917 236175
rect 94945 236147 94979 236175
rect 95007 236147 95041 236175
rect 95069 236147 95103 236175
rect 95131 236147 110277 236175
rect 110305 236147 110339 236175
rect 110367 236147 110401 236175
rect 110429 236147 110463 236175
rect 110491 236147 125637 236175
rect 125665 236147 125699 236175
rect 125727 236147 125761 236175
rect 125789 236147 125823 236175
rect 125851 236147 140997 236175
rect 141025 236147 141059 236175
rect 141087 236147 141121 236175
rect 141149 236147 141183 236175
rect 141211 236147 156357 236175
rect 156385 236147 156419 236175
rect 156447 236147 156481 236175
rect 156509 236147 156543 236175
rect 156571 236147 171717 236175
rect 171745 236147 171779 236175
rect 171807 236147 171841 236175
rect 171869 236147 171903 236175
rect 171931 236147 187077 236175
rect 187105 236147 187139 236175
rect 187167 236147 187201 236175
rect 187229 236147 187263 236175
rect 187291 236147 202437 236175
rect 202465 236147 202499 236175
rect 202527 236147 202561 236175
rect 202589 236147 202623 236175
rect 202651 236147 217797 236175
rect 217825 236147 217859 236175
rect 217887 236147 217921 236175
rect 217949 236147 217983 236175
rect 218011 236147 233157 236175
rect 233185 236147 233219 236175
rect 233247 236147 233281 236175
rect 233309 236147 233343 236175
rect 233371 236147 248517 236175
rect 248545 236147 248579 236175
rect 248607 236147 248641 236175
rect 248669 236147 248703 236175
rect 248731 236147 263877 236175
rect 263905 236147 263939 236175
rect 263967 236147 264001 236175
rect 264029 236147 264063 236175
rect 264091 236147 279237 236175
rect 279265 236147 279299 236175
rect 279327 236147 279361 236175
rect 279389 236147 279423 236175
rect 279451 236147 294597 236175
rect 294625 236147 294659 236175
rect 294687 236147 294721 236175
rect 294749 236147 294783 236175
rect 294811 236147 298248 236175
rect 298276 236147 298310 236175
rect 298338 236147 298372 236175
rect 298400 236147 298434 236175
rect 298462 236147 298990 236175
rect -958 236113 298990 236147
rect -958 236085 -430 236113
rect -402 236085 -368 236113
rect -340 236085 -306 236113
rect -278 236085 -244 236113
rect -216 236085 2757 236113
rect 2785 236085 2819 236113
rect 2847 236085 2881 236113
rect 2909 236085 2943 236113
rect 2971 236085 18117 236113
rect 18145 236085 18179 236113
rect 18207 236085 18241 236113
rect 18269 236085 18303 236113
rect 18331 236085 33477 236113
rect 33505 236085 33539 236113
rect 33567 236085 33601 236113
rect 33629 236085 33663 236113
rect 33691 236085 48837 236113
rect 48865 236085 48899 236113
rect 48927 236085 48961 236113
rect 48989 236085 49023 236113
rect 49051 236085 64197 236113
rect 64225 236085 64259 236113
rect 64287 236085 64321 236113
rect 64349 236085 64383 236113
rect 64411 236085 79557 236113
rect 79585 236085 79619 236113
rect 79647 236085 79681 236113
rect 79709 236085 79743 236113
rect 79771 236085 94917 236113
rect 94945 236085 94979 236113
rect 95007 236085 95041 236113
rect 95069 236085 95103 236113
rect 95131 236085 110277 236113
rect 110305 236085 110339 236113
rect 110367 236085 110401 236113
rect 110429 236085 110463 236113
rect 110491 236085 125637 236113
rect 125665 236085 125699 236113
rect 125727 236085 125761 236113
rect 125789 236085 125823 236113
rect 125851 236085 140997 236113
rect 141025 236085 141059 236113
rect 141087 236085 141121 236113
rect 141149 236085 141183 236113
rect 141211 236085 156357 236113
rect 156385 236085 156419 236113
rect 156447 236085 156481 236113
rect 156509 236085 156543 236113
rect 156571 236085 171717 236113
rect 171745 236085 171779 236113
rect 171807 236085 171841 236113
rect 171869 236085 171903 236113
rect 171931 236085 187077 236113
rect 187105 236085 187139 236113
rect 187167 236085 187201 236113
rect 187229 236085 187263 236113
rect 187291 236085 202437 236113
rect 202465 236085 202499 236113
rect 202527 236085 202561 236113
rect 202589 236085 202623 236113
rect 202651 236085 217797 236113
rect 217825 236085 217859 236113
rect 217887 236085 217921 236113
rect 217949 236085 217983 236113
rect 218011 236085 233157 236113
rect 233185 236085 233219 236113
rect 233247 236085 233281 236113
rect 233309 236085 233343 236113
rect 233371 236085 248517 236113
rect 248545 236085 248579 236113
rect 248607 236085 248641 236113
rect 248669 236085 248703 236113
rect 248731 236085 263877 236113
rect 263905 236085 263939 236113
rect 263967 236085 264001 236113
rect 264029 236085 264063 236113
rect 264091 236085 279237 236113
rect 279265 236085 279299 236113
rect 279327 236085 279361 236113
rect 279389 236085 279423 236113
rect 279451 236085 294597 236113
rect 294625 236085 294659 236113
rect 294687 236085 294721 236113
rect 294749 236085 294783 236113
rect 294811 236085 298248 236113
rect 298276 236085 298310 236113
rect 298338 236085 298372 236113
rect 298400 236085 298434 236113
rect 298462 236085 298990 236113
rect -958 236051 298990 236085
rect -958 236023 -430 236051
rect -402 236023 -368 236051
rect -340 236023 -306 236051
rect -278 236023 -244 236051
rect -216 236023 2757 236051
rect 2785 236023 2819 236051
rect 2847 236023 2881 236051
rect 2909 236023 2943 236051
rect 2971 236023 18117 236051
rect 18145 236023 18179 236051
rect 18207 236023 18241 236051
rect 18269 236023 18303 236051
rect 18331 236023 33477 236051
rect 33505 236023 33539 236051
rect 33567 236023 33601 236051
rect 33629 236023 33663 236051
rect 33691 236023 48837 236051
rect 48865 236023 48899 236051
rect 48927 236023 48961 236051
rect 48989 236023 49023 236051
rect 49051 236023 64197 236051
rect 64225 236023 64259 236051
rect 64287 236023 64321 236051
rect 64349 236023 64383 236051
rect 64411 236023 79557 236051
rect 79585 236023 79619 236051
rect 79647 236023 79681 236051
rect 79709 236023 79743 236051
rect 79771 236023 94917 236051
rect 94945 236023 94979 236051
rect 95007 236023 95041 236051
rect 95069 236023 95103 236051
rect 95131 236023 110277 236051
rect 110305 236023 110339 236051
rect 110367 236023 110401 236051
rect 110429 236023 110463 236051
rect 110491 236023 125637 236051
rect 125665 236023 125699 236051
rect 125727 236023 125761 236051
rect 125789 236023 125823 236051
rect 125851 236023 140997 236051
rect 141025 236023 141059 236051
rect 141087 236023 141121 236051
rect 141149 236023 141183 236051
rect 141211 236023 156357 236051
rect 156385 236023 156419 236051
rect 156447 236023 156481 236051
rect 156509 236023 156543 236051
rect 156571 236023 171717 236051
rect 171745 236023 171779 236051
rect 171807 236023 171841 236051
rect 171869 236023 171903 236051
rect 171931 236023 187077 236051
rect 187105 236023 187139 236051
rect 187167 236023 187201 236051
rect 187229 236023 187263 236051
rect 187291 236023 202437 236051
rect 202465 236023 202499 236051
rect 202527 236023 202561 236051
rect 202589 236023 202623 236051
rect 202651 236023 217797 236051
rect 217825 236023 217859 236051
rect 217887 236023 217921 236051
rect 217949 236023 217983 236051
rect 218011 236023 233157 236051
rect 233185 236023 233219 236051
rect 233247 236023 233281 236051
rect 233309 236023 233343 236051
rect 233371 236023 248517 236051
rect 248545 236023 248579 236051
rect 248607 236023 248641 236051
rect 248669 236023 248703 236051
rect 248731 236023 263877 236051
rect 263905 236023 263939 236051
rect 263967 236023 264001 236051
rect 264029 236023 264063 236051
rect 264091 236023 279237 236051
rect 279265 236023 279299 236051
rect 279327 236023 279361 236051
rect 279389 236023 279423 236051
rect 279451 236023 294597 236051
rect 294625 236023 294659 236051
rect 294687 236023 294721 236051
rect 294749 236023 294783 236051
rect 294811 236023 298248 236051
rect 298276 236023 298310 236051
rect 298338 236023 298372 236051
rect 298400 236023 298434 236051
rect 298462 236023 298990 236051
rect -958 235989 298990 236023
rect -958 235961 -430 235989
rect -402 235961 -368 235989
rect -340 235961 -306 235989
rect -278 235961 -244 235989
rect -216 235961 2757 235989
rect 2785 235961 2819 235989
rect 2847 235961 2881 235989
rect 2909 235961 2943 235989
rect 2971 235961 18117 235989
rect 18145 235961 18179 235989
rect 18207 235961 18241 235989
rect 18269 235961 18303 235989
rect 18331 235961 33477 235989
rect 33505 235961 33539 235989
rect 33567 235961 33601 235989
rect 33629 235961 33663 235989
rect 33691 235961 48837 235989
rect 48865 235961 48899 235989
rect 48927 235961 48961 235989
rect 48989 235961 49023 235989
rect 49051 235961 64197 235989
rect 64225 235961 64259 235989
rect 64287 235961 64321 235989
rect 64349 235961 64383 235989
rect 64411 235961 79557 235989
rect 79585 235961 79619 235989
rect 79647 235961 79681 235989
rect 79709 235961 79743 235989
rect 79771 235961 94917 235989
rect 94945 235961 94979 235989
rect 95007 235961 95041 235989
rect 95069 235961 95103 235989
rect 95131 235961 110277 235989
rect 110305 235961 110339 235989
rect 110367 235961 110401 235989
rect 110429 235961 110463 235989
rect 110491 235961 125637 235989
rect 125665 235961 125699 235989
rect 125727 235961 125761 235989
rect 125789 235961 125823 235989
rect 125851 235961 140997 235989
rect 141025 235961 141059 235989
rect 141087 235961 141121 235989
rect 141149 235961 141183 235989
rect 141211 235961 156357 235989
rect 156385 235961 156419 235989
rect 156447 235961 156481 235989
rect 156509 235961 156543 235989
rect 156571 235961 171717 235989
rect 171745 235961 171779 235989
rect 171807 235961 171841 235989
rect 171869 235961 171903 235989
rect 171931 235961 187077 235989
rect 187105 235961 187139 235989
rect 187167 235961 187201 235989
rect 187229 235961 187263 235989
rect 187291 235961 202437 235989
rect 202465 235961 202499 235989
rect 202527 235961 202561 235989
rect 202589 235961 202623 235989
rect 202651 235961 217797 235989
rect 217825 235961 217859 235989
rect 217887 235961 217921 235989
rect 217949 235961 217983 235989
rect 218011 235961 233157 235989
rect 233185 235961 233219 235989
rect 233247 235961 233281 235989
rect 233309 235961 233343 235989
rect 233371 235961 248517 235989
rect 248545 235961 248579 235989
rect 248607 235961 248641 235989
rect 248669 235961 248703 235989
rect 248731 235961 263877 235989
rect 263905 235961 263939 235989
rect 263967 235961 264001 235989
rect 264029 235961 264063 235989
rect 264091 235961 279237 235989
rect 279265 235961 279299 235989
rect 279327 235961 279361 235989
rect 279389 235961 279423 235989
rect 279451 235961 294597 235989
rect 294625 235961 294659 235989
rect 294687 235961 294721 235989
rect 294749 235961 294783 235989
rect 294811 235961 298248 235989
rect 298276 235961 298310 235989
rect 298338 235961 298372 235989
rect 298400 235961 298434 235989
rect 298462 235961 298990 235989
rect -958 235913 298990 235961
rect -958 230175 298990 230223
rect -958 230147 -910 230175
rect -882 230147 -848 230175
rect -820 230147 -786 230175
rect -758 230147 -724 230175
rect -696 230147 4617 230175
rect 4645 230147 4679 230175
rect 4707 230147 4741 230175
rect 4769 230147 4803 230175
rect 4831 230147 19977 230175
rect 20005 230147 20039 230175
rect 20067 230147 20101 230175
rect 20129 230147 20163 230175
rect 20191 230147 35337 230175
rect 35365 230147 35399 230175
rect 35427 230147 35461 230175
rect 35489 230147 35523 230175
rect 35551 230147 50697 230175
rect 50725 230147 50759 230175
rect 50787 230147 50821 230175
rect 50849 230147 50883 230175
rect 50911 230147 66057 230175
rect 66085 230147 66119 230175
rect 66147 230147 66181 230175
rect 66209 230147 66243 230175
rect 66271 230147 81417 230175
rect 81445 230147 81479 230175
rect 81507 230147 81541 230175
rect 81569 230147 81603 230175
rect 81631 230147 96777 230175
rect 96805 230147 96839 230175
rect 96867 230147 96901 230175
rect 96929 230147 96963 230175
rect 96991 230147 112137 230175
rect 112165 230147 112199 230175
rect 112227 230147 112261 230175
rect 112289 230147 112323 230175
rect 112351 230147 127497 230175
rect 127525 230147 127559 230175
rect 127587 230147 127621 230175
rect 127649 230147 127683 230175
rect 127711 230147 142857 230175
rect 142885 230147 142919 230175
rect 142947 230147 142981 230175
rect 143009 230147 143043 230175
rect 143071 230147 158217 230175
rect 158245 230147 158279 230175
rect 158307 230147 158341 230175
rect 158369 230147 158403 230175
rect 158431 230147 173577 230175
rect 173605 230147 173639 230175
rect 173667 230147 173701 230175
rect 173729 230147 173763 230175
rect 173791 230147 188937 230175
rect 188965 230147 188999 230175
rect 189027 230147 189061 230175
rect 189089 230147 189123 230175
rect 189151 230147 204297 230175
rect 204325 230147 204359 230175
rect 204387 230147 204421 230175
rect 204449 230147 204483 230175
rect 204511 230147 219657 230175
rect 219685 230147 219719 230175
rect 219747 230147 219781 230175
rect 219809 230147 219843 230175
rect 219871 230147 235017 230175
rect 235045 230147 235079 230175
rect 235107 230147 235141 230175
rect 235169 230147 235203 230175
rect 235231 230147 250377 230175
rect 250405 230147 250439 230175
rect 250467 230147 250501 230175
rect 250529 230147 250563 230175
rect 250591 230147 265737 230175
rect 265765 230147 265799 230175
rect 265827 230147 265861 230175
rect 265889 230147 265923 230175
rect 265951 230147 281097 230175
rect 281125 230147 281159 230175
rect 281187 230147 281221 230175
rect 281249 230147 281283 230175
rect 281311 230147 296457 230175
rect 296485 230147 296519 230175
rect 296547 230147 296581 230175
rect 296609 230147 296643 230175
rect 296671 230147 298728 230175
rect 298756 230147 298790 230175
rect 298818 230147 298852 230175
rect 298880 230147 298914 230175
rect 298942 230147 298990 230175
rect -958 230113 298990 230147
rect -958 230085 -910 230113
rect -882 230085 -848 230113
rect -820 230085 -786 230113
rect -758 230085 -724 230113
rect -696 230085 4617 230113
rect 4645 230085 4679 230113
rect 4707 230085 4741 230113
rect 4769 230085 4803 230113
rect 4831 230085 19977 230113
rect 20005 230085 20039 230113
rect 20067 230085 20101 230113
rect 20129 230085 20163 230113
rect 20191 230085 35337 230113
rect 35365 230085 35399 230113
rect 35427 230085 35461 230113
rect 35489 230085 35523 230113
rect 35551 230085 50697 230113
rect 50725 230085 50759 230113
rect 50787 230085 50821 230113
rect 50849 230085 50883 230113
rect 50911 230085 66057 230113
rect 66085 230085 66119 230113
rect 66147 230085 66181 230113
rect 66209 230085 66243 230113
rect 66271 230085 81417 230113
rect 81445 230085 81479 230113
rect 81507 230085 81541 230113
rect 81569 230085 81603 230113
rect 81631 230085 96777 230113
rect 96805 230085 96839 230113
rect 96867 230085 96901 230113
rect 96929 230085 96963 230113
rect 96991 230085 112137 230113
rect 112165 230085 112199 230113
rect 112227 230085 112261 230113
rect 112289 230085 112323 230113
rect 112351 230085 127497 230113
rect 127525 230085 127559 230113
rect 127587 230085 127621 230113
rect 127649 230085 127683 230113
rect 127711 230085 142857 230113
rect 142885 230085 142919 230113
rect 142947 230085 142981 230113
rect 143009 230085 143043 230113
rect 143071 230085 158217 230113
rect 158245 230085 158279 230113
rect 158307 230085 158341 230113
rect 158369 230085 158403 230113
rect 158431 230085 173577 230113
rect 173605 230085 173639 230113
rect 173667 230085 173701 230113
rect 173729 230085 173763 230113
rect 173791 230085 188937 230113
rect 188965 230085 188999 230113
rect 189027 230085 189061 230113
rect 189089 230085 189123 230113
rect 189151 230085 204297 230113
rect 204325 230085 204359 230113
rect 204387 230085 204421 230113
rect 204449 230085 204483 230113
rect 204511 230085 219657 230113
rect 219685 230085 219719 230113
rect 219747 230085 219781 230113
rect 219809 230085 219843 230113
rect 219871 230085 235017 230113
rect 235045 230085 235079 230113
rect 235107 230085 235141 230113
rect 235169 230085 235203 230113
rect 235231 230085 250377 230113
rect 250405 230085 250439 230113
rect 250467 230085 250501 230113
rect 250529 230085 250563 230113
rect 250591 230085 265737 230113
rect 265765 230085 265799 230113
rect 265827 230085 265861 230113
rect 265889 230085 265923 230113
rect 265951 230085 281097 230113
rect 281125 230085 281159 230113
rect 281187 230085 281221 230113
rect 281249 230085 281283 230113
rect 281311 230085 296457 230113
rect 296485 230085 296519 230113
rect 296547 230085 296581 230113
rect 296609 230085 296643 230113
rect 296671 230085 298728 230113
rect 298756 230085 298790 230113
rect 298818 230085 298852 230113
rect 298880 230085 298914 230113
rect 298942 230085 298990 230113
rect -958 230051 298990 230085
rect -958 230023 -910 230051
rect -882 230023 -848 230051
rect -820 230023 -786 230051
rect -758 230023 -724 230051
rect -696 230023 4617 230051
rect 4645 230023 4679 230051
rect 4707 230023 4741 230051
rect 4769 230023 4803 230051
rect 4831 230023 19977 230051
rect 20005 230023 20039 230051
rect 20067 230023 20101 230051
rect 20129 230023 20163 230051
rect 20191 230023 35337 230051
rect 35365 230023 35399 230051
rect 35427 230023 35461 230051
rect 35489 230023 35523 230051
rect 35551 230023 50697 230051
rect 50725 230023 50759 230051
rect 50787 230023 50821 230051
rect 50849 230023 50883 230051
rect 50911 230023 66057 230051
rect 66085 230023 66119 230051
rect 66147 230023 66181 230051
rect 66209 230023 66243 230051
rect 66271 230023 81417 230051
rect 81445 230023 81479 230051
rect 81507 230023 81541 230051
rect 81569 230023 81603 230051
rect 81631 230023 96777 230051
rect 96805 230023 96839 230051
rect 96867 230023 96901 230051
rect 96929 230023 96963 230051
rect 96991 230023 112137 230051
rect 112165 230023 112199 230051
rect 112227 230023 112261 230051
rect 112289 230023 112323 230051
rect 112351 230023 127497 230051
rect 127525 230023 127559 230051
rect 127587 230023 127621 230051
rect 127649 230023 127683 230051
rect 127711 230023 142857 230051
rect 142885 230023 142919 230051
rect 142947 230023 142981 230051
rect 143009 230023 143043 230051
rect 143071 230023 158217 230051
rect 158245 230023 158279 230051
rect 158307 230023 158341 230051
rect 158369 230023 158403 230051
rect 158431 230023 173577 230051
rect 173605 230023 173639 230051
rect 173667 230023 173701 230051
rect 173729 230023 173763 230051
rect 173791 230023 188937 230051
rect 188965 230023 188999 230051
rect 189027 230023 189061 230051
rect 189089 230023 189123 230051
rect 189151 230023 204297 230051
rect 204325 230023 204359 230051
rect 204387 230023 204421 230051
rect 204449 230023 204483 230051
rect 204511 230023 219657 230051
rect 219685 230023 219719 230051
rect 219747 230023 219781 230051
rect 219809 230023 219843 230051
rect 219871 230023 235017 230051
rect 235045 230023 235079 230051
rect 235107 230023 235141 230051
rect 235169 230023 235203 230051
rect 235231 230023 250377 230051
rect 250405 230023 250439 230051
rect 250467 230023 250501 230051
rect 250529 230023 250563 230051
rect 250591 230023 265737 230051
rect 265765 230023 265799 230051
rect 265827 230023 265861 230051
rect 265889 230023 265923 230051
rect 265951 230023 281097 230051
rect 281125 230023 281159 230051
rect 281187 230023 281221 230051
rect 281249 230023 281283 230051
rect 281311 230023 296457 230051
rect 296485 230023 296519 230051
rect 296547 230023 296581 230051
rect 296609 230023 296643 230051
rect 296671 230023 298728 230051
rect 298756 230023 298790 230051
rect 298818 230023 298852 230051
rect 298880 230023 298914 230051
rect 298942 230023 298990 230051
rect -958 229989 298990 230023
rect -958 229961 -910 229989
rect -882 229961 -848 229989
rect -820 229961 -786 229989
rect -758 229961 -724 229989
rect -696 229961 4617 229989
rect 4645 229961 4679 229989
rect 4707 229961 4741 229989
rect 4769 229961 4803 229989
rect 4831 229961 19977 229989
rect 20005 229961 20039 229989
rect 20067 229961 20101 229989
rect 20129 229961 20163 229989
rect 20191 229961 35337 229989
rect 35365 229961 35399 229989
rect 35427 229961 35461 229989
rect 35489 229961 35523 229989
rect 35551 229961 50697 229989
rect 50725 229961 50759 229989
rect 50787 229961 50821 229989
rect 50849 229961 50883 229989
rect 50911 229961 66057 229989
rect 66085 229961 66119 229989
rect 66147 229961 66181 229989
rect 66209 229961 66243 229989
rect 66271 229961 81417 229989
rect 81445 229961 81479 229989
rect 81507 229961 81541 229989
rect 81569 229961 81603 229989
rect 81631 229961 96777 229989
rect 96805 229961 96839 229989
rect 96867 229961 96901 229989
rect 96929 229961 96963 229989
rect 96991 229961 112137 229989
rect 112165 229961 112199 229989
rect 112227 229961 112261 229989
rect 112289 229961 112323 229989
rect 112351 229961 127497 229989
rect 127525 229961 127559 229989
rect 127587 229961 127621 229989
rect 127649 229961 127683 229989
rect 127711 229961 142857 229989
rect 142885 229961 142919 229989
rect 142947 229961 142981 229989
rect 143009 229961 143043 229989
rect 143071 229961 158217 229989
rect 158245 229961 158279 229989
rect 158307 229961 158341 229989
rect 158369 229961 158403 229989
rect 158431 229961 173577 229989
rect 173605 229961 173639 229989
rect 173667 229961 173701 229989
rect 173729 229961 173763 229989
rect 173791 229961 188937 229989
rect 188965 229961 188999 229989
rect 189027 229961 189061 229989
rect 189089 229961 189123 229989
rect 189151 229961 204297 229989
rect 204325 229961 204359 229989
rect 204387 229961 204421 229989
rect 204449 229961 204483 229989
rect 204511 229961 219657 229989
rect 219685 229961 219719 229989
rect 219747 229961 219781 229989
rect 219809 229961 219843 229989
rect 219871 229961 235017 229989
rect 235045 229961 235079 229989
rect 235107 229961 235141 229989
rect 235169 229961 235203 229989
rect 235231 229961 250377 229989
rect 250405 229961 250439 229989
rect 250467 229961 250501 229989
rect 250529 229961 250563 229989
rect 250591 229961 265737 229989
rect 265765 229961 265799 229989
rect 265827 229961 265861 229989
rect 265889 229961 265923 229989
rect 265951 229961 281097 229989
rect 281125 229961 281159 229989
rect 281187 229961 281221 229989
rect 281249 229961 281283 229989
rect 281311 229961 296457 229989
rect 296485 229961 296519 229989
rect 296547 229961 296581 229989
rect 296609 229961 296643 229989
rect 296671 229961 298728 229989
rect 298756 229961 298790 229989
rect 298818 229961 298852 229989
rect 298880 229961 298914 229989
rect 298942 229961 298990 229989
rect -958 229913 298990 229961
rect -958 227175 298990 227223
rect -958 227147 -430 227175
rect -402 227147 -368 227175
rect -340 227147 -306 227175
rect -278 227147 -244 227175
rect -216 227147 2757 227175
rect 2785 227147 2819 227175
rect 2847 227147 2881 227175
rect 2909 227147 2943 227175
rect 2971 227147 18117 227175
rect 18145 227147 18179 227175
rect 18207 227147 18241 227175
rect 18269 227147 18303 227175
rect 18331 227147 33477 227175
rect 33505 227147 33539 227175
rect 33567 227147 33601 227175
rect 33629 227147 33663 227175
rect 33691 227147 48837 227175
rect 48865 227147 48899 227175
rect 48927 227147 48961 227175
rect 48989 227147 49023 227175
rect 49051 227147 64197 227175
rect 64225 227147 64259 227175
rect 64287 227147 64321 227175
rect 64349 227147 64383 227175
rect 64411 227147 79557 227175
rect 79585 227147 79619 227175
rect 79647 227147 79681 227175
rect 79709 227147 79743 227175
rect 79771 227147 94917 227175
rect 94945 227147 94979 227175
rect 95007 227147 95041 227175
rect 95069 227147 95103 227175
rect 95131 227147 110277 227175
rect 110305 227147 110339 227175
rect 110367 227147 110401 227175
rect 110429 227147 110463 227175
rect 110491 227147 125637 227175
rect 125665 227147 125699 227175
rect 125727 227147 125761 227175
rect 125789 227147 125823 227175
rect 125851 227147 140997 227175
rect 141025 227147 141059 227175
rect 141087 227147 141121 227175
rect 141149 227147 141183 227175
rect 141211 227147 156357 227175
rect 156385 227147 156419 227175
rect 156447 227147 156481 227175
rect 156509 227147 156543 227175
rect 156571 227147 171717 227175
rect 171745 227147 171779 227175
rect 171807 227147 171841 227175
rect 171869 227147 171903 227175
rect 171931 227147 187077 227175
rect 187105 227147 187139 227175
rect 187167 227147 187201 227175
rect 187229 227147 187263 227175
rect 187291 227147 202437 227175
rect 202465 227147 202499 227175
rect 202527 227147 202561 227175
rect 202589 227147 202623 227175
rect 202651 227147 217797 227175
rect 217825 227147 217859 227175
rect 217887 227147 217921 227175
rect 217949 227147 217983 227175
rect 218011 227147 233157 227175
rect 233185 227147 233219 227175
rect 233247 227147 233281 227175
rect 233309 227147 233343 227175
rect 233371 227147 248517 227175
rect 248545 227147 248579 227175
rect 248607 227147 248641 227175
rect 248669 227147 248703 227175
rect 248731 227147 263877 227175
rect 263905 227147 263939 227175
rect 263967 227147 264001 227175
rect 264029 227147 264063 227175
rect 264091 227147 279237 227175
rect 279265 227147 279299 227175
rect 279327 227147 279361 227175
rect 279389 227147 279423 227175
rect 279451 227147 294597 227175
rect 294625 227147 294659 227175
rect 294687 227147 294721 227175
rect 294749 227147 294783 227175
rect 294811 227147 298248 227175
rect 298276 227147 298310 227175
rect 298338 227147 298372 227175
rect 298400 227147 298434 227175
rect 298462 227147 298990 227175
rect -958 227113 298990 227147
rect -958 227085 -430 227113
rect -402 227085 -368 227113
rect -340 227085 -306 227113
rect -278 227085 -244 227113
rect -216 227085 2757 227113
rect 2785 227085 2819 227113
rect 2847 227085 2881 227113
rect 2909 227085 2943 227113
rect 2971 227085 18117 227113
rect 18145 227085 18179 227113
rect 18207 227085 18241 227113
rect 18269 227085 18303 227113
rect 18331 227085 33477 227113
rect 33505 227085 33539 227113
rect 33567 227085 33601 227113
rect 33629 227085 33663 227113
rect 33691 227085 48837 227113
rect 48865 227085 48899 227113
rect 48927 227085 48961 227113
rect 48989 227085 49023 227113
rect 49051 227085 64197 227113
rect 64225 227085 64259 227113
rect 64287 227085 64321 227113
rect 64349 227085 64383 227113
rect 64411 227085 79557 227113
rect 79585 227085 79619 227113
rect 79647 227085 79681 227113
rect 79709 227085 79743 227113
rect 79771 227085 94917 227113
rect 94945 227085 94979 227113
rect 95007 227085 95041 227113
rect 95069 227085 95103 227113
rect 95131 227085 110277 227113
rect 110305 227085 110339 227113
rect 110367 227085 110401 227113
rect 110429 227085 110463 227113
rect 110491 227085 125637 227113
rect 125665 227085 125699 227113
rect 125727 227085 125761 227113
rect 125789 227085 125823 227113
rect 125851 227085 140997 227113
rect 141025 227085 141059 227113
rect 141087 227085 141121 227113
rect 141149 227085 141183 227113
rect 141211 227085 156357 227113
rect 156385 227085 156419 227113
rect 156447 227085 156481 227113
rect 156509 227085 156543 227113
rect 156571 227085 171717 227113
rect 171745 227085 171779 227113
rect 171807 227085 171841 227113
rect 171869 227085 171903 227113
rect 171931 227085 187077 227113
rect 187105 227085 187139 227113
rect 187167 227085 187201 227113
rect 187229 227085 187263 227113
rect 187291 227085 202437 227113
rect 202465 227085 202499 227113
rect 202527 227085 202561 227113
rect 202589 227085 202623 227113
rect 202651 227085 217797 227113
rect 217825 227085 217859 227113
rect 217887 227085 217921 227113
rect 217949 227085 217983 227113
rect 218011 227085 233157 227113
rect 233185 227085 233219 227113
rect 233247 227085 233281 227113
rect 233309 227085 233343 227113
rect 233371 227085 248517 227113
rect 248545 227085 248579 227113
rect 248607 227085 248641 227113
rect 248669 227085 248703 227113
rect 248731 227085 263877 227113
rect 263905 227085 263939 227113
rect 263967 227085 264001 227113
rect 264029 227085 264063 227113
rect 264091 227085 279237 227113
rect 279265 227085 279299 227113
rect 279327 227085 279361 227113
rect 279389 227085 279423 227113
rect 279451 227085 294597 227113
rect 294625 227085 294659 227113
rect 294687 227085 294721 227113
rect 294749 227085 294783 227113
rect 294811 227085 298248 227113
rect 298276 227085 298310 227113
rect 298338 227085 298372 227113
rect 298400 227085 298434 227113
rect 298462 227085 298990 227113
rect -958 227051 298990 227085
rect -958 227023 -430 227051
rect -402 227023 -368 227051
rect -340 227023 -306 227051
rect -278 227023 -244 227051
rect -216 227023 2757 227051
rect 2785 227023 2819 227051
rect 2847 227023 2881 227051
rect 2909 227023 2943 227051
rect 2971 227023 18117 227051
rect 18145 227023 18179 227051
rect 18207 227023 18241 227051
rect 18269 227023 18303 227051
rect 18331 227023 33477 227051
rect 33505 227023 33539 227051
rect 33567 227023 33601 227051
rect 33629 227023 33663 227051
rect 33691 227023 48837 227051
rect 48865 227023 48899 227051
rect 48927 227023 48961 227051
rect 48989 227023 49023 227051
rect 49051 227023 64197 227051
rect 64225 227023 64259 227051
rect 64287 227023 64321 227051
rect 64349 227023 64383 227051
rect 64411 227023 79557 227051
rect 79585 227023 79619 227051
rect 79647 227023 79681 227051
rect 79709 227023 79743 227051
rect 79771 227023 94917 227051
rect 94945 227023 94979 227051
rect 95007 227023 95041 227051
rect 95069 227023 95103 227051
rect 95131 227023 110277 227051
rect 110305 227023 110339 227051
rect 110367 227023 110401 227051
rect 110429 227023 110463 227051
rect 110491 227023 125637 227051
rect 125665 227023 125699 227051
rect 125727 227023 125761 227051
rect 125789 227023 125823 227051
rect 125851 227023 140997 227051
rect 141025 227023 141059 227051
rect 141087 227023 141121 227051
rect 141149 227023 141183 227051
rect 141211 227023 156357 227051
rect 156385 227023 156419 227051
rect 156447 227023 156481 227051
rect 156509 227023 156543 227051
rect 156571 227023 171717 227051
rect 171745 227023 171779 227051
rect 171807 227023 171841 227051
rect 171869 227023 171903 227051
rect 171931 227023 187077 227051
rect 187105 227023 187139 227051
rect 187167 227023 187201 227051
rect 187229 227023 187263 227051
rect 187291 227023 202437 227051
rect 202465 227023 202499 227051
rect 202527 227023 202561 227051
rect 202589 227023 202623 227051
rect 202651 227023 217797 227051
rect 217825 227023 217859 227051
rect 217887 227023 217921 227051
rect 217949 227023 217983 227051
rect 218011 227023 233157 227051
rect 233185 227023 233219 227051
rect 233247 227023 233281 227051
rect 233309 227023 233343 227051
rect 233371 227023 248517 227051
rect 248545 227023 248579 227051
rect 248607 227023 248641 227051
rect 248669 227023 248703 227051
rect 248731 227023 263877 227051
rect 263905 227023 263939 227051
rect 263967 227023 264001 227051
rect 264029 227023 264063 227051
rect 264091 227023 279237 227051
rect 279265 227023 279299 227051
rect 279327 227023 279361 227051
rect 279389 227023 279423 227051
rect 279451 227023 294597 227051
rect 294625 227023 294659 227051
rect 294687 227023 294721 227051
rect 294749 227023 294783 227051
rect 294811 227023 298248 227051
rect 298276 227023 298310 227051
rect 298338 227023 298372 227051
rect 298400 227023 298434 227051
rect 298462 227023 298990 227051
rect -958 226989 298990 227023
rect -958 226961 -430 226989
rect -402 226961 -368 226989
rect -340 226961 -306 226989
rect -278 226961 -244 226989
rect -216 226961 2757 226989
rect 2785 226961 2819 226989
rect 2847 226961 2881 226989
rect 2909 226961 2943 226989
rect 2971 226961 18117 226989
rect 18145 226961 18179 226989
rect 18207 226961 18241 226989
rect 18269 226961 18303 226989
rect 18331 226961 33477 226989
rect 33505 226961 33539 226989
rect 33567 226961 33601 226989
rect 33629 226961 33663 226989
rect 33691 226961 48837 226989
rect 48865 226961 48899 226989
rect 48927 226961 48961 226989
rect 48989 226961 49023 226989
rect 49051 226961 64197 226989
rect 64225 226961 64259 226989
rect 64287 226961 64321 226989
rect 64349 226961 64383 226989
rect 64411 226961 79557 226989
rect 79585 226961 79619 226989
rect 79647 226961 79681 226989
rect 79709 226961 79743 226989
rect 79771 226961 94917 226989
rect 94945 226961 94979 226989
rect 95007 226961 95041 226989
rect 95069 226961 95103 226989
rect 95131 226961 110277 226989
rect 110305 226961 110339 226989
rect 110367 226961 110401 226989
rect 110429 226961 110463 226989
rect 110491 226961 125637 226989
rect 125665 226961 125699 226989
rect 125727 226961 125761 226989
rect 125789 226961 125823 226989
rect 125851 226961 140997 226989
rect 141025 226961 141059 226989
rect 141087 226961 141121 226989
rect 141149 226961 141183 226989
rect 141211 226961 156357 226989
rect 156385 226961 156419 226989
rect 156447 226961 156481 226989
rect 156509 226961 156543 226989
rect 156571 226961 171717 226989
rect 171745 226961 171779 226989
rect 171807 226961 171841 226989
rect 171869 226961 171903 226989
rect 171931 226961 187077 226989
rect 187105 226961 187139 226989
rect 187167 226961 187201 226989
rect 187229 226961 187263 226989
rect 187291 226961 202437 226989
rect 202465 226961 202499 226989
rect 202527 226961 202561 226989
rect 202589 226961 202623 226989
rect 202651 226961 217797 226989
rect 217825 226961 217859 226989
rect 217887 226961 217921 226989
rect 217949 226961 217983 226989
rect 218011 226961 233157 226989
rect 233185 226961 233219 226989
rect 233247 226961 233281 226989
rect 233309 226961 233343 226989
rect 233371 226961 248517 226989
rect 248545 226961 248579 226989
rect 248607 226961 248641 226989
rect 248669 226961 248703 226989
rect 248731 226961 263877 226989
rect 263905 226961 263939 226989
rect 263967 226961 264001 226989
rect 264029 226961 264063 226989
rect 264091 226961 279237 226989
rect 279265 226961 279299 226989
rect 279327 226961 279361 226989
rect 279389 226961 279423 226989
rect 279451 226961 294597 226989
rect 294625 226961 294659 226989
rect 294687 226961 294721 226989
rect 294749 226961 294783 226989
rect 294811 226961 298248 226989
rect 298276 226961 298310 226989
rect 298338 226961 298372 226989
rect 298400 226961 298434 226989
rect 298462 226961 298990 226989
rect -958 226913 298990 226961
rect -958 221175 298990 221223
rect -958 221147 -910 221175
rect -882 221147 -848 221175
rect -820 221147 -786 221175
rect -758 221147 -724 221175
rect -696 221147 4617 221175
rect 4645 221147 4679 221175
rect 4707 221147 4741 221175
rect 4769 221147 4803 221175
rect 4831 221147 19977 221175
rect 20005 221147 20039 221175
rect 20067 221147 20101 221175
rect 20129 221147 20163 221175
rect 20191 221147 35337 221175
rect 35365 221147 35399 221175
rect 35427 221147 35461 221175
rect 35489 221147 35523 221175
rect 35551 221147 50697 221175
rect 50725 221147 50759 221175
rect 50787 221147 50821 221175
rect 50849 221147 50883 221175
rect 50911 221147 66057 221175
rect 66085 221147 66119 221175
rect 66147 221147 66181 221175
rect 66209 221147 66243 221175
rect 66271 221147 81417 221175
rect 81445 221147 81479 221175
rect 81507 221147 81541 221175
rect 81569 221147 81603 221175
rect 81631 221147 96777 221175
rect 96805 221147 96839 221175
rect 96867 221147 96901 221175
rect 96929 221147 96963 221175
rect 96991 221147 112137 221175
rect 112165 221147 112199 221175
rect 112227 221147 112261 221175
rect 112289 221147 112323 221175
rect 112351 221147 127497 221175
rect 127525 221147 127559 221175
rect 127587 221147 127621 221175
rect 127649 221147 127683 221175
rect 127711 221147 142857 221175
rect 142885 221147 142919 221175
rect 142947 221147 142981 221175
rect 143009 221147 143043 221175
rect 143071 221147 158217 221175
rect 158245 221147 158279 221175
rect 158307 221147 158341 221175
rect 158369 221147 158403 221175
rect 158431 221147 173577 221175
rect 173605 221147 173639 221175
rect 173667 221147 173701 221175
rect 173729 221147 173763 221175
rect 173791 221147 188937 221175
rect 188965 221147 188999 221175
rect 189027 221147 189061 221175
rect 189089 221147 189123 221175
rect 189151 221147 204297 221175
rect 204325 221147 204359 221175
rect 204387 221147 204421 221175
rect 204449 221147 204483 221175
rect 204511 221147 219657 221175
rect 219685 221147 219719 221175
rect 219747 221147 219781 221175
rect 219809 221147 219843 221175
rect 219871 221147 235017 221175
rect 235045 221147 235079 221175
rect 235107 221147 235141 221175
rect 235169 221147 235203 221175
rect 235231 221147 250377 221175
rect 250405 221147 250439 221175
rect 250467 221147 250501 221175
rect 250529 221147 250563 221175
rect 250591 221147 265737 221175
rect 265765 221147 265799 221175
rect 265827 221147 265861 221175
rect 265889 221147 265923 221175
rect 265951 221147 281097 221175
rect 281125 221147 281159 221175
rect 281187 221147 281221 221175
rect 281249 221147 281283 221175
rect 281311 221147 296457 221175
rect 296485 221147 296519 221175
rect 296547 221147 296581 221175
rect 296609 221147 296643 221175
rect 296671 221147 298728 221175
rect 298756 221147 298790 221175
rect 298818 221147 298852 221175
rect 298880 221147 298914 221175
rect 298942 221147 298990 221175
rect -958 221113 298990 221147
rect -958 221085 -910 221113
rect -882 221085 -848 221113
rect -820 221085 -786 221113
rect -758 221085 -724 221113
rect -696 221085 4617 221113
rect 4645 221085 4679 221113
rect 4707 221085 4741 221113
rect 4769 221085 4803 221113
rect 4831 221085 19977 221113
rect 20005 221085 20039 221113
rect 20067 221085 20101 221113
rect 20129 221085 20163 221113
rect 20191 221085 35337 221113
rect 35365 221085 35399 221113
rect 35427 221085 35461 221113
rect 35489 221085 35523 221113
rect 35551 221085 50697 221113
rect 50725 221085 50759 221113
rect 50787 221085 50821 221113
rect 50849 221085 50883 221113
rect 50911 221085 66057 221113
rect 66085 221085 66119 221113
rect 66147 221085 66181 221113
rect 66209 221085 66243 221113
rect 66271 221085 81417 221113
rect 81445 221085 81479 221113
rect 81507 221085 81541 221113
rect 81569 221085 81603 221113
rect 81631 221085 96777 221113
rect 96805 221085 96839 221113
rect 96867 221085 96901 221113
rect 96929 221085 96963 221113
rect 96991 221085 112137 221113
rect 112165 221085 112199 221113
rect 112227 221085 112261 221113
rect 112289 221085 112323 221113
rect 112351 221085 127497 221113
rect 127525 221085 127559 221113
rect 127587 221085 127621 221113
rect 127649 221085 127683 221113
rect 127711 221085 142857 221113
rect 142885 221085 142919 221113
rect 142947 221085 142981 221113
rect 143009 221085 143043 221113
rect 143071 221085 158217 221113
rect 158245 221085 158279 221113
rect 158307 221085 158341 221113
rect 158369 221085 158403 221113
rect 158431 221085 173577 221113
rect 173605 221085 173639 221113
rect 173667 221085 173701 221113
rect 173729 221085 173763 221113
rect 173791 221085 188937 221113
rect 188965 221085 188999 221113
rect 189027 221085 189061 221113
rect 189089 221085 189123 221113
rect 189151 221085 204297 221113
rect 204325 221085 204359 221113
rect 204387 221085 204421 221113
rect 204449 221085 204483 221113
rect 204511 221085 219657 221113
rect 219685 221085 219719 221113
rect 219747 221085 219781 221113
rect 219809 221085 219843 221113
rect 219871 221085 235017 221113
rect 235045 221085 235079 221113
rect 235107 221085 235141 221113
rect 235169 221085 235203 221113
rect 235231 221085 250377 221113
rect 250405 221085 250439 221113
rect 250467 221085 250501 221113
rect 250529 221085 250563 221113
rect 250591 221085 265737 221113
rect 265765 221085 265799 221113
rect 265827 221085 265861 221113
rect 265889 221085 265923 221113
rect 265951 221085 281097 221113
rect 281125 221085 281159 221113
rect 281187 221085 281221 221113
rect 281249 221085 281283 221113
rect 281311 221085 296457 221113
rect 296485 221085 296519 221113
rect 296547 221085 296581 221113
rect 296609 221085 296643 221113
rect 296671 221085 298728 221113
rect 298756 221085 298790 221113
rect 298818 221085 298852 221113
rect 298880 221085 298914 221113
rect 298942 221085 298990 221113
rect -958 221051 298990 221085
rect -958 221023 -910 221051
rect -882 221023 -848 221051
rect -820 221023 -786 221051
rect -758 221023 -724 221051
rect -696 221023 4617 221051
rect 4645 221023 4679 221051
rect 4707 221023 4741 221051
rect 4769 221023 4803 221051
rect 4831 221023 19977 221051
rect 20005 221023 20039 221051
rect 20067 221023 20101 221051
rect 20129 221023 20163 221051
rect 20191 221023 35337 221051
rect 35365 221023 35399 221051
rect 35427 221023 35461 221051
rect 35489 221023 35523 221051
rect 35551 221023 50697 221051
rect 50725 221023 50759 221051
rect 50787 221023 50821 221051
rect 50849 221023 50883 221051
rect 50911 221023 66057 221051
rect 66085 221023 66119 221051
rect 66147 221023 66181 221051
rect 66209 221023 66243 221051
rect 66271 221023 81417 221051
rect 81445 221023 81479 221051
rect 81507 221023 81541 221051
rect 81569 221023 81603 221051
rect 81631 221023 96777 221051
rect 96805 221023 96839 221051
rect 96867 221023 96901 221051
rect 96929 221023 96963 221051
rect 96991 221023 112137 221051
rect 112165 221023 112199 221051
rect 112227 221023 112261 221051
rect 112289 221023 112323 221051
rect 112351 221023 127497 221051
rect 127525 221023 127559 221051
rect 127587 221023 127621 221051
rect 127649 221023 127683 221051
rect 127711 221023 142857 221051
rect 142885 221023 142919 221051
rect 142947 221023 142981 221051
rect 143009 221023 143043 221051
rect 143071 221023 158217 221051
rect 158245 221023 158279 221051
rect 158307 221023 158341 221051
rect 158369 221023 158403 221051
rect 158431 221023 173577 221051
rect 173605 221023 173639 221051
rect 173667 221023 173701 221051
rect 173729 221023 173763 221051
rect 173791 221023 188937 221051
rect 188965 221023 188999 221051
rect 189027 221023 189061 221051
rect 189089 221023 189123 221051
rect 189151 221023 204297 221051
rect 204325 221023 204359 221051
rect 204387 221023 204421 221051
rect 204449 221023 204483 221051
rect 204511 221023 219657 221051
rect 219685 221023 219719 221051
rect 219747 221023 219781 221051
rect 219809 221023 219843 221051
rect 219871 221023 235017 221051
rect 235045 221023 235079 221051
rect 235107 221023 235141 221051
rect 235169 221023 235203 221051
rect 235231 221023 250377 221051
rect 250405 221023 250439 221051
rect 250467 221023 250501 221051
rect 250529 221023 250563 221051
rect 250591 221023 265737 221051
rect 265765 221023 265799 221051
rect 265827 221023 265861 221051
rect 265889 221023 265923 221051
rect 265951 221023 281097 221051
rect 281125 221023 281159 221051
rect 281187 221023 281221 221051
rect 281249 221023 281283 221051
rect 281311 221023 296457 221051
rect 296485 221023 296519 221051
rect 296547 221023 296581 221051
rect 296609 221023 296643 221051
rect 296671 221023 298728 221051
rect 298756 221023 298790 221051
rect 298818 221023 298852 221051
rect 298880 221023 298914 221051
rect 298942 221023 298990 221051
rect -958 220989 298990 221023
rect -958 220961 -910 220989
rect -882 220961 -848 220989
rect -820 220961 -786 220989
rect -758 220961 -724 220989
rect -696 220961 4617 220989
rect 4645 220961 4679 220989
rect 4707 220961 4741 220989
rect 4769 220961 4803 220989
rect 4831 220961 19977 220989
rect 20005 220961 20039 220989
rect 20067 220961 20101 220989
rect 20129 220961 20163 220989
rect 20191 220961 35337 220989
rect 35365 220961 35399 220989
rect 35427 220961 35461 220989
rect 35489 220961 35523 220989
rect 35551 220961 50697 220989
rect 50725 220961 50759 220989
rect 50787 220961 50821 220989
rect 50849 220961 50883 220989
rect 50911 220961 66057 220989
rect 66085 220961 66119 220989
rect 66147 220961 66181 220989
rect 66209 220961 66243 220989
rect 66271 220961 81417 220989
rect 81445 220961 81479 220989
rect 81507 220961 81541 220989
rect 81569 220961 81603 220989
rect 81631 220961 96777 220989
rect 96805 220961 96839 220989
rect 96867 220961 96901 220989
rect 96929 220961 96963 220989
rect 96991 220961 112137 220989
rect 112165 220961 112199 220989
rect 112227 220961 112261 220989
rect 112289 220961 112323 220989
rect 112351 220961 127497 220989
rect 127525 220961 127559 220989
rect 127587 220961 127621 220989
rect 127649 220961 127683 220989
rect 127711 220961 142857 220989
rect 142885 220961 142919 220989
rect 142947 220961 142981 220989
rect 143009 220961 143043 220989
rect 143071 220961 158217 220989
rect 158245 220961 158279 220989
rect 158307 220961 158341 220989
rect 158369 220961 158403 220989
rect 158431 220961 173577 220989
rect 173605 220961 173639 220989
rect 173667 220961 173701 220989
rect 173729 220961 173763 220989
rect 173791 220961 188937 220989
rect 188965 220961 188999 220989
rect 189027 220961 189061 220989
rect 189089 220961 189123 220989
rect 189151 220961 204297 220989
rect 204325 220961 204359 220989
rect 204387 220961 204421 220989
rect 204449 220961 204483 220989
rect 204511 220961 219657 220989
rect 219685 220961 219719 220989
rect 219747 220961 219781 220989
rect 219809 220961 219843 220989
rect 219871 220961 235017 220989
rect 235045 220961 235079 220989
rect 235107 220961 235141 220989
rect 235169 220961 235203 220989
rect 235231 220961 250377 220989
rect 250405 220961 250439 220989
rect 250467 220961 250501 220989
rect 250529 220961 250563 220989
rect 250591 220961 265737 220989
rect 265765 220961 265799 220989
rect 265827 220961 265861 220989
rect 265889 220961 265923 220989
rect 265951 220961 281097 220989
rect 281125 220961 281159 220989
rect 281187 220961 281221 220989
rect 281249 220961 281283 220989
rect 281311 220961 296457 220989
rect 296485 220961 296519 220989
rect 296547 220961 296581 220989
rect 296609 220961 296643 220989
rect 296671 220961 298728 220989
rect 298756 220961 298790 220989
rect 298818 220961 298852 220989
rect 298880 220961 298914 220989
rect 298942 220961 298990 220989
rect -958 220913 298990 220961
rect -958 218175 298990 218223
rect -958 218147 -430 218175
rect -402 218147 -368 218175
rect -340 218147 -306 218175
rect -278 218147 -244 218175
rect -216 218147 2757 218175
rect 2785 218147 2819 218175
rect 2847 218147 2881 218175
rect 2909 218147 2943 218175
rect 2971 218147 18117 218175
rect 18145 218147 18179 218175
rect 18207 218147 18241 218175
rect 18269 218147 18303 218175
rect 18331 218147 33477 218175
rect 33505 218147 33539 218175
rect 33567 218147 33601 218175
rect 33629 218147 33663 218175
rect 33691 218147 48837 218175
rect 48865 218147 48899 218175
rect 48927 218147 48961 218175
rect 48989 218147 49023 218175
rect 49051 218147 64197 218175
rect 64225 218147 64259 218175
rect 64287 218147 64321 218175
rect 64349 218147 64383 218175
rect 64411 218147 79557 218175
rect 79585 218147 79619 218175
rect 79647 218147 79681 218175
rect 79709 218147 79743 218175
rect 79771 218147 94917 218175
rect 94945 218147 94979 218175
rect 95007 218147 95041 218175
rect 95069 218147 95103 218175
rect 95131 218147 110277 218175
rect 110305 218147 110339 218175
rect 110367 218147 110401 218175
rect 110429 218147 110463 218175
rect 110491 218147 125637 218175
rect 125665 218147 125699 218175
rect 125727 218147 125761 218175
rect 125789 218147 125823 218175
rect 125851 218147 140997 218175
rect 141025 218147 141059 218175
rect 141087 218147 141121 218175
rect 141149 218147 141183 218175
rect 141211 218147 156357 218175
rect 156385 218147 156419 218175
rect 156447 218147 156481 218175
rect 156509 218147 156543 218175
rect 156571 218147 171717 218175
rect 171745 218147 171779 218175
rect 171807 218147 171841 218175
rect 171869 218147 171903 218175
rect 171931 218147 187077 218175
rect 187105 218147 187139 218175
rect 187167 218147 187201 218175
rect 187229 218147 187263 218175
rect 187291 218147 202437 218175
rect 202465 218147 202499 218175
rect 202527 218147 202561 218175
rect 202589 218147 202623 218175
rect 202651 218147 217797 218175
rect 217825 218147 217859 218175
rect 217887 218147 217921 218175
rect 217949 218147 217983 218175
rect 218011 218147 233157 218175
rect 233185 218147 233219 218175
rect 233247 218147 233281 218175
rect 233309 218147 233343 218175
rect 233371 218147 248517 218175
rect 248545 218147 248579 218175
rect 248607 218147 248641 218175
rect 248669 218147 248703 218175
rect 248731 218147 263877 218175
rect 263905 218147 263939 218175
rect 263967 218147 264001 218175
rect 264029 218147 264063 218175
rect 264091 218147 279237 218175
rect 279265 218147 279299 218175
rect 279327 218147 279361 218175
rect 279389 218147 279423 218175
rect 279451 218147 294597 218175
rect 294625 218147 294659 218175
rect 294687 218147 294721 218175
rect 294749 218147 294783 218175
rect 294811 218147 298248 218175
rect 298276 218147 298310 218175
rect 298338 218147 298372 218175
rect 298400 218147 298434 218175
rect 298462 218147 298990 218175
rect -958 218113 298990 218147
rect -958 218085 -430 218113
rect -402 218085 -368 218113
rect -340 218085 -306 218113
rect -278 218085 -244 218113
rect -216 218085 2757 218113
rect 2785 218085 2819 218113
rect 2847 218085 2881 218113
rect 2909 218085 2943 218113
rect 2971 218085 18117 218113
rect 18145 218085 18179 218113
rect 18207 218085 18241 218113
rect 18269 218085 18303 218113
rect 18331 218085 33477 218113
rect 33505 218085 33539 218113
rect 33567 218085 33601 218113
rect 33629 218085 33663 218113
rect 33691 218085 48837 218113
rect 48865 218085 48899 218113
rect 48927 218085 48961 218113
rect 48989 218085 49023 218113
rect 49051 218085 64197 218113
rect 64225 218085 64259 218113
rect 64287 218085 64321 218113
rect 64349 218085 64383 218113
rect 64411 218085 79557 218113
rect 79585 218085 79619 218113
rect 79647 218085 79681 218113
rect 79709 218085 79743 218113
rect 79771 218085 94917 218113
rect 94945 218085 94979 218113
rect 95007 218085 95041 218113
rect 95069 218085 95103 218113
rect 95131 218085 110277 218113
rect 110305 218085 110339 218113
rect 110367 218085 110401 218113
rect 110429 218085 110463 218113
rect 110491 218085 125637 218113
rect 125665 218085 125699 218113
rect 125727 218085 125761 218113
rect 125789 218085 125823 218113
rect 125851 218085 140997 218113
rect 141025 218085 141059 218113
rect 141087 218085 141121 218113
rect 141149 218085 141183 218113
rect 141211 218085 156357 218113
rect 156385 218085 156419 218113
rect 156447 218085 156481 218113
rect 156509 218085 156543 218113
rect 156571 218085 171717 218113
rect 171745 218085 171779 218113
rect 171807 218085 171841 218113
rect 171869 218085 171903 218113
rect 171931 218085 187077 218113
rect 187105 218085 187139 218113
rect 187167 218085 187201 218113
rect 187229 218085 187263 218113
rect 187291 218085 202437 218113
rect 202465 218085 202499 218113
rect 202527 218085 202561 218113
rect 202589 218085 202623 218113
rect 202651 218085 217797 218113
rect 217825 218085 217859 218113
rect 217887 218085 217921 218113
rect 217949 218085 217983 218113
rect 218011 218085 233157 218113
rect 233185 218085 233219 218113
rect 233247 218085 233281 218113
rect 233309 218085 233343 218113
rect 233371 218085 248517 218113
rect 248545 218085 248579 218113
rect 248607 218085 248641 218113
rect 248669 218085 248703 218113
rect 248731 218085 263877 218113
rect 263905 218085 263939 218113
rect 263967 218085 264001 218113
rect 264029 218085 264063 218113
rect 264091 218085 279237 218113
rect 279265 218085 279299 218113
rect 279327 218085 279361 218113
rect 279389 218085 279423 218113
rect 279451 218085 294597 218113
rect 294625 218085 294659 218113
rect 294687 218085 294721 218113
rect 294749 218085 294783 218113
rect 294811 218085 298248 218113
rect 298276 218085 298310 218113
rect 298338 218085 298372 218113
rect 298400 218085 298434 218113
rect 298462 218085 298990 218113
rect -958 218051 298990 218085
rect -958 218023 -430 218051
rect -402 218023 -368 218051
rect -340 218023 -306 218051
rect -278 218023 -244 218051
rect -216 218023 2757 218051
rect 2785 218023 2819 218051
rect 2847 218023 2881 218051
rect 2909 218023 2943 218051
rect 2971 218023 18117 218051
rect 18145 218023 18179 218051
rect 18207 218023 18241 218051
rect 18269 218023 18303 218051
rect 18331 218023 33477 218051
rect 33505 218023 33539 218051
rect 33567 218023 33601 218051
rect 33629 218023 33663 218051
rect 33691 218023 48837 218051
rect 48865 218023 48899 218051
rect 48927 218023 48961 218051
rect 48989 218023 49023 218051
rect 49051 218023 64197 218051
rect 64225 218023 64259 218051
rect 64287 218023 64321 218051
rect 64349 218023 64383 218051
rect 64411 218023 79557 218051
rect 79585 218023 79619 218051
rect 79647 218023 79681 218051
rect 79709 218023 79743 218051
rect 79771 218023 94917 218051
rect 94945 218023 94979 218051
rect 95007 218023 95041 218051
rect 95069 218023 95103 218051
rect 95131 218023 110277 218051
rect 110305 218023 110339 218051
rect 110367 218023 110401 218051
rect 110429 218023 110463 218051
rect 110491 218023 125637 218051
rect 125665 218023 125699 218051
rect 125727 218023 125761 218051
rect 125789 218023 125823 218051
rect 125851 218023 140997 218051
rect 141025 218023 141059 218051
rect 141087 218023 141121 218051
rect 141149 218023 141183 218051
rect 141211 218023 156357 218051
rect 156385 218023 156419 218051
rect 156447 218023 156481 218051
rect 156509 218023 156543 218051
rect 156571 218023 171717 218051
rect 171745 218023 171779 218051
rect 171807 218023 171841 218051
rect 171869 218023 171903 218051
rect 171931 218023 187077 218051
rect 187105 218023 187139 218051
rect 187167 218023 187201 218051
rect 187229 218023 187263 218051
rect 187291 218023 202437 218051
rect 202465 218023 202499 218051
rect 202527 218023 202561 218051
rect 202589 218023 202623 218051
rect 202651 218023 217797 218051
rect 217825 218023 217859 218051
rect 217887 218023 217921 218051
rect 217949 218023 217983 218051
rect 218011 218023 233157 218051
rect 233185 218023 233219 218051
rect 233247 218023 233281 218051
rect 233309 218023 233343 218051
rect 233371 218023 248517 218051
rect 248545 218023 248579 218051
rect 248607 218023 248641 218051
rect 248669 218023 248703 218051
rect 248731 218023 263877 218051
rect 263905 218023 263939 218051
rect 263967 218023 264001 218051
rect 264029 218023 264063 218051
rect 264091 218023 279237 218051
rect 279265 218023 279299 218051
rect 279327 218023 279361 218051
rect 279389 218023 279423 218051
rect 279451 218023 294597 218051
rect 294625 218023 294659 218051
rect 294687 218023 294721 218051
rect 294749 218023 294783 218051
rect 294811 218023 298248 218051
rect 298276 218023 298310 218051
rect 298338 218023 298372 218051
rect 298400 218023 298434 218051
rect 298462 218023 298990 218051
rect -958 217989 298990 218023
rect -958 217961 -430 217989
rect -402 217961 -368 217989
rect -340 217961 -306 217989
rect -278 217961 -244 217989
rect -216 217961 2757 217989
rect 2785 217961 2819 217989
rect 2847 217961 2881 217989
rect 2909 217961 2943 217989
rect 2971 217961 18117 217989
rect 18145 217961 18179 217989
rect 18207 217961 18241 217989
rect 18269 217961 18303 217989
rect 18331 217961 33477 217989
rect 33505 217961 33539 217989
rect 33567 217961 33601 217989
rect 33629 217961 33663 217989
rect 33691 217961 48837 217989
rect 48865 217961 48899 217989
rect 48927 217961 48961 217989
rect 48989 217961 49023 217989
rect 49051 217961 64197 217989
rect 64225 217961 64259 217989
rect 64287 217961 64321 217989
rect 64349 217961 64383 217989
rect 64411 217961 79557 217989
rect 79585 217961 79619 217989
rect 79647 217961 79681 217989
rect 79709 217961 79743 217989
rect 79771 217961 94917 217989
rect 94945 217961 94979 217989
rect 95007 217961 95041 217989
rect 95069 217961 95103 217989
rect 95131 217961 110277 217989
rect 110305 217961 110339 217989
rect 110367 217961 110401 217989
rect 110429 217961 110463 217989
rect 110491 217961 125637 217989
rect 125665 217961 125699 217989
rect 125727 217961 125761 217989
rect 125789 217961 125823 217989
rect 125851 217961 140997 217989
rect 141025 217961 141059 217989
rect 141087 217961 141121 217989
rect 141149 217961 141183 217989
rect 141211 217961 156357 217989
rect 156385 217961 156419 217989
rect 156447 217961 156481 217989
rect 156509 217961 156543 217989
rect 156571 217961 171717 217989
rect 171745 217961 171779 217989
rect 171807 217961 171841 217989
rect 171869 217961 171903 217989
rect 171931 217961 187077 217989
rect 187105 217961 187139 217989
rect 187167 217961 187201 217989
rect 187229 217961 187263 217989
rect 187291 217961 202437 217989
rect 202465 217961 202499 217989
rect 202527 217961 202561 217989
rect 202589 217961 202623 217989
rect 202651 217961 217797 217989
rect 217825 217961 217859 217989
rect 217887 217961 217921 217989
rect 217949 217961 217983 217989
rect 218011 217961 233157 217989
rect 233185 217961 233219 217989
rect 233247 217961 233281 217989
rect 233309 217961 233343 217989
rect 233371 217961 248517 217989
rect 248545 217961 248579 217989
rect 248607 217961 248641 217989
rect 248669 217961 248703 217989
rect 248731 217961 263877 217989
rect 263905 217961 263939 217989
rect 263967 217961 264001 217989
rect 264029 217961 264063 217989
rect 264091 217961 279237 217989
rect 279265 217961 279299 217989
rect 279327 217961 279361 217989
rect 279389 217961 279423 217989
rect 279451 217961 294597 217989
rect 294625 217961 294659 217989
rect 294687 217961 294721 217989
rect 294749 217961 294783 217989
rect 294811 217961 298248 217989
rect 298276 217961 298310 217989
rect 298338 217961 298372 217989
rect 298400 217961 298434 217989
rect 298462 217961 298990 217989
rect -958 217913 298990 217961
rect -958 212175 298990 212223
rect -958 212147 -910 212175
rect -882 212147 -848 212175
rect -820 212147 -786 212175
rect -758 212147 -724 212175
rect -696 212147 4617 212175
rect 4645 212147 4679 212175
rect 4707 212147 4741 212175
rect 4769 212147 4803 212175
rect 4831 212147 19977 212175
rect 20005 212147 20039 212175
rect 20067 212147 20101 212175
rect 20129 212147 20163 212175
rect 20191 212147 35337 212175
rect 35365 212147 35399 212175
rect 35427 212147 35461 212175
rect 35489 212147 35523 212175
rect 35551 212147 50697 212175
rect 50725 212147 50759 212175
rect 50787 212147 50821 212175
rect 50849 212147 50883 212175
rect 50911 212147 66057 212175
rect 66085 212147 66119 212175
rect 66147 212147 66181 212175
rect 66209 212147 66243 212175
rect 66271 212147 81417 212175
rect 81445 212147 81479 212175
rect 81507 212147 81541 212175
rect 81569 212147 81603 212175
rect 81631 212147 96777 212175
rect 96805 212147 96839 212175
rect 96867 212147 96901 212175
rect 96929 212147 96963 212175
rect 96991 212147 112137 212175
rect 112165 212147 112199 212175
rect 112227 212147 112261 212175
rect 112289 212147 112323 212175
rect 112351 212147 127497 212175
rect 127525 212147 127559 212175
rect 127587 212147 127621 212175
rect 127649 212147 127683 212175
rect 127711 212147 142857 212175
rect 142885 212147 142919 212175
rect 142947 212147 142981 212175
rect 143009 212147 143043 212175
rect 143071 212147 158217 212175
rect 158245 212147 158279 212175
rect 158307 212147 158341 212175
rect 158369 212147 158403 212175
rect 158431 212147 173577 212175
rect 173605 212147 173639 212175
rect 173667 212147 173701 212175
rect 173729 212147 173763 212175
rect 173791 212147 188937 212175
rect 188965 212147 188999 212175
rect 189027 212147 189061 212175
rect 189089 212147 189123 212175
rect 189151 212147 204297 212175
rect 204325 212147 204359 212175
rect 204387 212147 204421 212175
rect 204449 212147 204483 212175
rect 204511 212147 219657 212175
rect 219685 212147 219719 212175
rect 219747 212147 219781 212175
rect 219809 212147 219843 212175
rect 219871 212147 235017 212175
rect 235045 212147 235079 212175
rect 235107 212147 235141 212175
rect 235169 212147 235203 212175
rect 235231 212147 250377 212175
rect 250405 212147 250439 212175
rect 250467 212147 250501 212175
rect 250529 212147 250563 212175
rect 250591 212147 265737 212175
rect 265765 212147 265799 212175
rect 265827 212147 265861 212175
rect 265889 212147 265923 212175
rect 265951 212147 281097 212175
rect 281125 212147 281159 212175
rect 281187 212147 281221 212175
rect 281249 212147 281283 212175
rect 281311 212147 296457 212175
rect 296485 212147 296519 212175
rect 296547 212147 296581 212175
rect 296609 212147 296643 212175
rect 296671 212147 298728 212175
rect 298756 212147 298790 212175
rect 298818 212147 298852 212175
rect 298880 212147 298914 212175
rect 298942 212147 298990 212175
rect -958 212113 298990 212147
rect -958 212085 -910 212113
rect -882 212085 -848 212113
rect -820 212085 -786 212113
rect -758 212085 -724 212113
rect -696 212085 4617 212113
rect 4645 212085 4679 212113
rect 4707 212085 4741 212113
rect 4769 212085 4803 212113
rect 4831 212085 19977 212113
rect 20005 212085 20039 212113
rect 20067 212085 20101 212113
rect 20129 212085 20163 212113
rect 20191 212085 35337 212113
rect 35365 212085 35399 212113
rect 35427 212085 35461 212113
rect 35489 212085 35523 212113
rect 35551 212085 50697 212113
rect 50725 212085 50759 212113
rect 50787 212085 50821 212113
rect 50849 212085 50883 212113
rect 50911 212085 66057 212113
rect 66085 212085 66119 212113
rect 66147 212085 66181 212113
rect 66209 212085 66243 212113
rect 66271 212085 81417 212113
rect 81445 212085 81479 212113
rect 81507 212085 81541 212113
rect 81569 212085 81603 212113
rect 81631 212085 96777 212113
rect 96805 212085 96839 212113
rect 96867 212085 96901 212113
rect 96929 212085 96963 212113
rect 96991 212085 112137 212113
rect 112165 212085 112199 212113
rect 112227 212085 112261 212113
rect 112289 212085 112323 212113
rect 112351 212085 127497 212113
rect 127525 212085 127559 212113
rect 127587 212085 127621 212113
rect 127649 212085 127683 212113
rect 127711 212085 142857 212113
rect 142885 212085 142919 212113
rect 142947 212085 142981 212113
rect 143009 212085 143043 212113
rect 143071 212085 158217 212113
rect 158245 212085 158279 212113
rect 158307 212085 158341 212113
rect 158369 212085 158403 212113
rect 158431 212085 173577 212113
rect 173605 212085 173639 212113
rect 173667 212085 173701 212113
rect 173729 212085 173763 212113
rect 173791 212085 188937 212113
rect 188965 212085 188999 212113
rect 189027 212085 189061 212113
rect 189089 212085 189123 212113
rect 189151 212085 204297 212113
rect 204325 212085 204359 212113
rect 204387 212085 204421 212113
rect 204449 212085 204483 212113
rect 204511 212085 219657 212113
rect 219685 212085 219719 212113
rect 219747 212085 219781 212113
rect 219809 212085 219843 212113
rect 219871 212085 235017 212113
rect 235045 212085 235079 212113
rect 235107 212085 235141 212113
rect 235169 212085 235203 212113
rect 235231 212085 250377 212113
rect 250405 212085 250439 212113
rect 250467 212085 250501 212113
rect 250529 212085 250563 212113
rect 250591 212085 265737 212113
rect 265765 212085 265799 212113
rect 265827 212085 265861 212113
rect 265889 212085 265923 212113
rect 265951 212085 281097 212113
rect 281125 212085 281159 212113
rect 281187 212085 281221 212113
rect 281249 212085 281283 212113
rect 281311 212085 296457 212113
rect 296485 212085 296519 212113
rect 296547 212085 296581 212113
rect 296609 212085 296643 212113
rect 296671 212085 298728 212113
rect 298756 212085 298790 212113
rect 298818 212085 298852 212113
rect 298880 212085 298914 212113
rect 298942 212085 298990 212113
rect -958 212051 298990 212085
rect -958 212023 -910 212051
rect -882 212023 -848 212051
rect -820 212023 -786 212051
rect -758 212023 -724 212051
rect -696 212023 4617 212051
rect 4645 212023 4679 212051
rect 4707 212023 4741 212051
rect 4769 212023 4803 212051
rect 4831 212023 19977 212051
rect 20005 212023 20039 212051
rect 20067 212023 20101 212051
rect 20129 212023 20163 212051
rect 20191 212023 35337 212051
rect 35365 212023 35399 212051
rect 35427 212023 35461 212051
rect 35489 212023 35523 212051
rect 35551 212023 50697 212051
rect 50725 212023 50759 212051
rect 50787 212023 50821 212051
rect 50849 212023 50883 212051
rect 50911 212023 66057 212051
rect 66085 212023 66119 212051
rect 66147 212023 66181 212051
rect 66209 212023 66243 212051
rect 66271 212023 81417 212051
rect 81445 212023 81479 212051
rect 81507 212023 81541 212051
rect 81569 212023 81603 212051
rect 81631 212023 96777 212051
rect 96805 212023 96839 212051
rect 96867 212023 96901 212051
rect 96929 212023 96963 212051
rect 96991 212023 112137 212051
rect 112165 212023 112199 212051
rect 112227 212023 112261 212051
rect 112289 212023 112323 212051
rect 112351 212023 127497 212051
rect 127525 212023 127559 212051
rect 127587 212023 127621 212051
rect 127649 212023 127683 212051
rect 127711 212023 142857 212051
rect 142885 212023 142919 212051
rect 142947 212023 142981 212051
rect 143009 212023 143043 212051
rect 143071 212023 158217 212051
rect 158245 212023 158279 212051
rect 158307 212023 158341 212051
rect 158369 212023 158403 212051
rect 158431 212023 173577 212051
rect 173605 212023 173639 212051
rect 173667 212023 173701 212051
rect 173729 212023 173763 212051
rect 173791 212023 188937 212051
rect 188965 212023 188999 212051
rect 189027 212023 189061 212051
rect 189089 212023 189123 212051
rect 189151 212023 204297 212051
rect 204325 212023 204359 212051
rect 204387 212023 204421 212051
rect 204449 212023 204483 212051
rect 204511 212023 219657 212051
rect 219685 212023 219719 212051
rect 219747 212023 219781 212051
rect 219809 212023 219843 212051
rect 219871 212023 235017 212051
rect 235045 212023 235079 212051
rect 235107 212023 235141 212051
rect 235169 212023 235203 212051
rect 235231 212023 250377 212051
rect 250405 212023 250439 212051
rect 250467 212023 250501 212051
rect 250529 212023 250563 212051
rect 250591 212023 265737 212051
rect 265765 212023 265799 212051
rect 265827 212023 265861 212051
rect 265889 212023 265923 212051
rect 265951 212023 281097 212051
rect 281125 212023 281159 212051
rect 281187 212023 281221 212051
rect 281249 212023 281283 212051
rect 281311 212023 296457 212051
rect 296485 212023 296519 212051
rect 296547 212023 296581 212051
rect 296609 212023 296643 212051
rect 296671 212023 298728 212051
rect 298756 212023 298790 212051
rect 298818 212023 298852 212051
rect 298880 212023 298914 212051
rect 298942 212023 298990 212051
rect -958 211989 298990 212023
rect -958 211961 -910 211989
rect -882 211961 -848 211989
rect -820 211961 -786 211989
rect -758 211961 -724 211989
rect -696 211961 4617 211989
rect 4645 211961 4679 211989
rect 4707 211961 4741 211989
rect 4769 211961 4803 211989
rect 4831 211961 19977 211989
rect 20005 211961 20039 211989
rect 20067 211961 20101 211989
rect 20129 211961 20163 211989
rect 20191 211961 35337 211989
rect 35365 211961 35399 211989
rect 35427 211961 35461 211989
rect 35489 211961 35523 211989
rect 35551 211961 50697 211989
rect 50725 211961 50759 211989
rect 50787 211961 50821 211989
rect 50849 211961 50883 211989
rect 50911 211961 66057 211989
rect 66085 211961 66119 211989
rect 66147 211961 66181 211989
rect 66209 211961 66243 211989
rect 66271 211961 81417 211989
rect 81445 211961 81479 211989
rect 81507 211961 81541 211989
rect 81569 211961 81603 211989
rect 81631 211961 96777 211989
rect 96805 211961 96839 211989
rect 96867 211961 96901 211989
rect 96929 211961 96963 211989
rect 96991 211961 112137 211989
rect 112165 211961 112199 211989
rect 112227 211961 112261 211989
rect 112289 211961 112323 211989
rect 112351 211961 127497 211989
rect 127525 211961 127559 211989
rect 127587 211961 127621 211989
rect 127649 211961 127683 211989
rect 127711 211961 142857 211989
rect 142885 211961 142919 211989
rect 142947 211961 142981 211989
rect 143009 211961 143043 211989
rect 143071 211961 158217 211989
rect 158245 211961 158279 211989
rect 158307 211961 158341 211989
rect 158369 211961 158403 211989
rect 158431 211961 173577 211989
rect 173605 211961 173639 211989
rect 173667 211961 173701 211989
rect 173729 211961 173763 211989
rect 173791 211961 188937 211989
rect 188965 211961 188999 211989
rect 189027 211961 189061 211989
rect 189089 211961 189123 211989
rect 189151 211961 204297 211989
rect 204325 211961 204359 211989
rect 204387 211961 204421 211989
rect 204449 211961 204483 211989
rect 204511 211961 219657 211989
rect 219685 211961 219719 211989
rect 219747 211961 219781 211989
rect 219809 211961 219843 211989
rect 219871 211961 235017 211989
rect 235045 211961 235079 211989
rect 235107 211961 235141 211989
rect 235169 211961 235203 211989
rect 235231 211961 250377 211989
rect 250405 211961 250439 211989
rect 250467 211961 250501 211989
rect 250529 211961 250563 211989
rect 250591 211961 265737 211989
rect 265765 211961 265799 211989
rect 265827 211961 265861 211989
rect 265889 211961 265923 211989
rect 265951 211961 281097 211989
rect 281125 211961 281159 211989
rect 281187 211961 281221 211989
rect 281249 211961 281283 211989
rect 281311 211961 296457 211989
rect 296485 211961 296519 211989
rect 296547 211961 296581 211989
rect 296609 211961 296643 211989
rect 296671 211961 298728 211989
rect 298756 211961 298790 211989
rect 298818 211961 298852 211989
rect 298880 211961 298914 211989
rect 298942 211961 298990 211989
rect -958 211913 298990 211961
rect -958 209175 298990 209223
rect -958 209147 -430 209175
rect -402 209147 -368 209175
rect -340 209147 -306 209175
rect -278 209147 -244 209175
rect -216 209147 2757 209175
rect 2785 209147 2819 209175
rect 2847 209147 2881 209175
rect 2909 209147 2943 209175
rect 2971 209147 18117 209175
rect 18145 209147 18179 209175
rect 18207 209147 18241 209175
rect 18269 209147 18303 209175
rect 18331 209147 33477 209175
rect 33505 209147 33539 209175
rect 33567 209147 33601 209175
rect 33629 209147 33663 209175
rect 33691 209147 48837 209175
rect 48865 209147 48899 209175
rect 48927 209147 48961 209175
rect 48989 209147 49023 209175
rect 49051 209147 64197 209175
rect 64225 209147 64259 209175
rect 64287 209147 64321 209175
rect 64349 209147 64383 209175
rect 64411 209147 79557 209175
rect 79585 209147 79619 209175
rect 79647 209147 79681 209175
rect 79709 209147 79743 209175
rect 79771 209147 94917 209175
rect 94945 209147 94979 209175
rect 95007 209147 95041 209175
rect 95069 209147 95103 209175
rect 95131 209147 110277 209175
rect 110305 209147 110339 209175
rect 110367 209147 110401 209175
rect 110429 209147 110463 209175
rect 110491 209147 125637 209175
rect 125665 209147 125699 209175
rect 125727 209147 125761 209175
rect 125789 209147 125823 209175
rect 125851 209147 140997 209175
rect 141025 209147 141059 209175
rect 141087 209147 141121 209175
rect 141149 209147 141183 209175
rect 141211 209147 156357 209175
rect 156385 209147 156419 209175
rect 156447 209147 156481 209175
rect 156509 209147 156543 209175
rect 156571 209147 171717 209175
rect 171745 209147 171779 209175
rect 171807 209147 171841 209175
rect 171869 209147 171903 209175
rect 171931 209147 187077 209175
rect 187105 209147 187139 209175
rect 187167 209147 187201 209175
rect 187229 209147 187263 209175
rect 187291 209147 202437 209175
rect 202465 209147 202499 209175
rect 202527 209147 202561 209175
rect 202589 209147 202623 209175
rect 202651 209147 217797 209175
rect 217825 209147 217859 209175
rect 217887 209147 217921 209175
rect 217949 209147 217983 209175
rect 218011 209147 233157 209175
rect 233185 209147 233219 209175
rect 233247 209147 233281 209175
rect 233309 209147 233343 209175
rect 233371 209147 248517 209175
rect 248545 209147 248579 209175
rect 248607 209147 248641 209175
rect 248669 209147 248703 209175
rect 248731 209147 263877 209175
rect 263905 209147 263939 209175
rect 263967 209147 264001 209175
rect 264029 209147 264063 209175
rect 264091 209147 279237 209175
rect 279265 209147 279299 209175
rect 279327 209147 279361 209175
rect 279389 209147 279423 209175
rect 279451 209147 294597 209175
rect 294625 209147 294659 209175
rect 294687 209147 294721 209175
rect 294749 209147 294783 209175
rect 294811 209147 298248 209175
rect 298276 209147 298310 209175
rect 298338 209147 298372 209175
rect 298400 209147 298434 209175
rect 298462 209147 298990 209175
rect -958 209113 298990 209147
rect -958 209085 -430 209113
rect -402 209085 -368 209113
rect -340 209085 -306 209113
rect -278 209085 -244 209113
rect -216 209085 2757 209113
rect 2785 209085 2819 209113
rect 2847 209085 2881 209113
rect 2909 209085 2943 209113
rect 2971 209085 18117 209113
rect 18145 209085 18179 209113
rect 18207 209085 18241 209113
rect 18269 209085 18303 209113
rect 18331 209085 33477 209113
rect 33505 209085 33539 209113
rect 33567 209085 33601 209113
rect 33629 209085 33663 209113
rect 33691 209085 48837 209113
rect 48865 209085 48899 209113
rect 48927 209085 48961 209113
rect 48989 209085 49023 209113
rect 49051 209085 64197 209113
rect 64225 209085 64259 209113
rect 64287 209085 64321 209113
rect 64349 209085 64383 209113
rect 64411 209085 79557 209113
rect 79585 209085 79619 209113
rect 79647 209085 79681 209113
rect 79709 209085 79743 209113
rect 79771 209085 94917 209113
rect 94945 209085 94979 209113
rect 95007 209085 95041 209113
rect 95069 209085 95103 209113
rect 95131 209085 110277 209113
rect 110305 209085 110339 209113
rect 110367 209085 110401 209113
rect 110429 209085 110463 209113
rect 110491 209085 125637 209113
rect 125665 209085 125699 209113
rect 125727 209085 125761 209113
rect 125789 209085 125823 209113
rect 125851 209085 140997 209113
rect 141025 209085 141059 209113
rect 141087 209085 141121 209113
rect 141149 209085 141183 209113
rect 141211 209085 156357 209113
rect 156385 209085 156419 209113
rect 156447 209085 156481 209113
rect 156509 209085 156543 209113
rect 156571 209085 171717 209113
rect 171745 209085 171779 209113
rect 171807 209085 171841 209113
rect 171869 209085 171903 209113
rect 171931 209085 187077 209113
rect 187105 209085 187139 209113
rect 187167 209085 187201 209113
rect 187229 209085 187263 209113
rect 187291 209085 202437 209113
rect 202465 209085 202499 209113
rect 202527 209085 202561 209113
rect 202589 209085 202623 209113
rect 202651 209085 217797 209113
rect 217825 209085 217859 209113
rect 217887 209085 217921 209113
rect 217949 209085 217983 209113
rect 218011 209085 233157 209113
rect 233185 209085 233219 209113
rect 233247 209085 233281 209113
rect 233309 209085 233343 209113
rect 233371 209085 248517 209113
rect 248545 209085 248579 209113
rect 248607 209085 248641 209113
rect 248669 209085 248703 209113
rect 248731 209085 263877 209113
rect 263905 209085 263939 209113
rect 263967 209085 264001 209113
rect 264029 209085 264063 209113
rect 264091 209085 279237 209113
rect 279265 209085 279299 209113
rect 279327 209085 279361 209113
rect 279389 209085 279423 209113
rect 279451 209085 294597 209113
rect 294625 209085 294659 209113
rect 294687 209085 294721 209113
rect 294749 209085 294783 209113
rect 294811 209085 298248 209113
rect 298276 209085 298310 209113
rect 298338 209085 298372 209113
rect 298400 209085 298434 209113
rect 298462 209085 298990 209113
rect -958 209051 298990 209085
rect -958 209023 -430 209051
rect -402 209023 -368 209051
rect -340 209023 -306 209051
rect -278 209023 -244 209051
rect -216 209023 2757 209051
rect 2785 209023 2819 209051
rect 2847 209023 2881 209051
rect 2909 209023 2943 209051
rect 2971 209023 18117 209051
rect 18145 209023 18179 209051
rect 18207 209023 18241 209051
rect 18269 209023 18303 209051
rect 18331 209023 33477 209051
rect 33505 209023 33539 209051
rect 33567 209023 33601 209051
rect 33629 209023 33663 209051
rect 33691 209023 48837 209051
rect 48865 209023 48899 209051
rect 48927 209023 48961 209051
rect 48989 209023 49023 209051
rect 49051 209023 64197 209051
rect 64225 209023 64259 209051
rect 64287 209023 64321 209051
rect 64349 209023 64383 209051
rect 64411 209023 79557 209051
rect 79585 209023 79619 209051
rect 79647 209023 79681 209051
rect 79709 209023 79743 209051
rect 79771 209023 94917 209051
rect 94945 209023 94979 209051
rect 95007 209023 95041 209051
rect 95069 209023 95103 209051
rect 95131 209023 110277 209051
rect 110305 209023 110339 209051
rect 110367 209023 110401 209051
rect 110429 209023 110463 209051
rect 110491 209023 125637 209051
rect 125665 209023 125699 209051
rect 125727 209023 125761 209051
rect 125789 209023 125823 209051
rect 125851 209023 140997 209051
rect 141025 209023 141059 209051
rect 141087 209023 141121 209051
rect 141149 209023 141183 209051
rect 141211 209023 156357 209051
rect 156385 209023 156419 209051
rect 156447 209023 156481 209051
rect 156509 209023 156543 209051
rect 156571 209023 171717 209051
rect 171745 209023 171779 209051
rect 171807 209023 171841 209051
rect 171869 209023 171903 209051
rect 171931 209023 187077 209051
rect 187105 209023 187139 209051
rect 187167 209023 187201 209051
rect 187229 209023 187263 209051
rect 187291 209023 202437 209051
rect 202465 209023 202499 209051
rect 202527 209023 202561 209051
rect 202589 209023 202623 209051
rect 202651 209023 217797 209051
rect 217825 209023 217859 209051
rect 217887 209023 217921 209051
rect 217949 209023 217983 209051
rect 218011 209023 233157 209051
rect 233185 209023 233219 209051
rect 233247 209023 233281 209051
rect 233309 209023 233343 209051
rect 233371 209023 248517 209051
rect 248545 209023 248579 209051
rect 248607 209023 248641 209051
rect 248669 209023 248703 209051
rect 248731 209023 263877 209051
rect 263905 209023 263939 209051
rect 263967 209023 264001 209051
rect 264029 209023 264063 209051
rect 264091 209023 279237 209051
rect 279265 209023 279299 209051
rect 279327 209023 279361 209051
rect 279389 209023 279423 209051
rect 279451 209023 294597 209051
rect 294625 209023 294659 209051
rect 294687 209023 294721 209051
rect 294749 209023 294783 209051
rect 294811 209023 298248 209051
rect 298276 209023 298310 209051
rect 298338 209023 298372 209051
rect 298400 209023 298434 209051
rect 298462 209023 298990 209051
rect -958 208989 298990 209023
rect -958 208961 -430 208989
rect -402 208961 -368 208989
rect -340 208961 -306 208989
rect -278 208961 -244 208989
rect -216 208961 2757 208989
rect 2785 208961 2819 208989
rect 2847 208961 2881 208989
rect 2909 208961 2943 208989
rect 2971 208961 18117 208989
rect 18145 208961 18179 208989
rect 18207 208961 18241 208989
rect 18269 208961 18303 208989
rect 18331 208961 33477 208989
rect 33505 208961 33539 208989
rect 33567 208961 33601 208989
rect 33629 208961 33663 208989
rect 33691 208961 48837 208989
rect 48865 208961 48899 208989
rect 48927 208961 48961 208989
rect 48989 208961 49023 208989
rect 49051 208961 64197 208989
rect 64225 208961 64259 208989
rect 64287 208961 64321 208989
rect 64349 208961 64383 208989
rect 64411 208961 79557 208989
rect 79585 208961 79619 208989
rect 79647 208961 79681 208989
rect 79709 208961 79743 208989
rect 79771 208961 94917 208989
rect 94945 208961 94979 208989
rect 95007 208961 95041 208989
rect 95069 208961 95103 208989
rect 95131 208961 110277 208989
rect 110305 208961 110339 208989
rect 110367 208961 110401 208989
rect 110429 208961 110463 208989
rect 110491 208961 125637 208989
rect 125665 208961 125699 208989
rect 125727 208961 125761 208989
rect 125789 208961 125823 208989
rect 125851 208961 140997 208989
rect 141025 208961 141059 208989
rect 141087 208961 141121 208989
rect 141149 208961 141183 208989
rect 141211 208961 156357 208989
rect 156385 208961 156419 208989
rect 156447 208961 156481 208989
rect 156509 208961 156543 208989
rect 156571 208961 171717 208989
rect 171745 208961 171779 208989
rect 171807 208961 171841 208989
rect 171869 208961 171903 208989
rect 171931 208961 187077 208989
rect 187105 208961 187139 208989
rect 187167 208961 187201 208989
rect 187229 208961 187263 208989
rect 187291 208961 202437 208989
rect 202465 208961 202499 208989
rect 202527 208961 202561 208989
rect 202589 208961 202623 208989
rect 202651 208961 217797 208989
rect 217825 208961 217859 208989
rect 217887 208961 217921 208989
rect 217949 208961 217983 208989
rect 218011 208961 233157 208989
rect 233185 208961 233219 208989
rect 233247 208961 233281 208989
rect 233309 208961 233343 208989
rect 233371 208961 248517 208989
rect 248545 208961 248579 208989
rect 248607 208961 248641 208989
rect 248669 208961 248703 208989
rect 248731 208961 263877 208989
rect 263905 208961 263939 208989
rect 263967 208961 264001 208989
rect 264029 208961 264063 208989
rect 264091 208961 279237 208989
rect 279265 208961 279299 208989
rect 279327 208961 279361 208989
rect 279389 208961 279423 208989
rect 279451 208961 294597 208989
rect 294625 208961 294659 208989
rect 294687 208961 294721 208989
rect 294749 208961 294783 208989
rect 294811 208961 298248 208989
rect 298276 208961 298310 208989
rect 298338 208961 298372 208989
rect 298400 208961 298434 208989
rect 298462 208961 298990 208989
rect -958 208913 298990 208961
rect -958 203175 298990 203223
rect -958 203147 -910 203175
rect -882 203147 -848 203175
rect -820 203147 -786 203175
rect -758 203147 -724 203175
rect -696 203147 4617 203175
rect 4645 203147 4679 203175
rect 4707 203147 4741 203175
rect 4769 203147 4803 203175
rect 4831 203147 19977 203175
rect 20005 203147 20039 203175
rect 20067 203147 20101 203175
rect 20129 203147 20163 203175
rect 20191 203147 35337 203175
rect 35365 203147 35399 203175
rect 35427 203147 35461 203175
rect 35489 203147 35523 203175
rect 35551 203147 50697 203175
rect 50725 203147 50759 203175
rect 50787 203147 50821 203175
rect 50849 203147 50883 203175
rect 50911 203147 66057 203175
rect 66085 203147 66119 203175
rect 66147 203147 66181 203175
rect 66209 203147 66243 203175
rect 66271 203147 81417 203175
rect 81445 203147 81479 203175
rect 81507 203147 81541 203175
rect 81569 203147 81603 203175
rect 81631 203147 96777 203175
rect 96805 203147 96839 203175
rect 96867 203147 96901 203175
rect 96929 203147 96963 203175
rect 96991 203147 112137 203175
rect 112165 203147 112199 203175
rect 112227 203147 112261 203175
rect 112289 203147 112323 203175
rect 112351 203147 127497 203175
rect 127525 203147 127559 203175
rect 127587 203147 127621 203175
rect 127649 203147 127683 203175
rect 127711 203147 142857 203175
rect 142885 203147 142919 203175
rect 142947 203147 142981 203175
rect 143009 203147 143043 203175
rect 143071 203147 158217 203175
rect 158245 203147 158279 203175
rect 158307 203147 158341 203175
rect 158369 203147 158403 203175
rect 158431 203147 173577 203175
rect 173605 203147 173639 203175
rect 173667 203147 173701 203175
rect 173729 203147 173763 203175
rect 173791 203147 188937 203175
rect 188965 203147 188999 203175
rect 189027 203147 189061 203175
rect 189089 203147 189123 203175
rect 189151 203147 204297 203175
rect 204325 203147 204359 203175
rect 204387 203147 204421 203175
rect 204449 203147 204483 203175
rect 204511 203147 219657 203175
rect 219685 203147 219719 203175
rect 219747 203147 219781 203175
rect 219809 203147 219843 203175
rect 219871 203147 235017 203175
rect 235045 203147 235079 203175
rect 235107 203147 235141 203175
rect 235169 203147 235203 203175
rect 235231 203147 250377 203175
rect 250405 203147 250439 203175
rect 250467 203147 250501 203175
rect 250529 203147 250563 203175
rect 250591 203147 265737 203175
rect 265765 203147 265799 203175
rect 265827 203147 265861 203175
rect 265889 203147 265923 203175
rect 265951 203147 281097 203175
rect 281125 203147 281159 203175
rect 281187 203147 281221 203175
rect 281249 203147 281283 203175
rect 281311 203147 296457 203175
rect 296485 203147 296519 203175
rect 296547 203147 296581 203175
rect 296609 203147 296643 203175
rect 296671 203147 298728 203175
rect 298756 203147 298790 203175
rect 298818 203147 298852 203175
rect 298880 203147 298914 203175
rect 298942 203147 298990 203175
rect -958 203113 298990 203147
rect -958 203085 -910 203113
rect -882 203085 -848 203113
rect -820 203085 -786 203113
rect -758 203085 -724 203113
rect -696 203085 4617 203113
rect 4645 203085 4679 203113
rect 4707 203085 4741 203113
rect 4769 203085 4803 203113
rect 4831 203085 19977 203113
rect 20005 203085 20039 203113
rect 20067 203085 20101 203113
rect 20129 203085 20163 203113
rect 20191 203085 35337 203113
rect 35365 203085 35399 203113
rect 35427 203085 35461 203113
rect 35489 203085 35523 203113
rect 35551 203085 50697 203113
rect 50725 203085 50759 203113
rect 50787 203085 50821 203113
rect 50849 203085 50883 203113
rect 50911 203085 66057 203113
rect 66085 203085 66119 203113
rect 66147 203085 66181 203113
rect 66209 203085 66243 203113
rect 66271 203085 81417 203113
rect 81445 203085 81479 203113
rect 81507 203085 81541 203113
rect 81569 203085 81603 203113
rect 81631 203085 96777 203113
rect 96805 203085 96839 203113
rect 96867 203085 96901 203113
rect 96929 203085 96963 203113
rect 96991 203085 112137 203113
rect 112165 203085 112199 203113
rect 112227 203085 112261 203113
rect 112289 203085 112323 203113
rect 112351 203085 127497 203113
rect 127525 203085 127559 203113
rect 127587 203085 127621 203113
rect 127649 203085 127683 203113
rect 127711 203085 142857 203113
rect 142885 203085 142919 203113
rect 142947 203085 142981 203113
rect 143009 203085 143043 203113
rect 143071 203085 158217 203113
rect 158245 203085 158279 203113
rect 158307 203085 158341 203113
rect 158369 203085 158403 203113
rect 158431 203085 173577 203113
rect 173605 203085 173639 203113
rect 173667 203085 173701 203113
rect 173729 203085 173763 203113
rect 173791 203085 188937 203113
rect 188965 203085 188999 203113
rect 189027 203085 189061 203113
rect 189089 203085 189123 203113
rect 189151 203085 204297 203113
rect 204325 203085 204359 203113
rect 204387 203085 204421 203113
rect 204449 203085 204483 203113
rect 204511 203085 219657 203113
rect 219685 203085 219719 203113
rect 219747 203085 219781 203113
rect 219809 203085 219843 203113
rect 219871 203085 235017 203113
rect 235045 203085 235079 203113
rect 235107 203085 235141 203113
rect 235169 203085 235203 203113
rect 235231 203085 250377 203113
rect 250405 203085 250439 203113
rect 250467 203085 250501 203113
rect 250529 203085 250563 203113
rect 250591 203085 265737 203113
rect 265765 203085 265799 203113
rect 265827 203085 265861 203113
rect 265889 203085 265923 203113
rect 265951 203085 281097 203113
rect 281125 203085 281159 203113
rect 281187 203085 281221 203113
rect 281249 203085 281283 203113
rect 281311 203085 296457 203113
rect 296485 203085 296519 203113
rect 296547 203085 296581 203113
rect 296609 203085 296643 203113
rect 296671 203085 298728 203113
rect 298756 203085 298790 203113
rect 298818 203085 298852 203113
rect 298880 203085 298914 203113
rect 298942 203085 298990 203113
rect -958 203051 298990 203085
rect -958 203023 -910 203051
rect -882 203023 -848 203051
rect -820 203023 -786 203051
rect -758 203023 -724 203051
rect -696 203023 4617 203051
rect 4645 203023 4679 203051
rect 4707 203023 4741 203051
rect 4769 203023 4803 203051
rect 4831 203023 19977 203051
rect 20005 203023 20039 203051
rect 20067 203023 20101 203051
rect 20129 203023 20163 203051
rect 20191 203023 35337 203051
rect 35365 203023 35399 203051
rect 35427 203023 35461 203051
rect 35489 203023 35523 203051
rect 35551 203023 50697 203051
rect 50725 203023 50759 203051
rect 50787 203023 50821 203051
rect 50849 203023 50883 203051
rect 50911 203023 66057 203051
rect 66085 203023 66119 203051
rect 66147 203023 66181 203051
rect 66209 203023 66243 203051
rect 66271 203023 81417 203051
rect 81445 203023 81479 203051
rect 81507 203023 81541 203051
rect 81569 203023 81603 203051
rect 81631 203023 96777 203051
rect 96805 203023 96839 203051
rect 96867 203023 96901 203051
rect 96929 203023 96963 203051
rect 96991 203023 112137 203051
rect 112165 203023 112199 203051
rect 112227 203023 112261 203051
rect 112289 203023 112323 203051
rect 112351 203023 127497 203051
rect 127525 203023 127559 203051
rect 127587 203023 127621 203051
rect 127649 203023 127683 203051
rect 127711 203023 142857 203051
rect 142885 203023 142919 203051
rect 142947 203023 142981 203051
rect 143009 203023 143043 203051
rect 143071 203023 158217 203051
rect 158245 203023 158279 203051
rect 158307 203023 158341 203051
rect 158369 203023 158403 203051
rect 158431 203023 173577 203051
rect 173605 203023 173639 203051
rect 173667 203023 173701 203051
rect 173729 203023 173763 203051
rect 173791 203023 188937 203051
rect 188965 203023 188999 203051
rect 189027 203023 189061 203051
rect 189089 203023 189123 203051
rect 189151 203023 204297 203051
rect 204325 203023 204359 203051
rect 204387 203023 204421 203051
rect 204449 203023 204483 203051
rect 204511 203023 219657 203051
rect 219685 203023 219719 203051
rect 219747 203023 219781 203051
rect 219809 203023 219843 203051
rect 219871 203023 235017 203051
rect 235045 203023 235079 203051
rect 235107 203023 235141 203051
rect 235169 203023 235203 203051
rect 235231 203023 250377 203051
rect 250405 203023 250439 203051
rect 250467 203023 250501 203051
rect 250529 203023 250563 203051
rect 250591 203023 265737 203051
rect 265765 203023 265799 203051
rect 265827 203023 265861 203051
rect 265889 203023 265923 203051
rect 265951 203023 281097 203051
rect 281125 203023 281159 203051
rect 281187 203023 281221 203051
rect 281249 203023 281283 203051
rect 281311 203023 296457 203051
rect 296485 203023 296519 203051
rect 296547 203023 296581 203051
rect 296609 203023 296643 203051
rect 296671 203023 298728 203051
rect 298756 203023 298790 203051
rect 298818 203023 298852 203051
rect 298880 203023 298914 203051
rect 298942 203023 298990 203051
rect -958 202989 298990 203023
rect -958 202961 -910 202989
rect -882 202961 -848 202989
rect -820 202961 -786 202989
rect -758 202961 -724 202989
rect -696 202961 4617 202989
rect 4645 202961 4679 202989
rect 4707 202961 4741 202989
rect 4769 202961 4803 202989
rect 4831 202961 19977 202989
rect 20005 202961 20039 202989
rect 20067 202961 20101 202989
rect 20129 202961 20163 202989
rect 20191 202961 35337 202989
rect 35365 202961 35399 202989
rect 35427 202961 35461 202989
rect 35489 202961 35523 202989
rect 35551 202961 50697 202989
rect 50725 202961 50759 202989
rect 50787 202961 50821 202989
rect 50849 202961 50883 202989
rect 50911 202961 66057 202989
rect 66085 202961 66119 202989
rect 66147 202961 66181 202989
rect 66209 202961 66243 202989
rect 66271 202961 81417 202989
rect 81445 202961 81479 202989
rect 81507 202961 81541 202989
rect 81569 202961 81603 202989
rect 81631 202961 96777 202989
rect 96805 202961 96839 202989
rect 96867 202961 96901 202989
rect 96929 202961 96963 202989
rect 96991 202961 112137 202989
rect 112165 202961 112199 202989
rect 112227 202961 112261 202989
rect 112289 202961 112323 202989
rect 112351 202961 127497 202989
rect 127525 202961 127559 202989
rect 127587 202961 127621 202989
rect 127649 202961 127683 202989
rect 127711 202961 142857 202989
rect 142885 202961 142919 202989
rect 142947 202961 142981 202989
rect 143009 202961 143043 202989
rect 143071 202961 158217 202989
rect 158245 202961 158279 202989
rect 158307 202961 158341 202989
rect 158369 202961 158403 202989
rect 158431 202961 173577 202989
rect 173605 202961 173639 202989
rect 173667 202961 173701 202989
rect 173729 202961 173763 202989
rect 173791 202961 188937 202989
rect 188965 202961 188999 202989
rect 189027 202961 189061 202989
rect 189089 202961 189123 202989
rect 189151 202961 204297 202989
rect 204325 202961 204359 202989
rect 204387 202961 204421 202989
rect 204449 202961 204483 202989
rect 204511 202961 219657 202989
rect 219685 202961 219719 202989
rect 219747 202961 219781 202989
rect 219809 202961 219843 202989
rect 219871 202961 235017 202989
rect 235045 202961 235079 202989
rect 235107 202961 235141 202989
rect 235169 202961 235203 202989
rect 235231 202961 250377 202989
rect 250405 202961 250439 202989
rect 250467 202961 250501 202989
rect 250529 202961 250563 202989
rect 250591 202961 265737 202989
rect 265765 202961 265799 202989
rect 265827 202961 265861 202989
rect 265889 202961 265923 202989
rect 265951 202961 281097 202989
rect 281125 202961 281159 202989
rect 281187 202961 281221 202989
rect 281249 202961 281283 202989
rect 281311 202961 296457 202989
rect 296485 202961 296519 202989
rect 296547 202961 296581 202989
rect 296609 202961 296643 202989
rect 296671 202961 298728 202989
rect 298756 202961 298790 202989
rect 298818 202961 298852 202989
rect 298880 202961 298914 202989
rect 298942 202961 298990 202989
rect -958 202913 298990 202961
rect -958 200175 298990 200223
rect -958 200147 -430 200175
rect -402 200147 -368 200175
rect -340 200147 -306 200175
rect -278 200147 -244 200175
rect -216 200147 2757 200175
rect 2785 200147 2819 200175
rect 2847 200147 2881 200175
rect 2909 200147 2943 200175
rect 2971 200147 18117 200175
rect 18145 200147 18179 200175
rect 18207 200147 18241 200175
rect 18269 200147 18303 200175
rect 18331 200147 33477 200175
rect 33505 200147 33539 200175
rect 33567 200147 33601 200175
rect 33629 200147 33663 200175
rect 33691 200147 48837 200175
rect 48865 200147 48899 200175
rect 48927 200147 48961 200175
rect 48989 200147 49023 200175
rect 49051 200147 64197 200175
rect 64225 200147 64259 200175
rect 64287 200147 64321 200175
rect 64349 200147 64383 200175
rect 64411 200147 79557 200175
rect 79585 200147 79619 200175
rect 79647 200147 79681 200175
rect 79709 200147 79743 200175
rect 79771 200147 94917 200175
rect 94945 200147 94979 200175
rect 95007 200147 95041 200175
rect 95069 200147 95103 200175
rect 95131 200147 110277 200175
rect 110305 200147 110339 200175
rect 110367 200147 110401 200175
rect 110429 200147 110463 200175
rect 110491 200147 125637 200175
rect 125665 200147 125699 200175
rect 125727 200147 125761 200175
rect 125789 200147 125823 200175
rect 125851 200147 140997 200175
rect 141025 200147 141059 200175
rect 141087 200147 141121 200175
rect 141149 200147 141183 200175
rect 141211 200147 156357 200175
rect 156385 200147 156419 200175
rect 156447 200147 156481 200175
rect 156509 200147 156543 200175
rect 156571 200147 171717 200175
rect 171745 200147 171779 200175
rect 171807 200147 171841 200175
rect 171869 200147 171903 200175
rect 171931 200147 187077 200175
rect 187105 200147 187139 200175
rect 187167 200147 187201 200175
rect 187229 200147 187263 200175
rect 187291 200147 202437 200175
rect 202465 200147 202499 200175
rect 202527 200147 202561 200175
rect 202589 200147 202623 200175
rect 202651 200147 217797 200175
rect 217825 200147 217859 200175
rect 217887 200147 217921 200175
rect 217949 200147 217983 200175
rect 218011 200147 233157 200175
rect 233185 200147 233219 200175
rect 233247 200147 233281 200175
rect 233309 200147 233343 200175
rect 233371 200147 248517 200175
rect 248545 200147 248579 200175
rect 248607 200147 248641 200175
rect 248669 200147 248703 200175
rect 248731 200147 263877 200175
rect 263905 200147 263939 200175
rect 263967 200147 264001 200175
rect 264029 200147 264063 200175
rect 264091 200147 279237 200175
rect 279265 200147 279299 200175
rect 279327 200147 279361 200175
rect 279389 200147 279423 200175
rect 279451 200147 294597 200175
rect 294625 200147 294659 200175
rect 294687 200147 294721 200175
rect 294749 200147 294783 200175
rect 294811 200147 298248 200175
rect 298276 200147 298310 200175
rect 298338 200147 298372 200175
rect 298400 200147 298434 200175
rect 298462 200147 298990 200175
rect -958 200113 298990 200147
rect -958 200085 -430 200113
rect -402 200085 -368 200113
rect -340 200085 -306 200113
rect -278 200085 -244 200113
rect -216 200085 2757 200113
rect 2785 200085 2819 200113
rect 2847 200085 2881 200113
rect 2909 200085 2943 200113
rect 2971 200085 18117 200113
rect 18145 200085 18179 200113
rect 18207 200085 18241 200113
rect 18269 200085 18303 200113
rect 18331 200085 33477 200113
rect 33505 200085 33539 200113
rect 33567 200085 33601 200113
rect 33629 200085 33663 200113
rect 33691 200085 48837 200113
rect 48865 200085 48899 200113
rect 48927 200085 48961 200113
rect 48989 200085 49023 200113
rect 49051 200085 64197 200113
rect 64225 200085 64259 200113
rect 64287 200085 64321 200113
rect 64349 200085 64383 200113
rect 64411 200085 79557 200113
rect 79585 200085 79619 200113
rect 79647 200085 79681 200113
rect 79709 200085 79743 200113
rect 79771 200085 94917 200113
rect 94945 200085 94979 200113
rect 95007 200085 95041 200113
rect 95069 200085 95103 200113
rect 95131 200085 110277 200113
rect 110305 200085 110339 200113
rect 110367 200085 110401 200113
rect 110429 200085 110463 200113
rect 110491 200085 125637 200113
rect 125665 200085 125699 200113
rect 125727 200085 125761 200113
rect 125789 200085 125823 200113
rect 125851 200085 140997 200113
rect 141025 200085 141059 200113
rect 141087 200085 141121 200113
rect 141149 200085 141183 200113
rect 141211 200085 156357 200113
rect 156385 200085 156419 200113
rect 156447 200085 156481 200113
rect 156509 200085 156543 200113
rect 156571 200085 171717 200113
rect 171745 200085 171779 200113
rect 171807 200085 171841 200113
rect 171869 200085 171903 200113
rect 171931 200085 187077 200113
rect 187105 200085 187139 200113
rect 187167 200085 187201 200113
rect 187229 200085 187263 200113
rect 187291 200085 202437 200113
rect 202465 200085 202499 200113
rect 202527 200085 202561 200113
rect 202589 200085 202623 200113
rect 202651 200085 217797 200113
rect 217825 200085 217859 200113
rect 217887 200085 217921 200113
rect 217949 200085 217983 200113
rect 218011 200085 233157 200113
rect 233185 200085 233219 200113
rect 233247 200085 233281 200113
rect 233309 200085 233343 200113
rect 233371 200085 248517 200113
rect 248545 200085 248579 200113
rect 248607 200085 248641 200113
rect 248669 200085 248703 200113
rect 248731 200085 263877 200113
rect 263905 200085 263939 200113
rect 263967 200085 264001 200113
rect 264029 200085 264063 200113
rect 264091 200085 279237 200113
rect 279265 200085 279299 200113
rect 279327 200085 279361 200113
rect 279389 200085 279423 200113
rect 279451 200085 294597 200113
rect 294625 200085 294659 200113
rect 294687 200085 294721 200113
rect 294749 200085 294783 200113
rect 294811 200085 298248 200113
rect 298276 200085 298310 200113
rect 298338 200085 298372 200113
rect 298400 200085 298434 200113
rect 298462 200085 298990 200113
rect -958 200051 298990 200085
rect -958 200023 -430 200051
rect -402 200023 -368 200051
rect -340 200023 -306 200051
rect -278 200023 -244 200051
rect -216 200023 2757 200051
rect 2785 200023 2819 200051
rect 2847 200023 2881 200051
rect 2909 200023 2943 200051
rect 2971 200023 18117 200051
rect 18145 200023 18179 200051
rect 18207 200023 18241 200051
rect 18269 200023 18303 200051
rect 18331 200023 33477 200051
rect 33505 200023 33539 200051
rect 33567 200023 33601 200051
rect 33629 200023 33663 200051
rect 33691 200023 48837 200051
rect 48865 200023 48899 200051
rect 48927 200023 48961 200051
rect 48989 200023 49023 200051
rect 49051 200023 64197 200051
rect 64225 200023 64259 200051
rect 64287 200023 64321 200051
rect 64349 200023 64383 200051
rect 64411 200023 79557 200051
rect 79585 200023 79619 200051
rect 79647 200023 79681 200051
rect 79709 200023 79743 200051
rect 79771 200023 94917 200051
rect 94945 200023 94979 200051
rect 95007 200023 95041 200051
rect 95069 200023 95103 200051
rect 95131 200023 110277 200051
rect 110305 200023 110339 200051
rect 110367 200023 110401 200051
rect 110429 200023 110463 200051
rect 110491 200023 125637 200051
rect 125665 200023 125699 200051
rect 125727 200023 125761 200051
rect 125789 200023 125823 200051
rect 125851 200023 140997 200051
rect 141025 200023 141059 200051
rect 141087 200023 141121 200051
rect 141149 200023 141183 200051
rect 141211 200023 156357 200051
rect 156385 200023 156419 200051
rect 156447 200023 156481 200051
rect 156509 200023 156543 200051
rect 156571 200023 171717 200051
rect 171745 200023 171779 200051
rect 171807 200023 171841 200051
rect 171869 200023 171903 200051
rect 171931 200023 187077 200051
rect 187105 200023 187139 200051
rect 187167 200023 187201 200051
rect 187229 200023 187263 200051
rect 187291 200023 202437 200051
rect 202465 200023 202499 200051
rect 202527 200023 202561 200051
rect 202589 200023 202623 200051
rect 202651 200023 217797 200051
rect 217825 200023 217859 200051
rect 217887 200023 217921 200051
rect 217949 200023 217983 200051
rect 218011 200023 233157 200051
rect 233185 200023 233219 200051
rect 233247 200023 233281 200051
rect 233309 200023 233343 200051
rect 233371 200023 248517 200051
rect 248545 200023 248579 200051
rect 248607 200023 248641 200051
rect 248669 200023 248703 200051
rect 248731 200023 263877 200051
rect 263905 200023 263939 200051
rect 263967 200023 264001 200051
rect 264029 200023 264063 200051
rect 264091 200023 279237 200051
rect 279265 200023 279299 200051
rect 279327 200023 279361 200051
rect 279389 200023 279423 200051
rect 279451 200023 294597 200051
rect 294625 200023 294659 200051
rect 294687 200023 294721 200051
rect 294749 200023 294783 200051
rect 294811 200023 298248 200051
rect 298276 200023 298310 200051
rect 298338 200023 298372 200051
rect 298400 200023 298434 200051
rect 298462 200023 298990 200051
rect -958 199989 298990 200023
rect -958 199961 -430 199989
rect -402 199961 -368 199989
rect -340 199961 -306 199989
rect -278 199961 -244 199989
rect -216 199961 2757 199989
rect 2785 199961 2819 199989
rect 2847 199961 2881 199989
rect 2909 199961 2943 199989
rect 2971 199961 18117 199989
rect 18145 199961 18179 199989
rect 18207 199961 18241 199989
rect 18269 199961 18303 199989
rect 18331 199961 33477 199989
rect 33505 199961 33539 199989
rect 33567 199961 33601 199989
rect 33629 199961 33663 199989
rect 33691 199961 48837 199989
rect 48865 199961 48899 199989
rect 48927 199961 48961 199989
rect 48989 199961 49023 199989
rect 49051 199961 64197 199989
rect 64225 199961 64259 199989
rect 64287 199961 64321 199989
rect 64349 199961 64383 199989
rect 64411 199961 79557 199989
rect 79585 199961 79619 199989
rect 79647 199961 79681 199989
rect 79709 199961 79743 199989
rect 79771 199961 94917 199989
rect 94945 199961 94979 199989
rect 95007 199961 95041 199989
rect 95069 199961 95103 199989
rect 95131 199961 110277 199989
rect 110305 199961 110339 199989
rect 110367 199961 110401 199989
rect 110429 199961 110463 199989
rect 110491 199961 125637 199989
rect 125665 199961 125699 199989
rect 125727 199961 125761 199989
rect 125789 199961 125823 199989
rect 125851 199961 140997 199989
rect 141025 199961 141059 199989
rect 141087 199961 141121 199989
rect 141149 199961 141183 199989
rect 141211 199961 156357 199989
rect 156385 199961 156419 199989
rect 156447 199961 156481 199989
rect 156509 199961 156543 199989
rect 156571 199961 171717 199989
rect 171745 199961 171779 199989
rect 171807 199961 171841 199989
rect 171869 199961 171903 199989
rect 171931 199961 187077 199989
rect 187105 199961 187139 199989
rect 187167 199961 187201 199989
rect 187229 199961 187263 199989
rect 187291 199961 202437 199989
rect 202465 199961 202499 199989
rect 202527 199961 202561 199989
rect 202589 199961 202623 199989
rect 202651 199961 217797 199989
rect 217825 199961 217859 199989
rect 217887 199961 217921 199989
rect 217949 199961 217983 199989
rect 218011 199961 233157 199989
rect 233185 199961 233219 199989
rect 233247 199961 233281 199989
rect 233309 199961 233343 199989
rect 233371 199961 248517 199989
rect 248545 199961 248579 199989
rect 248607 199961 248641 199989
rect 248669 199961 248703 199989
rect 248731 199961 263877 199989
rect 263905 199961 263939 199989
rect 263967 199961 264001 199989
rect 264029 199961 264063 199989
rect 264091 199961 279237 199989
rect 279265 199961 279299 199989
rect 279327 199961 279361 199989
rect 279389 199961 279423 199989
rect 279451 199961 294597 199989
rect 294625 199961 294659 199989
rect 294687 199961 294721 199989
rect 294749 199961 294783 199989
rect 294811 199961 298248 199989
rect 298276 199961 298310 199989
rect 298338 199961 298372 199989
rect 298400 199961 298434 199989
rect 298462 199961 298990 199989
rect -958 199913 298990 199961
rect -958 194175 298990 194223
rect -958 194147 -910 194175
rect -882 194147 -848 194175
rect -820 194147 -786 194175
rect -758 194147 -724 194175
rect -696 194147 4617 194175
rect 4645 194147 4679 194175
rect 4707 194147 4741 194175
rect 4769 194147 4803 194175
rect 4831 194147 19977 194175
rect 20005 194147 20039 194175
rect 20067 194147 20101 194175
rect 20129 194147 20163 194175
rect 20191 194147 35337 194175
rect 35365 194147 35399 194175
rect 35427 194147 35461 194175
rect 35489 194147 35523 194175
rect 35551 194147 50697 194175
rect 50725 194147 50759 194175
rect 50787 194147 50821 194175
rect 50849 194147 50883 194175
rect 50911 194147 66057 194175
rect 66085 194147 66119 194175
rect 66147 194147 66181 194175
rect 66209 194147 66243 194175
rect 66271 194147 81417 194175
rect 81445 194147 81479 194175
rect 81507 194147 81541 194175
rect 81569 194147 81603 194175
rect 81631 194147 96777 194175
rect 96805 194147 96839 194175
rect 96867 194147 96901 194175
rect 96929 194147 96963 194175
rect 96991 194147 112137 194175
rect 112165 194147 112199 194175
rect 112227 194147 112261 194175
rect 112289 194147 112323 194175
rect 112351 194147 127497 194175
rect 127525 194147 127559 194175
rect 127587 194147 127621 194175
rect 127649 194147 127683 194175
rect 127711 194147 142857 194175
rect 142885 194147 142919 194175
rect 142947 194147 142981 194175
rect 143009 194147 143043 194175
rect 143071 194147 158217 194175
rect 158245 194147 158279 194175
rect 158307 194147 158341 194175
rect 158369 194147 158403 194175
rect 158431 194147 173577 194175
rect 173605 194147 173639 194175
rect 173667 194147 173701 194175
rect 173729 194147 173763 194175
rect 173791 194147 188937 194175
rect 188965 194147 188999 194175
rect 189027 194147 189061 194175
rect 189089 194147 189123 194175
rect 189151 194147 204297 194175
rect 204325 194147 204359 194175
rect 204387 194147 204421 194175
rect 204449 194147 204483 194175
rect 204511 194147 219657 194175
rect 219685 194147 219719 194175
rect 219747 194147 219781 194175
rect 219809 194147 219843 194175
rect 219871 194147 235017 194175
rect 235045 194147 235079 194175
rect 235107 194147 235141 194175
rect 235169 194147 235203 194175
rect 235231 194147 250377 194175
rect 250405 194147 250439 194175
rect 250467 194147 250501 194175
rect 250529 194147 250563 194175
rect 250591 194147 265737 194175
rect 265765 194147 265799 194175
rect 265827 194147 265861 194175
rect 265889 194147 265923 194175
rect 265951 194147 281097 194175
rect 281125 194147 281159 194175
rect 281187 194147 281221 194175
rect 281249 194147 281283 194175
rect 281311 194147 296457 194175
rect 296485 194147 296519 194175
rect 296547 194147 296581 194175
rect 296609 194147 296643 194175
rect 296671 194147 298728 194175
rect 298756 194147 298790 194175
rect 298818 194147 298852 194175
rect 298880 194147 298914 194175
rect 298942 194147 298990 194175
rect -958 194113 298990 194147
rect -958 194085 -910 194113
rect -882 194085 -848 194113
rect -820 194085 -786 194113
rect -758 194085 -724 194113
rect -696 194085 4617 194113
rect 4645 194085 4679 194113
rect 4707 194085 4741 194113
rect 4769 194085 4803 194113
rect 4831 194085 19977 194113
rect 20005 194085 20039 194113
rect 20067 194085 20101 194113
rect 20129 194085 20163 194113
rect 20191 194085 35337 194113
rect 35365 194085 35399 194113
rect 35427 194085 35461 194113
rect 35489 194085 35523 194113
rect 35551 194085 50697 194113
rect 50725 194085 50759 194113
rect 50787 194085 50821 194113
rect 50849 194085 50883 194113
rect 50911 194085 66057 194113
rect 66085 194085 66119 194113
rect 66147 194085 66181 194113
rect 66209 194085 66243 194113
rect 66271 194085 81417 194113
rect 81445 194085 81479 194113
rect 81507 194085 81541 194113
rect 81569 194085 81603 194113
rect 81631 194085 96777 194113
rect 96805 194085 96839 194113
rect 96867 194085 96901 194113
rect 96929 194085 96963 194113
rect 96991 194085 112137 194113
rect 112165 194085 112199 194113
rect 112227 194085 112261 194113
rect 112289 194085 112323 194113
rect 112351 194085 127497 194113
rect 127525 194085 127559 194113
rect 127587 194085 127621 194113
rect 127649 194085 127683 194113
rect 127711 194085 142857 194113
rect 142885 194085 142919 194113
rect 142947 194085 142981 194113
rect 143009 194085 143043 194113
rect 143071 194085 158217 194113
rect 158245 194085 158279 194113
rect 158307 194085 158341 194113
rect 158369 194085 158403 194113
rect 158431 194085 173577 194113
rect 173605 194085 173639 194113
rect 173667 194085 173701 194113
rect 173729 194085 173763 194113
rect 173791 194085 188937 194113
rect 188965 194085 188999 194113
rect 189027 194085 189061 194113
rect 189089 194085 189123 194113
rect 189151 194085 204297 194113
rect 204325 194085 204359 194113
rect 204387 194085 204421 194113
rect 204449 194085 204483 194113
rect 204511 194085 219657 194113
rect 219685 194085 219719 194113
rect 219747 194085 219781 194113
rect 219809 194085 219843 194113
rect 219871 194085 235017 194113
rect 235045 194085 235079 194113
rect 235107 194085 235141 194113
rect 235169 194085 235203 194113
rect 235231 194085 250377 194113
rect 250405 194085 250439 194113
rect 250467 194085 250501 194113
rect 250529 194085 250563 194113
rect 250591 194085 265737 194113
rect 265765 194085 265799 194113
rect 265827 194085 265861 194113
rect 265889 194085 265923 194113
rect 265951 194085 281097 194113
rect 281125 194085 281159 194113
rect 281187 194085 281221 194113
rect 281249 194085 281283 194113
rect 281311 194085 296457 194113
rect 296485 194085 296519 194113
rect 296547 194085 296581 194113
rect 296609 194085 296643 194113
rect 296671 194085 298728 194113
rect 298756 194085 298790 194113
rect 298818 194085 298852 194113
rect 298880 194085 298914 194113
rect 298942 194085 298990 194113
rect -958 194051 298990 194085
rect -958 194023 -910 194051
rect -882 194023 -848 194051
rect -820 194023 -786 194051
rect -758 194023 -724 194051
rect -696 194023 4617 194051
rect 4645 194023 4679 194051
rect 4707 194023 4741 194051
rect 4769 194023 4803 194051
rect 4831 194023 19977 194051
rect 20005 194023 20039 194051
rect 20067 194023 20101 194051
rect 20129 194023 20163 194051
rect 20191 194023 35337 194051
rect 35365 194023 35399 194051
rect 35427 194023 35461 194051
rect 35489 194023 35523 194051
rect 35551 194023 50697 194051
rect 50725 194023 50759 194051
rect 50787 194023 50821 194051
rect 50849 194023 50883 194051
rect 50911 194023 66057 194051
rect 66085 194023 66119 194051
rect 66147 194023 66181 194051
rect 66209 194023 66243 194051
rect 66271 194023 81417 194051
rect 81445 194023 81479 194051
rect 81507 194023 81541 194051
rect 81569 194023 81603 194051
rect 81631 194023 96777 194051
rect 96805 194023 96839 194051
rect 96867 194023 96901 194051
rect 96929 194023 96963 194051
rect 96991 194023 112137 194051
rect 112165 194023 112199 194051
rect 112227 194023 112261 194051
rect 112289 194023 112323 194051
rect 112351 194023 127497 194051
rect 127525 194023 127559 194051
rect 127587 194023 127621 194051
rect 127649 194023 127683 194051
rect 127711 194023 142857 194051
rect 142885 194023 142919 194051
rect 142947 194023 142981 194051
rect 143009 194023 143043 194051
rect 143071 194023 158217 194051
rect 158245 194023 158279 194051
rect 158307 194023 158341 194051
rect 158369 194023 158403 194051
rect 158431 194023 173577 194051
rect 173605 194023 173639 194051
rect 173667 194023 173701 194051
rect 173729 194023 173763 194051
rect 173791 194023 188937 194051
rect 188965 194023 188999 194051
rect 189027 194023 189061 194051
rect 189089 194023 189123 194051
rect 189151 194023 204297 194051
rect 204325 194023 204359 194051
rect 204387 194023 204421 194051
rect 204449 194023 204483 194051
rect 204511 194023 219657 194051
rect 219685 194023 219719 194051
rect 219747 194023 219781 194051
rect 219809 194023 219843 194051
rect 219871 194023 235017 194051
rect 235045 194023 235079 194051
rect 235107 194023 235141 194051
rect 235169 194023 235203 194051
rect 235231 194023 250377 194051
rect 250405 194023 250439 194051
rect 250467 194023 250501 194051
rect 250529 194023 250563 194051
rect 250591 194023 265737 194051
rect 265765 194023 265799 194051
rect 265827 194023 265861 194051
rect 265889 194023 265923 194051
rect 265951 194023 281097 194051
rect 281125 194023 281159 194051
rect 281187 194023 281221 194051
rect 281249 194023 281283 194051
rect 281311 194023 296457 194051
rect 296485 194023 296519 194051
rect 296547 194023 296581 194051
rect 296609 194023 296643 194051
rect 296671 194023 298728 194051
rect 298756 194023 298790 194051
rect 298818 194023 298852 194051
rect 298880 194023 298914 194051
rect 298942 194023 298990 194051
rect -958 193989 298990 194023
rect -958 193961 -910 193989
rect -882 193961 -848 193989
rect -820 193961 -786 193989
rect -758 193961 -724 193989
rect -696 193961 4617 193989
rect 4645 193961 4679 193989
rect 4707 193961 4741 193989
rect 4769 193961 4803 193989
rect 4831 193961 19977 193989
rect 20005 193961 20039 193989
rect 20067 193961 20101 193989
rect 20129 193961 20163 193989
rect 20191 193961 35337 193989
rect 35365 193961 35399 193989
rect 35427 193961 35461 193989
rect 35489 193961 35523 193989
rect 35551 193961 50697 193989
rect 50725 193961 50759 193989
rect 50787 193961 50821 193989
rect 50849 193961 50883 193989
rect 50911 193961 66057 193989
rect 66085 193961 66119 193989
rect 66147 193961 66181 193989
rect 66209 193961 66243 193989
rect 66271 193961 81417 193989
rect 81445 193961 81479 193989
rect 81507 193961 81541 193989
rect 81569 193961 81603 193989
rect 81631 193961 96777 193989
rect 96805 193961 96839 193989
rect 96867 193961 96901 193989
rect 96929 193961 96963 193989
rect 96991 193961 112137 193989
rect 112165 193961 112199 193989
rect 112227 193961 112261 193989
rect 112289 193961 112323 193989
rect 112351 193961 127497 193989
rect 127525 193961 127559 193989
rect 127587 193961 127621 193989
rect 127649 193961 127683 193989
rect 127711 193961 142857 193989
rect 142885 193961 142919 193989
rect 142947 193961 142981 193989
rect 143009 193961 143043 193989
rect 143071 193961 158217 193989
rect 158245 193961 158279 193989
rect 158307 193961 158341 193989
rect 158369 193961 158403 193989
rect 158431 193961 173577 193989
rect 173605 193961 173639 193989
rect 173667 193961 173701 193989
rect 173729 193961 173763 193989
rect 173791 193961 188937 193989
rect 188965 193961 188999 193989
rect 189027 193961 189061 193989
rect 189089 193961 189123 193989
rect 189151 193961 204297 193989
rect 204325 193961 204359 193989
rect 204387 193961 204421 193989
rect 204449 193961 204483 193989
rect 204511 193961 219657 193989
rect 219685 193961 219719 193989
rect 219747 193961 219781 193989
rect 219809 193961 219843 193989
rect 219871 193961 235017 193989
rect 235045 193961 235079 193989
rect 235107 193961 235141 193989
rect 235169 193961 235203 193989
rect 235231 193961 250377 193989
rect 250405 193961 250439 193989
rect 250467 193961 250501 193989
rect 250529 193961 250563 193989
rect 250591 193961 265737 193989
rect 265765 193961 265799 193989
rect 265827 193961 265861 193989
rect 265889 193961 265923 193989
rect 265951 193961 281097 193989
rect 281125 193961 281159 193989
rect 281187 193961 281221 193989
rect 281249 193961 281283 193989
rect 281311 193961 296457 193989
rect 296485 193961 296519 193989
rect 296547 193961 296581 193989
rect 296609 193961 296643 193989
rect 296671 193961 298728 193989
rect 298756 193961 298790 193989
rect 298818 193961 298852 193989
rect 298880 193961 298914 193989
rect 298942 193961 298990 193989
rect -958 193913 298990 193961
rect -958 191175 298990 191223
rect -958 191147 -430 191175
rect -402 191147 -368 191175
rect -340 191147 -306 191175
rect -278 191147 -244 191175
rect -216 191147 2757 191175
rect 2785 191147 2819 191175
rect 2847 191147 2881 191175
rect 2909 191147 2943 191175
rect 2971 191147 18117 191175
rect 18145 191147 18179 191175
rect 18207 191147 18241 191175
rect 18269 191147 18303 191175
rect 18331 191147 33477 191175
rect 33505 191147 33539 191175
rect 33567 191147 33601 191175
rect 33629 191147 33663 191175
rect 33691 191147 48837 191175
rect 48865 191147 48899 191175
rect 48927 191147 48961 191175
rect 48989 191147 49023 191175
rect 49051 191147 64197 191175
rect 64225 191147 64259 191175
rect 64287 191147 64321 191175
rect 64349 191147 64383 191175
rect 64411 191147 79557 191175
rect 79585 191147 79619 191175
rect 79647 191147 79681 191175
rect 79709 191147 79743 191175
rect 79771 191147 94917 191175
rect 94945 191147 94979 191175
rect 95007 191147 95041 191175
rect 95069 191147 95103 191175
rect 95131 191147 110277 191175
rect 110305 191147 110339 191175
rect 110367 191147 110401 191175
rect 110429 191147 110463 191175
rect 110491 191147 125637 191175
rect 125665 191147 125699 191175
rect 125727 191147 125761 191175
rect 125789 191147 125823 191175
rect 125851 191147 140997 191175
rect 141025 191147 141059 191175
rect 141087 191147 141121 191175
rect 141149 191147 141183 191175
rect 141211 191147 156357 191175
rect 156385 191147 156419 191175
rect 156447 191147 156481 191175
rect 156509 191147 156543 191175
rect 156571 191147 171717 191175
rect 171745 191147 171779 191175
rect 171807 191147 171841 191175
rect 171869 191147 171903 191175
rect 171931 191147 187077 191175
rect 187105 191147 187139 191175
rect 187167 191147 187201 191175
rect 187229 191147 187263 191175
rect 187291 191147 202437 191175
rect 202465 191147 202499 191175
rect 202527 191147 202561 191175
rect 202589 191147 202623 191175
rect 202651 191147 217797 191175
rect 217825 191147 217859 191175
rect 217887 191147 217921 191175
rect 217949 191147 217983 191175
rect 218011 191147 233157 191175
rect 233185 191147 233219 191175
rect 233247 191147 233281 191175
rect 233309 191147 233343 191175
rect 233371 191147 248517 191175
rect 248545 191147 248579 191175
rect 248607 191147 248641 191175
rect 248669 191147 248703 191175
rect 248731 191147 263877 191175
rect 263905 191147 263939 191175
rect 263967 191147 264001 191175
rect 264029 191147 264063 191175
rect 264091 191147 279237 191175
rect 279265 191147 279299 191175
rect 279327 191147 279361 191175
rect 279389 191147 279423 191175
rect 279451 191147 294597 191175
rect 294625 191147 294659 191175
rect 294687 191147 294721 191175
rect 294749 191147 294783 191175
rect 294811 191147 298248 191175
rect 298276 191147 298310 191175
rect 298338 191147 298372 191175
rect 298400 191147 298434 191175
rect 298462 191147 298990 191175
rect -958 191113 298990 191147
rect -958 191085 -430 191113
rect -402 191085 -368 191113
rect -340 191085 -306 191113
rect -278 191085 -244 191113
rect -216 191085 2757 191113
rect 2785 191085 2819 191113
rect 2847 191085 2881 191113
rect 2909 191085 2943 191113
rect 2971 191085 18117 191113
rect 18145 191085 18179 191113
rect 18207 191085 18241 191113
rect 18269 191085 18303 191113
rect 18331 191085 33477 191113
rect 33505 191085 33539 191113
rect 33567 191085 33601 191113
rect 33629 191085 33663 191113
rect 33691 191085 48837 191113
rect 48865 191085 48899 191113
rect 48927 191085 48961 191113
rect 48989 191085 49023 191113
rect 49051 191085 64197 191113
rect 64225 191085 64259 191113
rect 64287 191085 64321 191113
rect 64349 191085 64383 191113
rect 64411 191085 79557 191113
rect 79585 191085 79619 191113
rect 79647 191085 79681 191113
rect 79709 191085 79743 191113
rect 79771 191085 94917 191113
rect 94945 191085 94979 191113
rect 95007 191085 95041 191113
rect 95069 191085 95103 191113
rect 95131 191085 110277 191113
rect 110305 191085 110339 191113
rect 110367 191085 110401 191113
rect 110429 191085 110463 191113
rect 110491 191085 125637 191113
rect 125665 191085 125699 191113
rect 125727 191085 125761 191113
rect 125789 191085 125823 191113
rect 125851 191085 140997 191113
rect 141025 191085 141059 191113
rect 141087 191085 141121 191113
rect 141149 191085 141183 191113
rect 141211 191085 156357 191113
rect 156385 191085 156419 191113
rect 156447 191085 156481 191113
rect 156509 191085 156543 191113
rect 156571 191085 171717 191113
rect 171745 191085 171779 191113
rect 171807 191085 171841 191113
rect 171869 191085 171903 191113
rect 171931 191085 187077 191113
rect 187105 191085 187139 191113
rect 187167 191085 187201 191113
rect 187229 191085 187263 191113
rect 187291 191085 202437 191113
rect 202465 191085 202499 191113
rect 202527 191085 202561 191113
rect 202589 191085 202623 191113
rect 202651 191085 217797 191113
rect 217825 191085 217859 191113
rect 217887 191085 217921 191113
rect 217949 191085 217983 191113
rect 218011 191085 233157 191113
rect 233185 191085 233219 191113
rect 233247 191085 233281 191113
rect 233309 191085 233343 191113
rect 233371 191085 248517 191113
rect 248545 191085 248579 191113
rect 248607 191085 248641 191113
rect 248669 191085 248703 191113
rect 248731 191085 263877 191113
rect 263905 191085 263939 191113
rect 263967 191085 264001 191113
rect 264029 191085 264063 191113
rect 264091 191085 279237 191113
rect 279265 191085 279299 191113
rect 279327 191085 279361 191113
rect 279389 191085 279423 191113
rect 279451 191085 294597 191113
rect 294625 191085 294659 191113
rect 294687 191085 294721 191113
rect 294749 191085 294783 191113
rect 294811 191085 298248 191113
rect 298276 191085 298310 191113
rect 298338 191085 298372 191113
rect 298400 191085 298434 191113
rect 298462 191085 298990 191113
rect -958 191051 298990 191085
rect -958 191023 -430 191051
rect -402 191023 -368 191051
rect -340 191023 -306 191051
rect -278 191023 -244 191051
rect -216 191023 2757 191051
rect 2785 191023 2819 191051
rect 2847 191023 2881 191051
rect 2909 191023 2943 191051
rect 2971 191023 18117 191051
rect 18145 191023 18179 191051
rect 18207 191023 18241 191051
rect 18269 191023 18303 191051
rect 18331 191023 33477 191051
rect 33505 191023 33539 191051
rect 33567 191023 33601 191051
rect 33629 191023 33663 191051
rect 33691 191023 48837 191051
rect 48865 191023 48899 191051
rect 48927 191023 48961 191051
rect 48989 191023 49023 191051
rect 49051 191023 64197 191051
rect 64225 191023 64259 191051
rect 64287 191023 64321 191051
rect 64349 191023 64383 191051
rect 64411 191023 79557 191051
rect 79585 191023 79619 191051
rect 79647 191023 79681 191051
rect 79709 191023 79743 191051
rect 79771 191023 94917 191051
rect 94945 191023 94979 191051
rect 95007 191023 95041 191051
rect 95069 191023 95103 191051
rect 95131 191023 110277 191051
rect 110305 191023 110339 191051
rect 110367 191023 110401 191051
rect 110429 191023 110463 191051
rect 110491 191023 125637 191051
rect 125665 191023 125699 191051
rect 125727 191023 125761 191051
rect 125789 191023 125823 191051
rect 125851 191023 140997 191051
rect 141025 191023 141059 191051
rect 141087 191023 141121 191051
rect 141149 191023 141183 191051
rect 141211 191023 156357 191051
rect 156385 191023 156419 191051
rect 156447 191023 156481 191051
rect 156509 191023 156543 191051
rect 156571 191023 171717 191051
rect 171745 191023 171779 191051
rect 171807 191023 171841 191051
rect 171869 191023 171903 191051
rect 171931 191023 187077 191051
rect 187105 191023 187139 191051
rect 187167 191023 187201 191051
rect 187229 191023 187263 191051
rect 187291 191023 202437 191051
rect 202465 191023 202499 191051
rect 202527 191023 202561 191051
rect 202589 191023 202623 191051
rect 202651 191023 217797 191051
rect 217825 191023 217859 191051
rect 217887 191023 217921 191051
rect 217949 191023 217983 191051
rect 218011 191023 233157 191051
rect 233185 191023 233219 191051
rect 233247 191023 233281 191051
rect 233309 191023 233343 191051
rect 233371 191023 248517 191051
rect 248545 191023 248579 191051
rect 248607 191023 248641 191051
rect 248669 191023 248703 191051
rect 248731 191023 263877 191051
rect 263905 191023 263939 191051
rect 263967 191023 264001 191051
rect 264029 191023 264063 191051
rect 264091 191023 279237 191051
rect 279265 191023 279299 191051
rect 279327 191023 279361 191051
rect 279389 191023 279423 191051
rect 279451 191023 294597 191051
rect 294625 191023 294659 191051
rect 294687 191023 294721 191051
rect 294749 191023 294783 191051
rect 294811 191023 298248 191051
rect 298276 191023 298310 191051
rect 298338 191023 298372 191051
rect 298400 191023 298434 191051
rect 298462 191023 298990 191051
rect -958 190989 298990 191023
rect -958 190961 -430 190989
rect -402 190961 -368 190989
rect -340 190961 -306 190989
rect -278 190961 -244 190989
rect -216 190961 2757 190989
rect 2785 190961 2819 190989
rect 2847 190961 2881 190989
rect 2909 190961 2943 190989
rect 2971 190961 18117 190989
rect 18145 190961 18179 190989
rect 18207 190961 18241 190989
rect 18269 190961 18303 190989
rect 18331 190961 33477 190989
rect 33505 190961 33539 190989
rect 33567 190961 33601 190989
rect 33629 190961 33663 190989
rect 33691 190961 48837 190989
rect 48865 190961 48899 190989
rect 48927 190961 48961 190989
rect 48989 190961 49023 190989
rect 49051 190961 64197 190989
rect 64225 190961 64259 190989
rect 64287 190961 64321 190989
rect 64349 190961 64383 190989
rect 64411 190961 79557 190989
rect 79585 190961 79619 190989
rect 79647 190961 79681 190989
rect 79709 190961 79743 190989
rect 79771 190961 94917 190989
rect 94945 190961 94979 190989
rect 95007 190961 95041 190989
rect 95069 190961 95103 190989
rect 95131 190961 110277 190989
rect 110305 190961 110339 190989
rect 110367 190961 110401 190989
rect 110429 190961 110463 190989
rect 110491 190961 125637 190989
rect 125665 190961 125699 190989
rect 125727 190961 125761 190989
rect 125789 190961 125823 190989
rect 125851 190961 140997 190989
rect 141025 190961 141059 190989
rect 141087 190961 141121 190989
rect 141149 190961 141183 190989
rect 141211 190961 156357 190989
rect 156385 190961 156419 190989
rect 156447 190961 156481 190989
rect 156509 190961 156543 190989
rect 156571 190961 171717 190989
rect 171745 190961 171779 190989
rect 171807 190961 171841 190989
rect 171869 190961 171903 190989
rect 171931 190961 187077 190989
rect 187105 190961 187139 190989
rect 187167 190961 187201 190989
rect 187229 190961 187263 190989
rect 187291 190961 202437 190989
rect 202465 190961 202499 190989
rect 202527 190961 202561 190989
rect 202589 190961 202623 190989
rect 202651 190961 217797 190989
rect 217825 190961 217859 190989
rect 217887 190961 217921 190989
rect 217949 190961 217983 190989
rect 218011 190961 233157 190989
rect 233185 190961 233219 190989
rect 233247 190961 233281 190989
rect 233309 190961 233343 190989
rect 233371 190961 248517 190989
rect 248545 190961 248579 190989
rect 248607 190961 248641 190989
rect 248669 190961 248703 190989
rect 248731 190961 263877 190989
rect 263905 190961 263939 190989
rect 263967 190961 264001 190989
rect 264029 190961 264063 190989
rect 264091 190961 279237 190989
rect 279265 190961 279299 190989
rect 279327 190961 279361 190989
rect 279389 190961 279423 190989
rect 279451 190961 294597 190989
rect 294625 190961 294659 190989
rect 294687 190961 294721 190989
rect 294749 190961 294783 190989
rect 294811 190961 298248 190989
rect 298276 190961 298310 190989
rect 298338 190961 298372 190989
rect 298400 190961 298434 190989
rect 298462 190961 298990 190989
rect -958 190913 298990 190961
rect -958 185175 298990 185223
rect -958 185147 -910 185175
rect -882 185147 -848 185175
rect -820 185147 -786 185175
rect -758 185147 -724 185175
rect -696 185147 4617 185175
rect 4645 185147 4679 185175
rect 4707 185147 4741 185175
rect 4769 185147 4803 185175
rect 4831 185147 19977 185175
rect 20005 185147 20039 185175
rect 20067 185147 20101 185175
rect 20129 185147 20163 185175
rect 20191 185147 35337 185175
rect 35365 185147 35399 185175
rect 35427 185147 35461 185175
rect 35489 185147 35523 185175
rect 35551 185147 50697 185175
rect 50725 185147 50759 185175
rect 50787 185147 50821 185175
rect 50849 185147 50883 185175
rect 50911 185147 66057 185175
rect 66085 185147 66119 185175
rect 66147 185147 66181 185175
rect 66209 185147 66243 185175
rect 66271 185147 81417 185175
rect 81445 185147 81479 185175
rect 81507 185147 81541 185175
rect 81569 185147 81603 185175
rect 81631 185147 96777 185175
rect 96805 185147 96839 185175
rect 96867 185147 96901 185175
rect 96929 185147 96963 185175
rect 96991 185147 112137 185175
rect 112165 185147 112199 185175
rect 112227 185147 112261 185175
rect 112289 185147 112323 185175
rect 112351 185147 127497 185175
rect 127525 185147 127559 185175
rect 127587 185147 127621 185175
rect 127649 185147 127683 185175
rect 127711 185147 142857 185175
rect 142885 185147 142919 185175
rect 142947 185147 142981 185175
rect 143009 185147 143043 185175
rect 143071 185147 158217 185175
rect 158245 185147 158279 185175
rect 158307 185147 158341 185175
rect 158369 185147 158403 185175
rect 158431 185147 173577 185175
rect 173605 185147 173639 185175
rect 173667 185147 173701 185175
rect 173729 185147 173763 185175
rect 173791 185147 188937 185175
rect 188965 185147 188999 185175
rect 189027 185147 189061 185175
rect 189089 185147 189123 185175
rect 189151 185147 204297 185175
rect 204325 185147 204359 185175
rect 204387 185147 204421 185175
rect 204449 185147 204483 185175
rect 204511 185147 219657 185175
rect 219685 185147 219719 185175
rect 219747 185147 219781 185175
rect 219809 185147 219843 185175
rect 219871 185147 235017 185175
rect 235045 185147 235079 185175
rect 235107 185147 235141 185175
rect 235169 185147 235203 185175
rect 235231 185147 250377 185175
rect 250405 185147 250439 185175
rect 250467 185147 250501 185175
rect 250529 185147 250563 185175
rect 250591 185147 265737 185175
rect 265765 185147 265799 185175
rect 265827 185147 265861 185175
rect 265889 185147 265923 185175
rect 265951 185147 281097 185175
rect 281125 185147 281159 185175
rect 281187 185147 281221 185175
rect 281249 185147 281283 185175
rect 281311 185147 296457 185175
rect 296485 185147 296519 185175
rect 296547 185147 296581 185175
rect 296609 185147 296643 185175
rect 296671 185147 298728 185175
rect 298756 185147 298790 185175
rect 298818 185147 298852 185175
rect 298880 185147 298914 185175
rect 298942 185147 298990 185175
rect -958 185113 298990 185147
rect -958 185085 -910 185113
rect -882 185085 -848 185113
rect -820 185085 -786 185113
rect -758 185085 -724 185113
rect -696 185085 4617 185113
rect 4645 185085 4679 185113
rect 4707 185085 4741 185113
rect 4769 185085 4803 185113
rect 4831 185085 19977 185113
rect 20005 185085 20039 185113
rect 20067 185085 20101 185113
rect 20129 185085 20163 185113
rect 20191 185085 35337 185113
rect 35365 185085 35399 185113
rect 35427 185085 35461 185113
rect 35489 185085 35523 185113
rect 35551 185085 50697 185113
rect 50725 185085 50759 185113
rect 50787 185085 50821 185113
rect 50849 185085 50883 185113
rect 50911 185085 66057 185113
rect 66085 185085 66119 185113
rect 66147 185085 66181 185113
rect 66209 185085 66243 185113
rect 66271 185085 81417 185113
rect 81445 185085 81479 185113
rect 81507 185085 81541 185113
rect 81569 185085 81603 185113
rect 81631 185085 96777 185113
rect 96805 185085 96839 185113
rect 96867 185085 96901 185113
rect 96929 185085 96963 185113
rect 96991 185085 112137 185113
rect 112165 185085 112199 185113
rect 112227 185085 112261 185113
rect 112289 185085 112323 185113
rect 112351 185085 127497 185113
rect 127525 185085 127559 185113
rect 127587 185085 127621 185113
rect 127649 185085 127683 185113
rect 127711 185085 142857 185113
rect 142885 185085 142919 185113
rect 142947 185085 142981 185113
rect 143009 185085 143043 185113
rect 143071 185085 158217 185113
rect 158245 185085 158279 185113
rect 158307 185085 158341 185113
rect 158369 185085 158403 185113
rect 158431 185085 173577 185113
rect 173605 185085 173639 185113
rect 173667 185085 173701 185113
rect 173729 185085 173763 185113
rect 173791 185085 188937 185113
rect 188965 185085 188999 185113
rect 189027 185085 189061 185113
rect 189089 185085 189123 185113
rect 189151 185085 204297 185113
rect 204325 185085 204359 185113
rect 204387 185085 204421 185113
rect 204449 185085 204483 185113
rect 204511 185085 219657 185113
rect 219685 185085 219719 185113
rect 219747 185085 219781 185113
rect 219809 185085 219843 185113
rect 219871 185085 235017 185113
rect 235045 185085 235079 185113
rect 235107 185085 235141 185113
rect 235169 185085 235203 185113
rect 235231 185085 250377 185113
rect 250405 185085 250439 185113
rect 250467 185085 250501 185113
rect 250529 185085 250563 185113
rect 250591 185085 265737 185113
rect 265765 185085 265799 185113
rect 265827 185085 265861 185113
rect 265889 185085 265923 185113
rect 265951 185085 281097 185113
rect 281125 185085 281159 185113
rect 281187 185085 281221 185113
rect 281249 185085 281283 185113
rect 281311 185085 296457 185113
rect 296485 185085 296519 185113
rect 296547 185085 296581 185113
rect 296609 185085 296643 185113
rect 296671 185085 298728 185113
rect 298756 185085 298790 185113
rect 298818 185085 298852 185113
rect 298880 185085 298914 185113
rect 298942 185085 298990 185113
rect -958 185051 298990 185085
rect -958 185023 -910 185051
rect -882 185023 -848 185051
rect -820 185023 -786 185051
rect -758 185023 -724 185051
rect -696 185023 4617 185051
rect 4645 185023 4679 185051
rect 4707 185023 4741 185051
rect 4769 185023 4803 185051
rect 4831 185023 19977 185051
rect 20005 185023 20039 185051
rect 20067 185023 20101 185051
rect 20129 185023 20163 185051
rect 20191 185023 35337 185051
rect 35365 185023 35399 185051
rect 35427 185023 35461 185051
rect 35489 185023 35523 185051
rect 35551 185023 50697 185051
rect 50725 185023 50759 185051
rect 50787 185023 50821 185051
rect 50849 185023 50883 185051
rect 50911 185023 66057 185051
rect 66085 185023 66119 185051
rect 66147 185023 66181 185051
rect 66209 185023 66243 185051
rect 66271 185023 81417 185051
rect 81445 185023 81479 185051
rect 81507 185023 81541 185051
rect 81569 185023 81603 185051
rect 81631 185023 96777 185051
rect 96805 185023 96839 185051
rect 96867 185023 96901 185051
rect 96929 185023 96963 185051
rect 96991 185023 112137 185051
rect 112165 185023 112199 185051
rect 112227 185023 112261 185051
rect 112289 185023 112323 185051
rect 112351 185023 127497 185051
rect 127525 185023 127559 185051
rect 127587 185023 127621 185051
rect 127649 185023 127683 185051
rect 127711 185023 142857 185051
rect 142885 185023 142919 185051
rect 142947 185023 142981 185051
rect 143009 185023 143043 185051
rect 143071 185023 158217 185051
rect 158245 185023 158279 185051
rect 158307 185023 158341 185051
rect 158369 185023 158403 185051
rect 158431 185023 173577 185051
rect 173605 185023 173639 185051
rect 173667 185023 173701 185051
rect 173729 185023 173763 185051
rect 173791 185023 188937 185051
rect 188965 185023 188999 185051
rect 189027 185023 189061 185051
rect 189089 185023 189123 185051
rect 189151 185023 204297 185051
rect 204325 185023 204359 185051
rect 204387 185023 204421 185051
rect 204449 185023 204483 185051
rect 204511 185023 219657 185051
rect 219685 185023 219719 185051
rect 219747 185023 219781 185051
rect 219809 185023 219843 185051
rect 219871 185023 235017 185051
rect 235045 185023 235079 185051
rect 235107 185023 235141 185051
rect 235169 185023 235203 185051
rect 235231 185023 250377 185051
rect 250405 185023 250439 185051
rect 250467 185023 250501 185051
rect 250529 185023 250563 185051
rect 250591 185023 265737 185051
rect 265765 185023 265799 185051
rect 265827 185023 265861 185051
rect 265889 185023 265923 185051
rect 265951 185023 281097 185051
rect 281125 185023 281159 185051
rect 281187 185023 281221 185051
rect 281249 185023 281283 185051
rect 281311 185023 296457 185051
rect 296485 185023 296519 185051
rect 296547 185023 296581 185051
rect 296609 185023 296643 185051
rect 296671 185023 298728 185051
rect 298756 185023 298790 185051
rect 298818 185023 298852 185051
rect 298880 185023 298914 185051
rect 298942 185023 298990 185051
rect -958 184989 298990 185023
rect -958 184961 -910 184989
rect -882 184961 -848 184989
rect -820 184961 -786 184989
rect -758 184961 -724 184989
rect -696 184961 4617 184989
rect 4645 184961 4679 184989
rect 4707 184961 4741 184989
rect 4769 184961 4803 184989
rect 4831 184961 19977 184989
rect 20005 184961 20039 184989
rect 20067 184961 20101 184989
rect 20129 184961 20163 184989
rect 20191 184961 35337 184989
rect 35365 184961 35399 184989
rect 35427 184961 35461 184989
rect 35489 184961 35523 184989
rect 35551 184961 50697 184989
rect 50725 184961 50759 184989
rect 50787 184961 50821 184989
rect 50849 184961 50883 184989
rect 50911 184961 66057 184989
rect 66085 184961 66119 184989
rect 66147 184961 66181 184989
rect 66209 184961 66243 184989
rect 66271 184961 81417 184989
rect 81445 184961 81479 184989
rect 81507 184961 81541 184989
rect 81569 184961 81603 184989
rect 81631 184961 96777 184989
rect 96805 184961 96839 184989
rect 96867 184961 96901 184989
rect 96929 184961 96963 184989
rect 96991 184961 112137 184989
rect 112165 184961 112199 184989
rect 112227 184961 112261 184989
rect 112289 184961 112323 184989
rect 112351 184961 127497 184989
rect 127525 184961 127559 184989
rect 127587 184961 127621 184989
rect 127649 184961 127683 184989
rect 127711 184961 142857 184989
rect 142885 184961 142919 184989
rect 142947 184961 142981 184989
rect 143009 184961 143043 184989
rect 143071 184961 158217 184989
rect 158245 184961 158279 184989
rect 158307 184961 158341 184989
rect 158369 184961 158403 184989
rect 158431 184961 173577 184989
rect 173605 184961 173639 184989
rect 173667 184961 173701 184989
rect 173729 184961 173763 184989
rect 173791 184961 188937 184989
rect 188965 184961 188999 184989
rect 189027 184961 189061 184989
rect 189089 184961 189123 184989
rect 189151 184961 204297 184989
rect 204325 184961 204359 184989
rect 204387 184961 204421 184989
rect 204449 184961 204483 184989
rect 204511 184961 219657 184989
rect 219685 184961 219719 184989
rect 219747 184961 219781 184989
rect 219809 184961 219843 184989
rect 219871 184961 235017 184989
rect 235045 184961 235079 184989
rect 235107 184961 235141 184989
rect 235169 184961 235203 184989
rect 235231 184961 250377 184989
rect 250405 184961 250439 184989
rect 250467 184961 250501 184989
rect 250529 184961 250563 184989
rect 250591 184961 265737 184989
rect 265765 184961 265799 184989
rect 265827 184961 265861 184989
rect 265889 184961 265923 184989
rect 265951 184961 281097 184989
rect 281125 184961 281159 184989
rect 281187 184961 281221 184989
rect 281249 184961 281283 184989
rect 281311 184961 296457 184989
rect 296485 184961 296519 184989
rect 296547 184961 296581 184989
rect 296609 184961 296643 184989
rect 296671 184961 298728 184989
rect 298756 184961 298790 184989
rect 298818 184961 298852 184989
rect 298880 184961 298914 184989
rect 298942 184961 298990 184989
rect -958 184913 298990 184961
rect -958 182175 298990 182223
rect -958 182147 -430 182175
rect -402 182147 -368 182175
rect -340 182147 -306 182175
rect -278 182147 -244 182175
rect -216 182147 2757 182175
rect 2785 182147 2819 182175
rect 2847 182147 2881 182175
rect 2909 182147 2943 182175
rect 2971 182147 18117 182175
rect 18145 182147 18179 182175
rect 18207 182147 18241 182175
rect 18269 182147 18303 182175
rect 18331 182147 33477 182175
rect 33505 182147 33539 182175
rect 33567 182147 33601 182175
rect 33629 182147 33663 182175
rect 33691 182147 48837 182175
rect 48865 182147 48899 182175
rect 48927 182147 48961 182175
rect 48989 182147 49023 182175
rect 49051 182147 64197 182175
rect 64225 182147 64259 182175
rect 64287 182147 64321 182175
rect 64349 182147 64383 182175
rect 64411 182147 79557 182175
rect 79585 182147 79619 182175
rect 79647 182147 79681 182175
rect 79709 182147 79743 182175
rect 79771 182147 94917 182175
rect 94945 182147 94979 182175
rect 95007 182147 95041 182175
rect 95069 182147 95103 182175
rect 95131 182147 110277 182175
rect 110305 182147 110339 182175
rect 110367 182147 110401 182175
rect 110429 182147 110463 182175
rect 110491 182147 125637 182175
rect 125665 182147 125699 182175
rect 125727 182147 125761 182175
rect 125789 182147 125823 182175
rect 125851 182147 140997 182175
rect 141025 182147 141059 182175
rect 141087 182147 141121 182175
rect 141149 182147 141183 182175
rect 141211 182147 156357 182175
rect 156385 182147 156419 182175
rect 156447 182147 156481 182175
rect 156509 182147 156543 182175
rect 156571 182147 171717 182175
rect 171745 182147 171779 182175
rect 171807 182147 171841 182175
rect 171869 182147 171903 182175
rect 171931 182147 187077 182175
rect 187105 182147 187139 182175
rect 187167 182147 187201 182175
rect 187229 182147 187263 182175
rect 187291 182147 202437 182175
rect 202465 182147 202499 182175
rect 202527 182147 202561 182175
rect 202589 182147 202623 182175
rect 202651 182147 217797 182175
rect 217825 182147 217859 182175
rect 217887 182147 217921 182175
rect 217949 182147 217983 182175
rect 218011 182147 233157 182175
rect 233185 182147 233219 182175
rect 233247 182147 233281 182175
rect 233309 182147 233343 182175
rect 233371 182147 248517 182175
rect 248545 182147 248579 182175
rect 248607 182147 248641 182175
rect 248669 182147 248703 182175
rect 248731 182147 263877 182175
rect 263905 182147 263939 182175
rect 263967 182147 264001 182175
rect 264029 182147 264063 182175
rect 264091 182147 279237 182175
rect 279265 182147 279299 182175
rect 279327 182147 279361 182175
rect 279389 182147 279423 182175
rect 279451 182147 294597 182175
rect 294625 182147 294659 182175
rect 294687 182147 294721 182175
rect 294749 182147 294783 182175
rect 294811 182147 298248 182175
rect 298276 182147 298310 182175
rect 298338 182147 298372 182175
rect 298400 182147 298434 182175
rect 298462 182147 298990 182175
rect -958 182113 298990 182147
rect -958 182085 -430 182113
rect -402 182085 -368 182113
rect -340 182085 -306 182113
rect -278 182085 -244 182113
rect -216 182085 2757 182113
rect 2785 182085 2819 182113
rect 2847 182085 2881 182113
rect 2909 182085 2943 182113
rect 2971 182085 18117 182113
rect 18145 182085 18179 182113
rect 18207 182085 18241 182113
rect 18269 182085 18303 182113
rect 18331 182085 33477 182113
rect 33505 182085 33539 182113
rect 33567 182085 33601 182113
rect 33629 182085 33663 182113
rect 33691 182085 48837 182113
rect 48865 182085 48899 182113
rect 48927 182085 48961 182113
rect 48989 182085 49023 182113
rect 49051 182085 64197 182113
rect 64225 182085 64259 182113
rect 64287 182085 64321 182113
rect 64349 182085 64383 182113
rect 64411 182085 79557 182113
rect 79585 182085 79619 182113
rect 79647 182085 79681 182113
rect 79709 182085 79743 182113
rect 79771 182085 94917 182113
rect 94945 182085 94979 182113
rect 95007 182085 95041 182113
rect 95069 182085 95103 182113
rect 95131 182085 110277 182113
rect 110305 182085 110339 182113
rect 110367 182085 110401 182113
rect 110429 182085 110463 182113
rect 110491 182085 125637 182113
rect 125665 182085 125699 182113
rect 125727 182085 125761 182113
rect 125789 182085 125823 182113
rect 125851 182085 140997 182113
rect 141025 182085 141059 182113
rect 141087 182085 141121 182113
rect 141149 182085 141183 182113
rect 141211 182085 156357 182113
rect 156385 182085 156419 182113
rect 156447 182085 156481 182113
rect 156509 182085 156543 182113
rect 156571 182085 171717 182113
rect 171745 182085 171779 182113
rect 171807 182085 171841 182113
rect 171869 182085 171903 182113
rect 171931 182085 187077 182113
rect 187105 182085 187139 182113
rect 187167 182085 187201 182113
rect 187229 182085 187263 182113
rect 187291 182085 202437 182113
rect 202465 182085 202499 182113
rect 202527 182085 202561 182113
rect 202589 182085 202623 182113
rect 202651 182085 217797 182113
rect 217825 182085 217859 182113
rect 217887 182085 217921 182113
rect 217949 182085 217983 182113
rect 218011 182085 233157 182113
rect 233185 182085 233219 182113
rect 233247 182085 233281 182113
rect 233309 182085 233343 182113
rect 233371 182085 248517 182113
rect 248545 182085 248579 182113
rect 248607 182085 248641 182113
rect 248669 182085 248703 182113
rect 248731 182085 263877 182113
rect 263905 182085 263939 182113
rect 263967 182085 264001 182113
rect 264029 182085 264063 182113
rect 264091 182085 279237 182113
rect 279265 182085 279299 182113
rect 279327 182085 279361 182113
rect 279389 182085 279423 182113
rect 279451 182085 294597 182113
rect 294625 182085 294659 182113
rect 294687 182085 294721 182113
rect 294749 182085 294783 182113
rect 294811 182085 298248 182113
rect 298276 182085 298310 182113
rect 298338 182085 298372 182113
rect 298400 182085 298434 182113
rect 298462 182085 298990 182113
rect -958 182051 298990 182085
rect -958 182023 -430 182051
rect -402 182023 -368 182051
rect -340 182023 -306 182051
rect -278 182023 -244 182051
rect -216 182023 2757 182051
rect 2785 182023 2819 182051
rect 2847 182023 2881 182051
rect 2909 182023 2943 182051
rect 2971 182023 18117 182051
rect 18145 182023 18179 182051
rect 18207 182023 18241 182051
rect 18269 182023 18303 182051
rect 18331 182023 33477 182051
rect 33505 182023 33539 182051
rect 33567 182023 33601 182051
rect 33629 182023 33663 182051
rect 33691 182023 48837 182051
rect 48865 182023 48899 182051
rect 48927 182023 48961 182051
rect 48989 182023 49023 182051
rect 49051 182023 64197 182051
rect 64225 182023 64259 182051
rect 64287 182023 64321 182051
rect 64349 182023 64383 182051
rect 64411 182023 79557 182051
rect 79585 182023 79619 182051
rect 79647 182023 79681 182051
rect 79709 182023 79743 182051
rect 79771 182023 94917 182051
rect 94945 182023 94979 182051
rect 95007 182023 95041 182051
rect 95069 182023 95103 182051
rect 95131 182023 110277 182051
rect 110305 182023 110339 182051
rect 110367 182023 110401 182051
rect 110429 182023 110463 182051
rect 110491 182023 125637 182051
rect 125665 182023 125699 182051
rect 125727 182023 125761 182051
rect 125789 182023 125823 182051
rect 125851 182023 140997 182051
rect 141025 182023 141059 182051
rect 141087 182023 141121 182051
rect 141149 182023 141183 182051
rect 141211 182023 156357 182051
rect 156385 182023 156419 182051
rect 156447 182023 156481 182051
rect 156509 182023 156543 182051
rect 156571 182023 171717 182051
rect 171745 182023 171779 182051
rect 171807 182023 171841 182051
rect 171869 182023 171903 182051
rect 171931 182023 187077 182051
rect 187105 182023 187139 182051
rect 187167 182023 187201 182051
rect 187229 182023 187263 182051
rect 187291 182023 202437 182051
rect 202465 182023 202499 182051
rect 202527 182023 202561 182051
rect 202589 182023 202623 182051
rect 202651 182023 217797 182051
rect 217825 182023 217859 182051
rect 217887 182023 217921 182051
rect 217949 182023 217983 182051
rect 218011 182023 233157 182051
rect 233185 182023 233219 182051
rect 233247 182023 233281 182051
rect 233309 182023 233343 182051
rect 233371 182023 248517 182051
rect 248545 182023 248579 182051
rect 248607 182023 248641 182051
rect 248669 182023 248703 182051
rect 248731 182023 263877 182051
rect 263905 182023 263939 182051
rect 263967 182023 264001 182051
rect 264029 182023 264063 182051
rect 264091 182023 279237 182051
rect 279265 182023 279299 182051
rect 279327 182023 279361 182051
rect 279389 182023 279423 182051
rect 279451 182023 294597 182051
rect 294625 182023 294659 182051
rect 294687 182023 294721 182051
rect 294749 182023 294783 182051
rect 294811 182023 298248 182051
rect 298276 182023 298310 182051
rect 298338 182023 298372 182051
rect 298400 182023 298434 182051
rect 298462 182023 298990 182051
rect -958 181989 298990 182023
rect -958 181961 -430 181989
rect -402 181961 -368 181989
rect -340 181961 -306 181989
rect -278 181961 -244 181989
rect -216 181961 2757 181989
rect 2785 181961 2819 181989
rect 2847 181961 2881 181989
rect 2909 181961 2943 181989
rect 2971 181961 18117 181989
rect 18145 181961 18179 181989
rect 18207 181961 18241 181989
rect 18269 181961 18303 181989
rect 18331 181961 33477 181989
rect 33505 181961 33539 181989
rect 33567 181961 33601 181989
rect 33629 181961 33663 181989
rect 33691 181961 48837 181989
rect 48865 181961 48899 181989
rect 48927 181961 48961 181989
rect 48989 181961 49023 181989
rect 49051 181961 64197 181989
rect 64225 181961 64259 181989
rect 64287 181961 64321 181989
rect 64349 181961 64383 181989
rect 64411 181961 79557 181989
rect 79585 181961 79619 181989
rect 79647 181961 79681 181989
rect 79709 181961 79743 181989
rect 79771 181961 94917 181989
rect 94945 181961 94979 181989
rect 95007 181961 95041 181989
rect 95069 181961 95103 181989
rect 95131 181961 110277 181989
rect 110305 181961 110339 181989
rect 110367 181961 110401 181989
rect 110429 181961 110463 181989
rect 110491 181961 125637 181989
rect 125665 181961 125699 181989
rect 125727 181961 125761 181989
rect 125789 181961 125823 181989
rect 125851 181961 140997 181989
rect 141025 181961 141059 181989
rect 141087 181961 141121 181989
rect 141149 181961 141183 181989
rect 141211 181961 156357 181989
rect 156385 181961 156419 181989
rect 156447 181961 156481 181989
rect 156509 181961 156543 181989
rect 156571 181961 171717 181989
rect 171745 181961 171779 181989
rect 171807 181961 171841 181989
rect 171869 181961 171903 181989
rect 171931 181961 187077 181989
rect 187105 181961 187139 181989
rect 187167 181961 187201 181989
rect 187229 181961 187263 181989
rect 187291 181961 202437 181989
rect 202465 181961 202499 181989
rect 202527 181961 202561 181989
rect 202589 181961 202623 181989
rect 202651 181961 217797 181989
rect 217825 181961 217859 181989
rect 217887 181961 217921 181989
rect 217949 181961 217983 181989
rect 218011 181961 233157 181989
rect 233185 181961 233219 181989
rect 233247 181961 233281 181989
rect 233309 181961 233343 181989
rect 233371 181961 248517 181989
rect 248545 181961 248579 181989
rect 248607 181961 248641 181989
rect 248669 181961 248703 181989
rect 248731 181961 263877 181989
rect 263905 181961 263939 181989
rect 263967 181961 264001 181989
rect 264029 181961 264063 181989
rect 264091 181961 279237 181989
rect 279265 181961 279299 181989
rect 279327 181961 279361 181989
rect 279389 181961 279423 181989
rect 279451 181961 294597 181989
rect 294625 181961 294659 181989
rect 294687 181961 294721 181989
rect 294749 181961 294783 181989
rect 294811 181961 298248 181989
rect 298276 181961 298310 181989
rect 298338 181961 298372 181989
rect 298400 181961 298434 181989
rect 298462 181961 298990 181989
rect -958 181913 298990 181961
rect -958 176175 298990 176223
rect -958 176147 -910 176175
rect -882 176147 -848 176175
rect -820 176147 -786 176175
rect -758 176147 -724 176175
rect -696 176147 4617 176175
rect 4645 176147 4679 176175
rect 4707 176147 4741 176175
rect 4769 176147 4803 176175
rect 4831 176147 19977 176175
rect 20005 176147 20039 176175
rect 20067 176147 20101 176175
rect 20129 176147 20163 176175
rect 20191 176147 35337 176175
rect 35365 176147 35399 176175
rect 35427 176147 35461 176175
rect 35489 176147 35523 176175
rect 35551 176147 50697 176175
rect 50725 176147 50759 176175
rect 50787 176147 50821 176175
rect 50849 176147 50883 176175
rect 50911 176147 66057 176175
rect 66085 176147 66119 176175
rect 66147 176147 66181 176175
rect 66209 176147 66243 176175
rect 66271 176147 81417 176175
rect 81445 176147 81479 176175
rect 81507 176147 81541 176175
rect 81569 176147 81603 176175
rect 81631 176147 96777 176175
rect 96805 176147 96839 176175
rect 96867 176147 96901 176175
rect 96929 176147 96963 176175
rect 96991 176147 112137 176175
rect 112165 176147 112199 176175
rect 112227 176147 112261 176175
rect 112289 176147 112323 176175
rect 112351 176147 127497 176175
rect 127525 176147 127559 176175
rect 127587 176147 127621 176175
rect 127649 176147 127683 176175
rect 127711 176147 142857 176175
rect 142885 176147 142919 176175
rect 142947 176147 142981 176175
rect 143009 176147 143043 176175
rect 143071 176147 158217 176175
rect 158245 176147 158279 176175
rect 158307 176147 158341 176175
rect 158369 176147 158403 176175
rect 158431 176147 173577 176175
rect 173605 176147 173639 176175
rect 173667 176147 173701 176175
rect 173729 176147 173763 176175
rect 173791 176147 188937 176175
rect 188965 176147 188999 176175
rect 189027 176147 189061 176175
rect 189089 176147 189123 176175
rect 189151 176147 204297 176175
rect 204325 176147 204359 176175
rect 204387 176147 204421 176175
rect 204449 176147 204483 176175
rect 204511 176147 219657 176175
rect 219685 176147 219719 176175
rect 219747 176147 219781 176175
rect 219809 176147 219843 176175
rect 219871 176147 235017 176175
rect 235045 176147 235079 176175
rect 235107 176147 235141 176175
rect 235169 176147 235203 176175
rect 235231 176147 250377 176175
rect 250405 176147 250439 176175
rect 250467 176147 250501 176175
rect 250529 176147 250563 176175
rect 250591 176147 265737 176175
rect 265765 176147 265799 176175
rect 265827 176147 265861 176175
rect 265889 176147 265923 176175
rect 265951 176147 281097 176175
rect 281125 176147 281159 176175
rect 281187 176147 281221 176175
rect 281249 176147 281283 176175
rect 281311 176147 296457 176175
rect 296485 176147 296519 176175
rect 296547 176147 296581 176175
rect 296609 176147 296643 176175
rect 296671 176147 298728 176175
rect 298756 176147 298790 176175
rect 298818 176147 298852 176175
rect 298880 176147 298914 176175
rect 298942 176147 298990 176175
rect -958 176113 298990 176147
rect -958 176085 -910 176113
rect -882 176085 -848 176113
rect -820 176085 -786 176113
rect -758 176085 -724 176113
rect -696 176085 4617 176113
rect 4645 176085 4679 176113
rect 4707 176085 4741 176113
rect 4769 176085 4803 176113
rect 4831 176085 19977 176113
rect 20005 176085 20039 176113
rect 20067 176085 20101 176113
rect 20129 176085 20163 176113
rect 20191 176085 35337 176113
rect 35365 176085 35399 176113
rect 35427 176085 35461 176113
rect 35489 176085 35523 176113
rect 35551 176085 50697 176113
rect 50725 176085 50759 176113
rect 50787 176085 50821 176113
rect 50849 176085 50883 176113
rect 50911 176085 66057 176113
rect 66085 176085 66119 176113
rect 66147 176085 66181 176113
rect 66209 176085 66243 176113
rect 66271 176085 81417 176113
rect 81445 176085 81479 176113
rect 81507 176085 81541 176113
rect 81569 176085 81603 176113
rect 81631 176085 96777 176113
rect 96805 176085 96839 176113
rect 96867 176085 96901 176113
rect 96929 176085 96963 176113
rect 96991 176085 112137 176113
rect 112165 176085 112199 176113
rect 112227 176085 112261 176113
rect 112289 176085 112323 176113
rect 112351 176085 127497 176113
rect 127525 176085 127559 176113
rect 127587 176085 127621 176113
rect 127649 176085 127683 176113
rect 127711 176085 142857 176113
rect 142885 176085 142919 176113
rect 142947 176085 142981 176113
rect 143009 176085 143043 176113
rect 143071 176085 158217 176113
rect 158245 176085 158279 176113
rect 158307 176085 158341 176113
rect 158369 176085 158403 176113
rect 158431 176085 173577 176113
rect 173605 176085 173639 176113
rect 173667 176085 173701 176113
rect 173729 176085 173763 176113
rect 173791 176085 188937 176113
rect 188965 176085 188999 176113
rect 189027 176085 189061 176113
rect 189089 176085 189123 176113
rect 189151 176085 204297 176113
rect 204325 176085 204359 176113
rect 204387 176085 204421 176113
rect 204449 176085 204483 176113
rect 204511 176085 219657 176113
rect 219685 176085 219719 176113
rect 219747 176085 219781 176113
rect 219809 176085 219843 176113
rect 219871 176085 235017 176113
rect 235045 176085 235079 176113
rect 235107 176085 235141 176113
rect 235169 176085 235203 176113
rect 235231 176085 250377 176113
rect 250405 176085 250439 176113
rect 250467 176085 250501 176113
rect 250529 176085 250563 176113
rect 250591 176085 265737 176113
rect 265765 176085 265799 176113
rect 265827 176085 265861 176113
rect 265889 176085 265923 176113
rect 265951 176085 281097 176113
rect 281125 176085 281159 176113
rect 281187 176085 281221 176113
rect 281249 176085 281283 176113
rect 281311 176085 296457 176113
rect 296485 176085 296519 176113
rect 296547 176085 296581 176113
rect 296609 176085 296643 176113
rect 296671 176085 298728 176113
rect 298756 176085 298790 176113
rect 298818 176085 298852 176113
rect 298880 176085 298914 176113
rect 298942 176085 298990 176113
rect -958 176051 298990 176085
rect -958 176023 -910 176051
rect -882 176023 -848 176051
rect -820 176023 -786 176051
rect -758 176023 -724 176051
rect -696 176023 4617 176051
rect 4645 176023 4679 176051
rect 4707 176023 4741 176051
rect 4769 176023 4803 176051
rect 4831 176023 19977 176051
rect 20005 176023 20039 176051
rect 20067 176023 20101 176051
rect 20129 176023 20163 176051
rect 20191 176023 35337 176051
rect 35365 176023 35399 176051
rect 35427 176023 35461 176051
rect 35489 176023 35523 176051
rect 35551 176023 50697 176051
rect 50725 176023 50759 176051
rect 50787 176023 50821 176051
rect 50849 176023 50883 176051
rect 50911 176023 66057 176051
rect 66085 176023 66119 176051
rect 66147 176023 66181 176051
rect 66209 176023 66243 176051
rect 66271 176023 81417 176051
rect 81445 176023 81479 176051
rect 81507 176023 81541 176051
rect 81569 176023 81603 176051
rect 81631 176023 96777 176051
rect 96805 176023 96839 176051
rect 96867 176023 96901 176051
rect 96929 176023 96963 176051
rect 96991 176023 112137 176051
rect 112165 176023 112199 176051
rect 112227 176023 112261 176051
rect 112289 176023 112323 176051
rect 112351 176023 127497 176051
rect 127525 176023 127559 176051
rect 127587 176023 127621 176051
rect 127649 176023 127683 176051
rect 127711 176023 142857 176051
rect 142885 176023 142919 176051
rect 142947 176023 142981 176051
rect 143009 176023 143043 176051
rect 143071 176023 158217 176051
rect 158245 176023 158279 176051
rect 158307 176023 158341 176051
rect 158369 176023 158403 176051
rect 158431 176023 173577 176051
rect 173605 176023 173639 176051
rect 173667 176023 173701 176051
rect 173729 176023 173763 176051
rect 173791 176023 188937 176051
rect 188965 176023 188999 176051
rect 189027 176023 189061 176051
rect 189089 176023 189123 176051
rect 189151 176023 204297 176051
rect 204325 176023 204359 176051
rect 204387 176023 204421 176051
rect 204449 176023 204483 176051
rect 204511 176023 219657 176051
rect 219685 176023 219719 176051
rect 219747 176023 219781 176051
rect 219809 176023 219843 176051
rect 219871 176023 235017 176051
rect 235045 176023 235079 176051
rect 235107 176023 235141 176051
rect 235169 176023 235203 176051
rect 235231 176023 250377 176051
rect 250405 176023 250439 176051
rect 250467 176023 250501 176051
rect 250529 176023 250563 176051
rect 250591 176023 265737 176051
rect 265765 176023 265799 176051
rect 265827 176023 265861 176051
rect 265889 176023 265923 176051
rect 265951 176023 281097 176051
rect 281125 176023 281159 176051
rect 281187 176023 281221 176051
rect 281249 176023 281283 176051
rect 281311 176023 296457 176051
rect 296485 176023 296519 176051
rect 296547 176023 296581 176051
rect 296609 176023 296643 176051
rect 296671 176023 298728 176051
rect 298756 176023 298790 176051
rect 298818 176023 298852 176051
rect 298880 176023 298914 176051
rect 298942 176023 298990 176051
rect -958 175989 298990 176023
rect -958 175961 -910 175989
rect -882 175961 -848 175989
rect -820 175961 -786 175989
rect -758 175961 -724 175989
rect -696 175961 4617 175989
rect 4645 175961 4679 175989
rect 4707 175961 4741 175989
rect 4769 175961 4803 175989
rect 4831 175961 19977 175989
rect 20005 175961 20039 175989
rect 20067 175961 20101 175989
rect 20129 175961 20163 175989
rect 20191 175961 35337 175989
rect 35365 175961 35399 175989
rect 35427 175961 35461 175989
rect 35489 175961 35523 175989
rect 35551 175961 50697 175989
rect 50725 175961 50759 175989
rect 50787 175961 50821 175989
rect 50849 175961 50883 175989
rect 50911 175961 66057 175989
rect 66085 175961 66119 175989
rect 66147 175961 66181 175989
rect 66209 175961 66243 175989
rect 66271 175961 81417 175989
rect 81445 175961 81479 175989
rect 81507 175961 81541 175989
rect 81569 175961 81603 175989
rect 81631 175961 96777 175989
rect 96805 175961 96839 175989
rect 96867 175961 96901 175989
rect 96929 175961 96963 175989
rect 96991 175961 112137 175989
rect 112165 175961 112199 175989
rect 112227 175961 112261 175989
rect 112289 175961 112323 175989
rect 112351 175961 127497 175989
rect 127525 175961 127559 175989
rect 127587 175961 127621 175989
rect 127649 175961 127683 175989
rect 127711 175961 142857 175989
rect 142885 175961 142919 175989
rect 142947 175961 142981 175989
rect 143009 175961 143043 175989
rect 143071 175961 158217 175989
rect 158245 175961 158279 175989
rect 158307 175961 158341 175989
rect 158369 175961 158403 175989
rect 158431 175961 173577 175989
rect 173605 175961 173639 175989
rect 173667 175961 173701 175989
rect 173729 175961 173763 175989
rect 173791 175961 188937 175989
rect 188965 175961 188999 175989
rect 189027 175961 189061 175989
rect 189089 175961 189123 175989
rect 189151 175961 204297 175989
rect 204325 175961 204359 175989
rect 204387 175961 204421 175989
rect 204449 175961 204483 175989
rect 204511 175961 219657 175989
rect 219685 175961 219719 175989
rect 219747 175961 219781 175989
rect 219809 175961 219843 175989
rect 219871 175961 235017 175989
rect 235045 175961 235079 175989
rect 235107 175961 235141 175989
rect 235169 175961 235203 175989
rect 235231 175961 250377 175989
rect 250405 175961 250439 175989
rect 250467 175961 250501 175989
rect 250529 175961 250563 175989
rect 250591 175961 265737 175989
rect 265765 175961 265799 175989
rect 265827 175961 265861 175989
rect 265889 175961 265923 175989
rect 265951 175961 281097 175989
rect 281125 175961 281159 175989
rect 281187 175961 281221 175989
rect 281249 175961 281283 175989
rect 281311 175961 296457 175989
rect 296485 175961 296519 175989
rect 296547 175961 296581 175989
rect 296609 175961 296643 175989
rect 296671 175961 298728 175989
rect 298756 175961 298790 175989
rect 298818 175961 298852 175989
rect 298880 175961 298914 175989
rect 298942 175961 298990 175989
rect -958 175913 298990 175961
rect -958 173175 298990 173223
rect -958 173147 -430 173175
rect -402 173147 -368 173175
rect -340 173147 -306 173175
rect -278 173147 -244 173175
rect -216 173147 2757 173175
rect 2785 173147 2819 173175
rect 2847 173147 2881 173175
rect 2909 173147 2943 173175
rect 2971 173147 8259 173175
rect 8287 173147 8321 173175
rect 8349 173147 18117 173175
rect 18145 173147 18179 173175
rect 18207 173147 18241 173175
rect 18269 173147 18303 173175
rect 18331 173147 23619 173175
rect 23647 173147 23681 173175
rect 23709 173147 33477 173175
rect 33505 173147 33539 173175
rect 33567 173147 33601 173175
rect 33629 173147 33663 173175
rect 33691 173147 38979 173175
rect 39007 173147 39041 173175
rect 39069 173147 48837 173175
rect 48865 173147 48899 173175
rect 48927 173147 48961 173175
rect 48989 173147 49023 173175
rect 49051 173147 54339 173175
rect 54367 173147 54401 173175
rect 54429 173147 64197 173175
rect 64225 173147 64259 173175
rect 64287 173147 64321 173175
rect 64349 173147 64383 173175
rect 64411 173147 69699 173175
rect 69727 173147 69761 173175
rect 69789 173147 79557 173175
rect 79585 173147 79619 173175
rect 79647 173147 79681 173175
rect 79709 173147 79743 173175
rect 79771 173147 85059 173175
rect 85087 173147 85121 173175
rect 85149 173147 94917 173175
rect 94945 173147 94979 173175
rect 95007 173147 95041 173175
rect 95069 173147 95103 173175
rect 95131 173147 100419 173175
rect 100447 173147 100481 173175
rect 100509 173147 110277 173175
rect 110305 173147 110339 173175
rect 110367 173147 110401 173175
rect 110429 173147 110463 173175
rect 110491 173147 115779 173175
rect 115807 173147 115841 173175
rect 115869 173147 125637 173175
rect 125665 173147 125699 173175
rect 125727 173147 125761 173175
rect 125789 173147 125823 173175
rect 125851 173147 131139 173175
rect 131167 173147 131201 173175
rect 131229 173147 140997 173175
rect 141025 173147 141059 173175
rect 141087 173147 141121 173175
rect 141149 173147 141183 173175
rect 141211 173147 146499 173175
rect 146527 173147 146561 173175
rect 146589 173147 156357 173175
rect 156385 173147 156419 173175
rect 156447 173147 156481 173175
rect 156509 173147 156543 173175
rect 156571 173147 161859 173175
rect 161887 173147 161921 173175
rect 161949 173147 171717 173175
rect 171745 173147 171779 173175
rect 171807 173147 171841 173175
rect 171869 173147 171903 173175
rect 171931 173147 177219 173175
rect 177247 173147 177281 173175
rect 177309 173147 187077 173175
rect 187105 173147 187139 173175
rect 187167 173147 187201 173175
rect 187229 173147 187263 173175
rect 187291 173147 192579 173175
rect 192607 173147 192641 173175
rect 192669 173147 202437 173175
rect 202465 173147 202499 173175
rect 202527 173147 202561 173175
rect 202589 173147 202623 173175
rect 202651 173147 207939 173175
rect 207967 173147 208001 173175
rect 208029 173147 217797 173175
rect 217825 173147 217859 173175
rect 217887 173147 217921 173175
rect 217949 173147 217983 173175
rect 218011 173147 223299 173175
rect 223327 173147 223361 173175
rect 223389 173147 233157 173175
rect 233185 173147 233219 173175
rect 233247 173147 233281 173175
rect 233309 173147 233343 173175
rect 233371 173147 238659 173175
rect 238687 173147 238721 173175
rect 238749 173147 248517 173175
rect 248545 173147 248579 173175
rect 248607 173147 248641 173175
rect 248669 173147 248703 173175
rect 248731 173147 254019 173175
rect 254047 173147 254081 173175
rect 254109 173147 263877 173175
rect 263905 173147 263939 173175
rect 263967 173147 264001 173175
rect 264029 173147 264063 173175
rect 264091 173147 269379 173175
rect 269407 173147 269441 173175
rect 269469 173147 279237 173175
rect 279265 173147 279299 173175
rect 279327 173147 279361 173175
rect 279389 173147 279423 173175
rect 279451 173147 284739 173175
rect 284767 173147 284801 173175
rect 284829 173147 294597 173175
rect 294625 173147 294659 173175
rect 294687 173147 294721 173175
rect 294749 173147 294783 173175
rect 294811 173147 298248 173175
rect 298276 173147 298310 173175
rect 298338 173147 298372 173175
rect 298400 173147 298434 173175
rect 298462 173147 298990 173175
rect -958 173113 298990 173147
rect -958 173085 -430 173113
rect -402 173085 -368 173113
rect -340 173085 -306 173113
rect -278 173085 -244 173113
rect -216 173085 2757 173113
rect 2785 173085 2819 173113
rect 2847 173085 2881 173113
rect 2909 173085 2943 173113
rect 2971 173085 8259 173113
rect 8287 173085 8321 173113
rect 8349 173085 18117 173113
rect 18145 173085 18179 173113
rect 18207 173085 18241 173113
rect 18269 173085 18303 173113
rect 18331 173085 23619 173113
rect 23647 173085 23681 173113
rect 23709 173085 33477 173113
rect 33505 173085 33539 173113
rect 33567 173085 33601 173113
rect 33629 173085 33663 173113
rect 33691 173085 38979 173113
rect 39007 173085 39041 173113
rect 39069 173085 48837 173113
rect 48865 173085 48899 173113
rect 48927 173085 48961 173113
rect 48989 173085 49023 173113
rect 49051 173085 54339 173113
rect 54367 173085 54401 173113
rect 54429 173085 64197 173113
rect 64225 173085 64259 173113
rect 64287 173085 64321 173113
rect 64349 173085 64383 173113
rect 64411 173085 69699 173113
rect 69727 173085 69761 173113
rect 69789 173085 79557 173113
rect 79585 173085 79619 173113
rect 79647 173085 79681 173113
rect 79709 173085 79743 173113
rect 79771 173085 85059 173113
rect 85087 173085 85121 173113
rect 85149 173085 94917 173113
rect 94945 173085 94979 173113
rect 95007 173085 95041 173113
rect 95069 173085 95103 173113
rect 95131 173085 100419 173113
rect 100447 173085 100481 173113
rect 100509 173085 110277 173113
rect 110305 173085 110339 173113
rect 110367 173085 110401 173113
rect 110429 173085 110463 173113
rect 110491 173085 115779 173113
rect 115807 173085 115841 173113
rect 115869 173085 125637 173113
rect 125665 173085 125699 173113
rect 125727 173085 125761 173113
rect 125789 173085 125823 173113
rect 125851 173085 131139 173113
rect 131167 173085 131201 173113
rect 131229 173085 140997 173113
rect 141025 173085 141059 173113
rect 141087 173085 141121 173113
rect 141149 173085 141183 173113
rect 141211 173085 146499 173113
rect 146527 173085 146561 173113
rect 146589 173085 156357 173113
rect 156385 173085 156419 173113
rect 156447 173085 156481 173113
rect 156509 173085 156543 173113
rect 156571 173085 161859 173113
rect 161887 173085 161921 173113
rect 161949 173085 171717 173113
rect 171745 173085 171779 173113
rect 171807 173085 171841 173113
rect 171869 173085 171903 173113
rect 171931 173085 177219 173113
rect 177247 173085 177281 173113
rect 177309 173085 187077 173113
rect 187105 173085 187139 173113
rect 187167 173085 187201 173113
rect 187229 173085 187263 173113
rect 187291 173085 192579 173113
rect 192607 173085 192641 173113
rect 192669 173085 202437 173113
rect 202465 173085 202499 173113
rect 202527 173085 202561 173113
rect 202589 173085 202623 173113
rect 202651 173085 207939 173113
rect 207967 173085 208001 173113
rect 208029 173085 217797 173113
rect 217825 173085 217859 173113
rect 217887 173085 217921 173113
rect 217949 173085 217983 173113
rect 218011 173085 223299 173113
rect 223327 173085 223361 173113
rect 223389 173085 233157 173113
rect 233185 173085 233219 173113
rect 233247 173085 233281 173113
rect 233309 173085 233343 173113
rect 233371 173085 238659 173113
rect 238687 173085 238721 173113
rect 238749 173085 248517 173113
rect 248545 173085 248579 173113
rect 248607 173085 248641 173113
rect 248669 173085 248703 173113
rect 248731 173085 254019 173113
rect 254047 173085 254081 173113
rect 254109 173085 263877 173113
rect 263905 173085 263939 173113
rect 263967 173085 264001 173113
rect 264029 173085 264063 173113
rect 264091 173085 269379 173113
rect 269407 173085 269441 173113
rect 269469 173085 279237 173113
rect 279265 173085 279299 173113
rect 279327 173085 279361 173113
rect 279389 173085 279423 173113
rect 279451 173085 284739 173113
rect 284767 173085 284801 173113
rect 284829 173085 294597 173113
rect 294625 173085 294659 173113
rect 294687 173085 294721 173113
rect 294749 173085 294783 173113
rect 294811 173085 298248 173113
rect 298276 173085 298310 173113
rect 298338 173085 298372 173113
rect 298400 173085 298434 173113
rect 298462 173085 298990 173113
rect -958 173051 298990 173085
rect -958 173023 -430 173051
rect -402 173023 -368 173051
rect -340 173023 -306 173051
rect -278 173023 -244 173051
rect -216 173023 2757 173051
rect 2785 173023 2819 173051
rect 2847 173023 2881 173051
rect 2909 173023 2943 173051
rect 2971 173023 8259 173051
rect 8287 173023 8321 173051
rect 8349 173023 18117 173051
rect 18145 173023 18179 173051
rect 18207 173023 18241 173051
rect 18269 173023 18303 173051
rect 18331 173023 23619 173051
rect 23647 173023 23681 173051
rect 23709 173023 33477 173051
rect 33505 173023 33539 173051
rect 33567 173023 33601 173051
rect 33629 173023 33663 173051
rect 33691 173023 38979 173051
rect 39007 173023 39041 173051
rect 39069 173023 48837 173051
rect 48865 173023 48899 173051
rect 48927 173023 48961 173051
rect 48989 173023 49023 173051
rect 49051 173023 54339 173051
rect 54367 173023 54401 173051
rect 54429 173023 64197 173051
rect 64225 173023 64259 173051
rect 64287 173023 64321 173051
rect 64349 173023 64383 173051
rect 64411 173023 69699 173051
rect 69727 173023 69761 173051
rect 69789 173023 79557 173051
rect 79585 173023 79619 173051
rect 79647 173023 79681 173051
rect 79709 173023 79743 173051
rect 79771 173023 85059 173051
rect 85087 173023 85121 173051
rect 85149 173023 94917 173051
rect 94945 173023 94979 173051
rect 95007 173023 95041 173051
rect 95069 173023 95103 173051
rect 95131 173023 100419 173051
rect 100447 173023 100481 173051
rect 100509 173023 110277 173051
rect 110305 173023 110339 173051
rect 110367 173023 110401 173051
rect 110429 173023 110463 173051
rect 110491 173023 115779 173051
rect 115807 173023 115841 173051
rect 115869 173023 125637 173051
rect 125665 173023 125699 173051
rect 125727 173023 125761 173051
rect 125789 173023 125823 173051
rect 125851 173023 131139 173051
rect 131167 173023 131201 173051
rect 131229 173023 140997 173051
rect 141025 173023 141059 173051
rect 141087 173023 141121 173051
rect 141149 173023 141183 173051
rect 141211 173023 146499 173051
rect 146527 173023 146561 173051
rect 146589 173023 156357 173051
rect 156385 173023 156419 173051
rect 156447 173023 156481 173051
rect 156509 173023 156543 173051
rect 156571 173023 161859 173051
rect 161887 173023 161921 173051
rect 161949 173023 171717 173051
rect 171745 173023 171779 173051
rect 171807 173023 171841 173051
rect 171869 173023 171903 173051
rect 171931 173023 177219 173051
rect 177247 173023 177281 173051
rect 177309 173023 187077 173051
rect 187105 173023 187139 173051
rect 187167 173023 187201 173051
rect 187229 173023 187263 173051
rect 187291 173023 192579 173051
rect 192607 173023 192641 173051
rect 192669 173023 202437 173051
rect 202465 173023 202499 173051
rect 202527 173023 202561 173051
rect 202589 173023 202623 173051
rect 202651 173023 207939 173051
rect 207967 173023 208001 173051
rect 208029 173023 217797 173051
rect 217825 173023 217859 173051
rect 217887 173023 217921 173051
rect 217949 173023 217983 173051
rect 218011 173023 223299 173051
rect 223327 173023 223361 173051
rect 223389 173023 233157 173051
rect 233185 173023 233219 173051
rect 233247 173023 233281 173051
rect 233309 173023 233343 173051
rect 233371 173023 238659 173051
rect 238687 173023 238721 173051
rect 238749 173023 248517 173051
rect 248545 173023 248579 173051
rect 248607 173023 248641 173051
rect 248669 173023 248703 173051
rect 248731 173023 254019 173051
rect 254047 173023 254081 173051
rect 254109 173023 263877 173051
rect 263905 173023 263939 173051
rect 263967 173023 264001 173051
rect 264029 173023 264063 173051
rect 264091 173023 269379 173051
rect 269407 173023 269441 173051
rect 269469 173023 279237 173051
rect 279265 173023 279299 173051
rect 279327 173023 279361 173051
rect 279389 173023 279423 173051
rect 279451 173023 284739 173051
rect 284767 173023 284801 173051
rect 284829 173023 294597 173051
rect 294625 173023 294659 173051
rect 294687 173023 294721 173051
rect 294749 173023 294783 173051
rect 294811 173023 298248 173051
rect 298276 173023 298310 173051
rect 298338 173023 298372 173051
rect 298400 173023 298434 173051
rect 298462 173023 298990 173051
rect -958 172989 298990 173023
rect -958 172961 -430 172989
rect -402 172961 -368 172989
rect -340 172961 -306 172989
rect -278 172961 -244 172989
rect -216 172961 2757 172989
rect 2785 172961 2819 172989
rect 2847 172961 2881 172989
rect 2909 172961 2943 172989
rect 2971 172961 8259 172989
rect 8287 172961 8321 172989
rect 8349 172961 18117 172989
rect 18145 172961 18179 172989
rect 18207 172961 18241 172989
rect 18269 172961 18303 172989
rect 18331 172961 23619 172989
rect 23647 172961 23681 172989
rect 23709 172961 33477 172989
rect 33505 172961 33539 172989
rect 33567 172961 33601 172989
rect 33629 172961 33663 172989
rect 33691 172961 38979 172989
rect 39007 172961 39041 172989
rect 39069 172961 48837 172989
rect 48865 172961 48899 172989
rect 48927 172961 48961 172989
rect 48989 172961 49023 172989
rect 49051 172961 54339 172989
rect 54367 172961 54401 172989
rect 54429 172961 64197 172989
rect 64225 172961 64259 172989
rect 64287 172961 64321 172989
rect 64349 172961 64383 172989
rect 64411 172961 69699 172989
rect 69727 172961 69761 172989
rect 69789 172961 79557 172989
rect 79585 172961 79619 172989
rect 79647 172961 79681 172989
rect 79709 172961 79743 172989
rect 79771 172961 85059 172989
rect 85087 172961 85121 172989
rect 85149 172961 94917 172989
rect 94945 172961 94979 172989
rect 95007 172961 95041 172989
rect 95069 172961 95103 172989
rect 95131 172961 100419 172989
rect 100447 172961 100481 172989
rect 100509 172961 110277 172989
rect 110305 172961 110339 172989
rect 110367 172961 110401 172989
rect 110429 172961 110463 172989
rect 110491 172961 115779 172989
rect 115807 172961 115841 172989
rect 115869 172961 125637 172989
rect 125665 172961 125699 172989
rect 125727 172961 125761 172989
rect 125789 172961 125823 172989
rect 125851 172961 131139 172989
rect 131167 172961 131201 172989
rect 131229 172961 140997 172989
rect 141025 172961 141059 172989
rect 141087 172961 141121 172989
rect 141149 172961 141183 172989
rect 141211 172961 146499 172989
rect 146527 172961 146561 172989
rect 146589 172961 156357 172989
rect 156385 172961 156419 172989
rect 156447 172961 156481 172989
rect 156509 172961 156543 172989
rect 156571 172961 161859 172989
rect 161887 172961 161921 172989
rect 161949 172961 171717 172989
rect 171745 172961 171779 172989
rect 171807 172961 171841 172989
rect 171869 172961 171903 172989
rect 171931 172961 177219 172989
rect 177247 172961 177281 172989
rect 177309 172961 187077 172989
rect 187105 172961 187139 172989
rect 187167 172961 187201 172989
rect 187229 172961 187263 172989
rect 187291 172961 192579 172989
rect 192607 172961 192641 172989
rect 192669 172961 202437 172989
rect 202465 172961 202499 172989
rect 202527 172961 202561 172989
rect 202589 172961 202623 172989
rect 202651 172961 207939 172989
rect 207967 172961 208001 172989
rect 208029 172961 217797 172989
rect 217825 172961 217859 172989
rect 217887 172961 217921 172989
rect 217949 172961 217983 172989
rect 218011 172961 223299 172989
rect 223327 172961 223361 172989
rect 223389 172961 233157 172989
rect 233185 172961 233219 172989
rect 233247 172961 233281 172989
rect 233309 172961 233343 172989
rect 233371 172961 238659 172989
rect 238687 172961 238721 172989
rect 238749 172961 248517 172989
rect 248545 172961 248579 172989
rect 248607 172961 248641 172989
rect 248669 172961 248703 172989
rect 248731 172961 254019 172989
rect 254047 172961 254081 172989
rect 254109 172961 263877 172989
rect 263905 172961 263939 172989
rect 263967 172961 264001 172989
rect 264029 172961 264063 172989
rect 264091 172961 269379 172989
rect 269407 172961 269441 172989
rect 269469 172961 279237 172989
rect 279265 172961 279299 172989
rect 279327 172961 279361 172989
rect 279389 172961 279423 172989
rect 279451 172961 284739 172989
rect 284767 172961 284801 172989
rect 284829 172961 294597 172989
rect 294625 172961 294659 172989
rect 294687 172961 294721 172989
rect 294749 172961 294783 172989
rect 294811 172961 298248 172989
rect 298276 172961 298310 172989
rect 298338 172961 298372 172989
rect 298400 172961 298434 172989
rect 298462 172961 298990 172989
rect -958 172913 298990 172961
rect -958 167175 298990 167223
rect -958 167147 -910 167175
rect -882 167147 -848 167175
rect -820 167147 -786 167175
rect -758 167147 -724 167175
rect -696 167147 4617 167175
rect 4645 167147 4679 167175
rect 4707 167147 4741 167175
rect 4769 167147 4803 167175
rect 4831 167147 15939 167175
rect 15967 167147 16001 167175
rect 16029 167147 19977 167175
rect 20005 167147 20039 167175
rect 20067 167147 20101 167175
rect 20129 167147 20163 167175
rect 20191 167147 31299 167175
rect 31327 167147 31361 167175
rect 31389 167147 35337 167175
rect 35365 167147 35399 167175
rect 35427 167147 35461 167175
rect 35489 167147 35523 167175
rect 35551 167147 46659 167175
rect 46687 167147 46721 167175
rect 46749 167147 50697 167175
rect 50725 167147 50759 167175
rect 50787 167147 50821 167175
rect 50849 167147 50883 167175
rect 50911 167147 62019 167175
rect 62047 167147 62081 167175
rect 62109 167147 66057 167175
rect 66085 167147 66119 167175
rect 66147 167147 66181 167175
rect 66209 167147 66243 167175
rect 66271 167147 77379 167175
rect 77407 167147 77441 167175
rect 77469 167147 81417 167175
rect 81445 167147 81479 167175
rect 81507 167147 81541 167175
rect 81569 167147 81603 167175
rect 81631 167147 92739 167175
rect 92767 167147 92801 167175
rect 92829 167147 96777 167175
rect 96805 167147 96839 167175
rect 96867 167147 96901 167175
rect 96929 167147 96963 167175
rect 96991 167147 108099 167175
rect 108127 167147 108161 167175
rect 108189 167147 112137 167175
rect 112165 167147 112199 167175
rect 112227 167147 112261 167175
rect 112289 167147 112323 167175
rect 112351 167147 123459 167175
rect 123487 167147 123521 167175
rect 123549 167147 127497 167175
rect 127525 167147 127559 167175
rect 127587 167147 127621 167175
rect 127649 167147 127683 167175
rect 127711 167147 138819 167175
rect 138847 167147 138881 167175
rect 138909 167147 142857 167175
rect 142885 167147 142919 167175
rect 142947 167147 142981 167175
rect 143009 167147 143043 167175
rect 143071 167147 154179 167175
rect 154207 167147 154241 167175
rect 154269 167147 158217 167175
rect 158245 167147 158279 167175
rect 158307 167147 158341 167175
rect 158369 167147 158403 167175
rect 158431 167147 169539 167175
rect 169567 167147 169601 167175
rect 169629 167147 173577 167175
rect 173605 167147 173639 167175
rect 173667 167147 173701 167175
rect 173729 167147 173763 167175
rect 173791 167147 184899 167175
rect 184927 167147 184961 167175
rect 184989 167147 188937 167175
rect 188965 167147 188999 167175
rect 189027 167147 189061 167175
rect 189089 167147 189123 167175
rect 189151 167147 200259 167175
rect 200287 167147 200321 167175
rect 200349 167147 204297 167175
rect 204325 167147 204359 167175
rect 204387 167147 204421 167175
rect 204449 167147 204483 167175
rect 204511 167147 215619 167175
rect 215647 167147 215681 167175
rect 215709 167147 219657 167175
rect 219685 167147 219719 167175
rect 219747 167147 219781 167175
rect 219809 167147 219843 167175
rect 219871 167147 230979 167175
rect 231007 167147 231041 167175
rect 231069 167147 235017 167175
rect 235045 167147 235079 167175
rect 235107 167147 235141 167175
rect 235169 167147 235203 167175
rect 235231 167147 246339 167175
rect 246367 167147 246401 167175
rect 246429 167147 250377 167175
rect 250405 167147 250439 167175
rect 250467 167147 250501 167175
rect 250529 167147 250563 167175
rect 250591 167147 261699 167175
rect 261727 167147 261761 167175
rect 261789 167147 265737 167175
rect 265765 167147 265799 167175
rect 265827 167147 265861 167175
rect 265889 167147 265923 167175
rect 265951 167147 277059 167175
rect 277087 167147 277121 167175
rect 277149 167147 281097 167175
rect 281125 167147 281159 167175
rect 281187 167147 281221 167175
rect 281249 167147 281283 167175
rect 281311 167147 296457 167175
rect 296485 167147 296519 167175
rect 296547 167147 296581 167175
rect 296609 167147 296643 167175
rect 296671 167147 298728 167175
rect 298756 167147 298790 167175
rect 298818 167147 298852 167175
rect 298880 167147 298914 167175
rect 298942 167147 298990 167175
rect -958 167113 298990 167147
rect -958 167085 -910 167113
rect -882 167085 -848 167113
rect -820 167085 -786 167113
rect -758 167085 -724 167113
rect -696 167085 4617 167113
rect 4645 167085 4679 167113
rect 4707 167085 4741 167113
rect 4769 167085 4803 167113
rect 4831 167085 15939 167113
rect 15967 167085 16001 167113
rect 16029 167085 19977 167113
rect 20005 167085 20039 167113
rect 20067 167085 20101 167113
rect 20129 167085 20163 167113
rect 20191 167085 31299 167113
rect 31327 167085 31361 167113
rect 31389 167085 35337 167113
rect 35365 167085 35399 167113
rect 35427 167085 35461 167113
rect 35489 167085 35523 167113
rect 35551 167085 46659 167113
rect 46687 167085 46721 167113
rect 46749 167085 50697 167113
rect 50725 167085 50759 167113
rect 50787 167085 50821 167113
rect 50849 167085 50883 167113
rect 50911 167085 62019 167113
rect 62047 167085 62081 167113
rect 62109 167085 66057 167113
rect 66085 167085 66119 167113
rect 66147 167085 66181 167113
rect 66209 167085 66243 167113
rect 66271 167085 77379 167113
rect 77407 167085 77441 167113
rect 77469 167085 81417 167113
rect 81445 167085 81479 167113
rect 81507 167085 81541 167113
rect 81569 167085 81603 167113
rect 81631 167085 92739 167113
rect 92767 167085 92801 167113
rect 92829 167085 96777 167113
rect 96805 167085 96839 167113
rect 96867 167085 96901 167113
rect 96929 167085 96963 167113
rect 96991 167085 108099 167113
rect 108127 167085 108161 167113
rect 108189 167085 112137 167113
rect 112165 167085 112199 167113
rect 112227 167085 112261 167113
rect 112289 167085 112323 167113
rect 112351 167085 123459 167113
rect 123487 167085 123521 167113
rect 123549 167085 127497 167113
rect 127525 167085 127559 167113
rect 127587 167085 127621 167113
rect 127649 167085 127683 167113
rect 127711 167085 138819 167113
rect 138847 167085 138881 167113
rect 138909 167085 142857 167113
rect 142885 167085 142919 167113
rect 142947 167085 142981 167113
rect 143009 167085 143043 167113
rect 143071 167085 154179 167113
rect 154207 167085 154241 167113
rect 154269 167085 158217 167113
rect 158245 167085 158279 167113
rect 158307 167085 158341 167113
rect 158369 167085 158403 167113
rect 158431 167085 169539 167113
rect 169567 167085 169601 167113
rect 169629 167085 173577 167113
rect 173605 167085 173639 167113
rect 173667 167085 173701 167113
rect 173729 167085 173763 167113
rect 173791 167085 184899 167113
rect 184927 167085 184961 167113
rect 184989 167085 188937 167113
rect 188965 167085 188999 167113
rect 189027 167085 189061 167113
rect 189089 167085 189123 167113
rect 189151 167085 200259 167113
rect 200287 167085 200321 167113
rect 200349 167085 204297 167113
rect 204325 167085 204359 167113
rect 204387 167085 204421 167113
rect 204449 167085 204483 167113
rect 204511 167085 215619 167113
rect 215647 167085 215681 167113
rect 215709 167085 219657 167113
rect 219685 167085 219719 167113
rect 219747 167085 219781 167113
rect 219809 167085 219843 167113
rect 219871 167085 230979 167113
rect 231007 167085 231041 167113
rect 231069 167085 235017 167113
rect 235045 167085 235079 167113
rect 235107 167085 235141 167113
rect 235169 167085 235203 167113
rect 235231 167085 246339 167113
rect 246367 167085 246401 167113
rect 246429 167085 250377 167113
rect 250405 167085 250439 167113
rect 250467 167085 250501 167113
rect 250529 167085 250563 167113
rect 250591 167085 261699 167113
rect 261727 167085 261761 167113
rect 261789 167085 265737 167113
rect 265765 167085 265799 167113
rect 265827 167085 265861 167113
rect 265889 167085 265923 167113
rect 265951 167085 277059 167113
rect 277087 167085 277121 167113
rect 277149 167085 281097 167113
rect 281125 167085 281159 167113
rect 281187 167085 281221 167113
rect 281249 167085 281283 167113
rect 281311 167085 296457 167113
rect 296485 167085 296519 167113
rect 296547 167085 296581 167113
rect 296609 167085 296643 167113
rect 296671 167085 298728 167113
rect 298756 167085 298790 167113
rect 298818 167085 298852 167113
rect 298880 167085 298914 167113
rect 298942 167085 298990 167113
rect -958 167051 298990 167085
rect -958 167023 -910 167051
rect -882 167023 -848 167051
rect -820 167023 -786 167051
rect -758 167023 -724 167051
rect -696 167023 4617 167051
rect 4645 167023 4679 167051
rect 4707 167023 4741 167051
rect 4769 167023 4803 167051
rect 4831 167023 15939 167051
rect 15967 167023 16001 167051
rect 16029 167023 19977 167051
rect 20005 167023 20039 167051
rect 20067 167023 20101 167051
rect 20129 167023 20163 167051
rect 20191 167023 31299 167051
rect 31327 167023 31361 167051
rect 31389 167023 35337 167051
rect 35365 167023 35399 167051
rect 35427 167023 35461 167051
rect 35489 167023 35523 167051
rect 35551 167023 46659 167051
rect 46687 167023 46721 167051
rect 46749 167023 50697 167051
rect 50725 167023 50759 167051
rect 50787 167023 50821 167051
rect 50849 167023 50883 167051
rect 50911 167023 62019 167051
rect 62047 167023 62081 167051
rect 62109 167023 66057 167051
rect 66085 167023 66119 167051
rect 66147 167023 66181 167051
rect 66209 167023 66243 167051
rect 66271 167023 77379 167051
rect 77407 167023 77441 167051
rect 77469 167023 81417 167051
rect 81445 167023 81479 167051
rect 81507 167023 81541 167051
rect 81569 167023 81603 167051
rect 81631 167023 92739 167051
rect 92767 167023 92801 167051
rect 92829 167023 96777 167051
rect 96805 167023 96839 167051
rect 96867 167023 96901 167051
rect 96929 167023 96963 167051
rect 96991 167023 108099 167051
rect 108127 167023 108161 167051
rect 108189 167023 112137 167051
rect 112165 167023 112199 167051
rect 112227 167023 112261 167051
rect 112289 167023 112323 167051
rect 112351 167023 123459 167051
rect 123487 167023 123521 167051
rect 123549 167023 127497 167051
rect 127525 167023 127559 167051
rect 127587 167023 127621 167051
rect 127649 167023 127683 167051
rect 127711 167023 138819 167051
rect 138847 167023 138881 167051
rect 138909 167023 142857 167051
rect 142885 167023 142919 167051
rect 142947 167023 142981 167051
rect 143009 167023 143043 167051
rect 143071 167023 154179 167051
rect 154207 167023 154241 167051
rect 154269 167023 158217 167051
rect 158245 167023 158279 167051
rect 158307 167023 158341 167051
rect 158369 167023 158403 167051
rect 158431 167023 169539 167051
rect 169567 167023 169601 167051
rect 169629 167023 173577 167051
rect 173605 167023 173639 167051
rect 173667 167023 173701 167051
rect 173729 167023 173763 167051
rect 173791 167023 184899 167051
rect 184927 167023 184961 167051
rect 184989 167023 188937 167051
rect 188965 167023 188999 167051
rect 189027 167023 189061 167051
rect 189089 167023 189123 167051
rect 189151 167023 200259 167051
rect 200287 167023 200321 167051
rect 200349 167023 204297 167051
rect 204325 167023 204359 167051
rect 204387 167023 204421 167051
rect 204449 167023 204483 167051
rect 204511 167023 215619 167051
rect 215647 167023 215681 167051
rect 215709 167023 219657 167051
rect 219685 167023 219719 167051
rect 219747 167023 219781 167051
rect 219809 167023 219843 167051
rect 219871 167023 230979 167051
rect 231007 167023 231041 167051
rect 231069 167023 235017 167051
rect 235045 167023 235079 167051
rect 235107 167023 235141 167051
rect 235169 167023 235203 167051
rect 235231 167023 246339 167051
rect 246367 167023 246401 167051
rect 246429 167023 250377 167051
rect 250405 167023 250439 167051
rect 250467 167023 250501 167051
rect 250529 167023 250563 167051
rect 250591 167023 261699 167051
rect 261727 167023 261761 167051
rect 261789 167023 265737 167051
rect 265765 167023 265799 167051
rect 265827 167023 265861 167051
rect 265889 167023 265923 167051
rect 265951 167023 277059 167051
rect 277087 167023 277121 167051
rect 277149 167023 281097 167051
rect 281125 167023 281159 167051
rect 281187 167023 281221 167051
rect 281249 167023 281283 167051
rect 281311 167023 296457 167051
rect 296485 167023 296519 167051
rect 296547 167023 296581 167051
rect 296609 167023 296643 167051
rect 296671 167023 298728 167051
rect 298756 167023 298790 167051
rect 298818 167023 298852 167051
rect 298880 167023 298914 167051
rect 298942 167023 298990 167051
rect -958 166989 298990 167023
rect -958 166961 -910 166989
rect -882 166961 -848 166989
rect -820 166961 -786 166989
rect -758 166961 -724 166989
rect -696 166961 4617 166989
rect 4645 166961 4679 166989
rect 4707 166961 4741 166989
rect 4769 166961 4803 166989
rect 4831 166961 15939 166989
rect 15967 166961 16001 166989
rect 16029 166961 19977 166989
rect 20005 166961 20039 166989
rect 20067 166961 20101 166989
rect 20129 166961 20163 166989
rect 20191 166961 31299 166989
rect 31327 166961 31361 166989
rect 31389 166961 35337 166989
rect 35365 166961 35399 166989
rect 35427 166961 35461 166989
rect 35489 166961 35523 166989
rect 35551 166961 46659 166989
rect 46687 166961 46721 166989
rect 46749 166961 50697 166989
rect 50725 166961 50759 166989
rect 50787 166961 50821 166989
rect 50849 166961 50883 166989
rect 50911 166961 62019 166989
rect 62047 166961 62081 166989
rect 62109 166961 66057 166989
rect 66085 166961 66119 166989
rect 66147 166961 66181 166989
rect 66209 166961 66243 166989
rect 66271 166961 77379 166989
rect 77407 166961 77441 166989
rect 77469 166961 81417 166989
rect 81445 166961 81479 166989
rect 81507 166961 81541 166989
rect 81569 166961 81603 166989
rect 81631 166961 92739 166989
rect 92767 166961 92801 166989
rect 92829 166961 96777 166989
rect 96805 166961 96839 166989
rect 96867 166961 96901 166989
rect 96929 166961 96963 166989
rect 96991 166961 108099 166989
rect 108127 166961 108161 166989
rect 108189 166961 112137 166989
rect 112165 166961 112199 166989
rect 112227 166961 112261 166989
rect 112289 166961 112323 166989
rect 112351 166961 123459 166989
rect 123487 166961 123521 166989
rect 123549 166961 127497 166989
rect 127525 166961 127559 166989
rect 127587 166961 127621 166989
rect 127649 166961 127683 166989
rect 127711 166961 138819 166989
rect 138847 166961 138881 166989
rect 138909 166961 142857 166989
rect 142885 166961 142919 166989
rect 142947 166961 142981 166989
rect 143009 166961 143043 166989
rect 143071 166961 154179 166989
rect 154207 166961 154241 166989
rect 154269 166961 158217 166989
rect 158245 166961 158279 166989
rect 158307 166961 158341 166989
rect 158369 166961 158403 166989
rect 158431 166961 169539 166989
rect 169567 166961 169601 166989
rect 169629 166961 173577 166989
rect 173605 166961 173639 166989
rect 173667 166961 173701 166989
rect 173729 166961 173763 166989
rect 173791 166961 184899 166989
rect 184927 166961 184961 166989
rect 184989 166961 188937 166989
rect 188965 166961 188999 166989
rect 189027 166961 189061 166989
rect 189089 166961 189123 166989
rect 189151 166961 200259 166989
rect 200287 166961 200321 166989
rect 200349 166961 204297 166989
rect 204325 166961 204359 166989
rect 204387 166961 204421 166989
rect 204449 166961 204483 166989
rect 204511 166961 215619 166989
rect 215647 166961 215681 166989
rect 215709 166961 219657 166989
rect 219685 166961 219719 166989
rect 219747 166961 219781 166989
rect 219809 166961 219843 166989
rect 219871 166961 230979 166989
rect 231007 166961 231041 166989
rect 231069 166961 235017 166989
rect 235045 166961 235079 166989
rect 235107 166961 235141 166989
rect 235169 166961 235203 166989
rect 235231 166961 246339 166989
rect 246367 166961 246401 166989
rect 246429 166961 250377 166989
rect 250405 166961 250439 166989
rect 250467 166961 250501 166989
rect 250529 166961 250563 166989
rect 250591 166961 261699 166989
rect 261727 166961 261761 166989
rect 261789 166961 265737 166989
rect 265765 166961 265799 166989
rect 265827 166961 265861 166989
rect 265889 166961 265923 166989
rect 265951 166961 277059 166989
rect 277087 166961 277121 166989
rect 277149 166961 281097 166989
rect 281125 166961 281159 166989
rect 281187 166961 281221 166989
rect 281249 166961 281283 166989
rect 281311 166961 296457 166989
rect 296485 166961 296519 166989
rect 296547 166961 296581 166989
rect 296609 166961 296643 166989
rect 296671 166961 298728 166989
rect 298756 166961 298790 166989
rect 298818 166961 298852 166989
rect 298880 166961 298914 166989
rect 298942 166961 298990 166989
rect -958 166913 298990 166961
rect -958 164175 298990 164223
rect -958 164147 -430 164175
rect -402 164147 -368 164175
rect -340 164147 -306 164175
rect -278 164147 -244 164175
rect -216 164147 2757 164175
rect 2785 164147 2819 164175
rect 2847 164147 2881 164175
rect 2909 164147 2943 164175
rect 2971 164147 8259 164175
rect 8287 164147 8321 164175
rect 8349 164147 18117 164175
rect 18145 164147 18179 164175
rect 18207 164147 18241 164175
rect 18269 164147 18303 164175
rect 18331 164147 23619 164175
rect 23647 164147 23681 164175
rect 23709 164147 33477 164175
rect 33505 164147 33539 164175
rect 33567 164147 33601 164175
rect 33629 164147 33663 164175
rect 33691 164147 38979 164175
rect 39007 164147 39041 164175
rect 39069 164147 48837 164175
rect 48865 164147 48899 164175
rect 48927 164147 48961 164175
rect 48989 164147 49023 164175
rect 49051 164147 54339 164175
rect 54367 164147 54401 164175
rect 54429 164147 64197 164175
rect 64225 164147 64259 164175
rect 64287 164147 64321 164175
rect 64349 164147 64383 164175
rect 64411 164147 69699 164175
rect 69727 164147 69761 164175
rect 69789 164147 79557 164175
rect 79585 164147 79619 164175
rect 79647 164147 79681 164175
rect 79709 164147 79743 164175
rect 79771 164147 85059 164175
rect 85087 164147 85121 164175
rect 85149 164147 94917 164175
rect 94945 164147 94979 164175
rect 95007 164147 95041 164175
rect 95069 164147 95103 164175
rect 95131 164147 100419 164175
rect 100447 164147 100481 164175
rect 100509 164147 110277 164175
rect 110305 164147 110339 164175
rect 110367 164147 110401 164175
rect 110429 164147 110463 164175
rect 110491 164147 115779 164175
rect 115807 164147 115841 164175
rect 115869 164147 125637 164175
rect 125665 164147 125699 164175
rect 125727 164147 125761 164175
rect 125789 164147 125823 164175
rect 125851 164147 131139 164175
rect 131167 164147 131201 164175
rect 131229 164147 140997 164175
rect 141025 164147 141059 164175
rect 141087 164147 141121 164175
rect 141149 164147 141183 164175
rect 141211 164147 146499 164175
rect 146527 164147 146561 164175
rect 146589 164147 156357 164175
rect 156385 164147 156419 164175
rect 156447 164147 156481 164175
rect 156509 164147 156543 164175
rect 156571 164147 161859 164175
rect 161887 164147 161921 164175
rect 161949 164147 171717 164175
rect 171745 164147 171779 164175
rect 171807 164147 171841 164175
rect 171869 164147 171903 164175
rect 171931 164147 177219 164175
rect 177247 164147 177281 164175
rect 177309 164147 187077 164175
rect 187105 164147 187139 164175
rect 187167 164147 187201 164175
rect 187229 164147 187263 164175
rect 187291 164147 192579 164175
rect 192607 164147 192641 164175
rect 192669 164147 202437 164175
rect 202465 164147 202499 164175
rect 202527 164147 202561 164175
rect 202589 164147 202623 164175
rect 202651 164147 207939 164175
rect 207967 164147 208001 164175
rect 208029 164147 217797 164175
rect 217825 164147 217859 164175
rect 217887 164147 217921 164175
rect 217949 164147 217983 164175
rect 218011 164147 223299 164175
rect 223327 164147 223361 164175
rect 223389 164147 233157 164175
rect 233185 164147 233219 164175
rect 233247 164147 233281 164175
rect 233309 164147 233343 164175
rect 233371 164147 238659 164175
rect 238687 164147 238721 164175
rect 238749 164147 248517 164175
rect 248545 164147 248579 164175
rect 248607 164147 248641 164175
rect 248669 164147 248703 164175
rect 248731 164147 254019 164175
rect 254047 164147 254081 164175
rect 254109 164147 263877 164175
rect 263905 164147 263939 164175
rect 263967 164147 264001 164175
rect 264029 164147 264063 164175
rect 264091 164147 269379 164175
rect 269407 164147 269441 164175
rect 269469 164147 279237 164175
rect 279265 164147 279299 164175
rect 279327 164147 279361 164175
rect 279389 164147 279423 164175
rect 279451 164147 284739 164175
rect 284767 164147 284801 164175
rect 284829 164147 294597 164175
rect 294625 164147 294659 164175
rect 294687 164147 294721 164175
rect 294749 164147 294783 164175
rect 294811 164147 298248 164175
rect 298276 164147 298310 164175
rect 298338 164147 298372 164175
rect 298400 164147 298434 164175
rect 298462 164147 298990 164175
rect -958 164113 298990 164147
rect -958 164085 -430 164113
rect -402 164085 -368 164113
rect -340 164085 -306 164113
rect -278 164085 -244 164113
rect -216 164085 2757 164113
rect 2785 164085 2819 164113
rect 2847 164085 2881 164113
rect 2909 164085 2943 164113
rect 2971 164085 8259 164113
rect 8287 164085 8321 164113
rect 8349 164085 18117 164113
rect 18145 164085 18179 164113
rect 18207 164085 18241 164113
rect 18269 164085 18303 164113
rect 18331 164085 23619 164113
rect 23647 164085 23681 164113
rect 23709 164085 33477 164113
rect 33505 164085 33539 164113
rect 33567 164085 33601 164113
rect 33629 164085 33663 164113
rect 33691 164085 38979 164113
rect 39007 164085 39041 164113
rect 39069 164085 48837 164113
rect 48865 164085 48899 164113
rect 48927 164085 48961 164113
rect 48989 164085 49023 164113
rect 49051 164085 54339 164113
rect 54367 164085 54401 164113
rect 54429 164085 64197 164113
rect 64225 164085 64259 164113
rect 64287 164085 64321 164113
rect 64349 164085 64383 164113
rect 64411 164085 69699 164113
rect 69727 164085 69761 164113
rect 69789 164085 79557 164113
rect 79585 164085 79619 164113
rect 79647 164085 79681 164113
rect 79709 164085 79743 164113
rect 79771 164085 85059 164113
rect 85087 164085 85121 164113
rect 85149 164085 94917 164113
rect 94945 164085 94979 164113
rect 95007 164085 95041 164113
rect 95069 164085 95103 164113
rect 95131 164085 100419 164113
rect 100447 164085 100481 164113
rect 100509 164085 110277 164113
rect 110305 164085 110339 164113
rect 110367 164085 110401 164113
rect 110429 164085 110463 164113
rect 110491 164085 115779 164113
rect 115807 164085 115841 164113
rect 115869 164085 125637 164113
rect 125665 164085 125699 164113
rect 125727 164085 125761 164113
rect 125789 164085 125823 164113
rect 125851 164085 131139 164113
rect 131167 164085 131201 164113
rect 131229 164085 140997 164113
rect 141025 164085 141059 164113
rect 141087 164085 141121 164113
rect 141149 164085 141183 164113
rect 141211 164085 146499 164113
rect 146527 164085 146561 164113
rect 146589 164085 156357 164113
rect 156385 164085 156419 164113
rect 156447 164085 156481 164113
rect 156509 164085 156543 164113
rect 156571 164085 161859 164113
rect 161887 164085 161921 164113
rect 161949 164085 171717 164113
rect 171745 164085 171779 164113
rect 171807 164085 171841 164113
rect 171869 164085 171903 164113
rect 171931 164085 177219 164113
rect 177247 164085 177281 164113
rect 177309 164085 187077 164113
rect 187105 164085 187139 164113
rect 187167 164085 187201 164113
rect 187229 164085 187263 164113
rect 187291 164085 192579 164113
rect 192607 164085 192641 164113
rect 192669 164085 202437 164113
rect 202465 164085 202499 164113
rect 202527 164085 202561 164113
rect 202589 164085 202623 164113
rect 202651 164085 207939 164113
rect 207967 164085 208001 164113
rect 208029 164085 217797 164113
rect 217825 164085 217859 164113
rect 217887 164085 217921 164113
rect 217949 164085 217983 164113
rect 218011 164085 223299 164113
rect 223327 164085 223361 164113
rect 223389 164085 233157 164113
rect 233185 164085 233219 164113
rect 233247 164085 233281 164113
rect 233309 164085 233343 164113
rect 233371 164085 238659 164113
rect 238687 164085 238721 164113
rect 238749 164085 248517 164113
rect 248545 164085 248579 164113
rect 248607 164085 248641 164113
rect 248669 164085 248703 164113
rect 248731 164085 254019 164113
rect 254047 164085 254081 164113
rect 254109 164085 263877 164113
rect 263905 164085 263939 164113
rect 263967 164085 264001 164113
rect 264029 164085 264063 164113
rect 264091 164085 269379 164113
rect 269407 164085 269441 164113
rect 269469 164085 279237 164113
rect 279265 164085 279299 164113
rect 279327 164085 279361 164113
rect 279389 164085 279423 164113
rect 279451 164085 284739 164113
rect 284767 164085 284801 164113
rect 284829 164085 294597 164113
rect 294625 164085 294659 164113
rect 294687 164085 294721 164113
rect 294749 164085 294783 164113
rect 294811 164085 298248 164113
rect 298276 164085 298310 164113
rect 298338 164085 298372 164113
rect 298400 164085 298434 164113
rect 298462 164085 298990 164113
rect -958 164051 298990 164085
rect -958 164023 -430 164051
rect -402 164023 -368 164051
rect -340 164023 -306 164051
rect -278 164023 -244 164051
rect -216 164023 2757 164051
rect 2785 164023 2819 164051
rect 2847 164023 2881 164051
rect 2909 164023 2943 164051
rect 2971 164023 8259 164051
rect 8287 164023 8321 164051
rect 8349 164023 18117 164051
rect 18145 164023 18179 164051
rect 18207 164023 18241 164051
rect 18269 164023 18303 164051
rect 18331 164023 23619 164051
rect 23647 164023 23681 164051
rect 23709 164023 33477 164051
rect 33505 164023 33539 164051
rect 33567 164023 33601 164051
rect 33629 164023 33663 164051
rect 33691 164023 38979 164051
rect 39007 164023 39041 164051
rect 39069 164023 48837 164051
rect 48865 164023 48899 164051
rect 48927 164023 48961 164051
rect 48989 164023 49023 164051
rect 49051 164023 54339 164051
rect 54367 164023 54401 164051
rect 54429 164023 64197 164051
rect 64225 164023 64259 164051
rect 64287 164023 64321 164051
rect 64349 164023 64383 164051
rect 64411 164023 69699 164051
rect 69727 164023 69761 164051
rect 69789 164023 79557 164051
rect 79585 164023 79619 164051
rect 79647 164023 79681 164051
rect 79709 164023 79743 164051
rect 79771 164023 85059 164051
rect 85087 164023 85121 164051
rect 85149 164023 94917 164051
rect 94945 164023 94979 164051
rect 95007 164023 95041 164051
rect 95069 164023 95103 164051
rect 95131 164023 100419 164051
rect 100447 164023 100481 164051
rect 100509 164023 110277 164051
rect 110305 164023 110339 164051
rect 110367 164023 110401 164051
rect 110429 164023 110463 164051
rect 110491 164023 115779 164051
rect 115807 164023 115841 164051
rect 115869 164023 125637 164051
rect 125665 164023 125699 164051
rect 125727 164023 125761 164051
rect 125789 164023 125823 164051
rect 125851 164023 131139 164051
rect 131167 164023 131201 164051
rect 131229 164023 140997 164051
rect 141025 164023 141059 164051
rect 141087 164023 141121 164051
rect 141149 164023 141183 164051
rect 141211 164023 146499 164051
rect 146527 164023 146561 164051
rect 146589 164023 156357 164051
rect 156385 164023 156419 164051
rect 156447 164023 156481 164051
rect 156509 164023 156543 164051
rect 156571 164023 161859 164051
rect 161887 164023 161921 164051
rect 161949 164023 171717 164051
rect 171745 164023 171779 164051
rect 171807 164023 171841 164051
rect 171869 164023 171903 164051
rect 171931 164023 177219 164051
rect 177247 164023 177281 164051
rect 177309 164023 187077 164051
rect 187105 164023 187139 164051
rect 187167 164023 187201 164051
rect 187229 164023 187263 164051
rect 187291 164023 192579 164051
rect 192607 164023 192641 164051
rect 192669 164023 202437 164051
rect 202465 164023 202499 164051
rect 202527 164023 202561 164051
rect 202589 164023 202623 164051
rect 202651 164023 207939 164051
rect 207967 164023 208001 164051
rect 208029 164023 217797 164051
rect 217825 164023 217859 164051
rect 217887 164023 217921 164051
rect 217949 164023 217983 164051
rect 218011 164023 223299 164051
rect 223327 164023 223361 164051
rect 223389 164023 233157 164051
rect 233185 164023 233219 164051
rect 233247 164023 233281 164051
rect 233309 164023 233343 164051
rect 233371 164023 238659 164051
rect 238687 164023 238721 164051
rect 238749 164023 248517 164051
rect 248545 164023 248579 164051
rect 248607 164023 248641 164051
rect 248669 164023 248703 164051
rect 248731 164023 254019 164051
rect 254047 164023 254081 164051
rect 254109 164023 263877 164051
rect 263905 164023 263939 164051
rect 263967 164023 264001 164051
rect 264029 164023 264063 164051
rect 264091 164023 269379 164051
rect 269407 164023 269441 164051
rect 269469 164023 279237 164051
rect 279265 164023 279299 164051
rect 279327 164023 279361 164051
rect 279389 164023 279423 164051
rect 279451 164023 284739 164051
rect 284767 164023 284801 164051
rect 284829 164023 294597 164051
rect 294625 164023 294659 164051
rect 294687 164023 294721 164051
rect 294749 164023 294783 164051
rect 294811 164023 298248 164051
rect 298276 164023 298310 164051
rect 298338 164023 298372 164051
rect 298400 164023 298434 164051
rect 298462 164023 298990 164051
rect -958 163989 298990 164023
rect -958 163961 -430 163989
rect -402 163961 -368 163989
rect -340 163961 -306 163989
rect -278 163961 -244 163989
rect -216 163961 2757 163989
rect 2785 163961 2819 163989
rect 2847 163961 2881 163989
rect 2909 163961 2943 163989
rect 2971 163961 8259 163989
rect 8287 163961 8321 163989
rect 8349 163961 18117 163989
rect 18145 163961 18179 163989
rect 18207 163961 18241 163989
rect 18269 163961 18303 163989
rect 18331 163961 23619 163989
rect 23647 163961 23681 163989
rect 23709 163961 33477 163989
rect 33505 163961 33539 163989
rect 33567 163961 33601 163989
rect 33629 163961 33663 163989
rect 33691 163961 38979 163989
rect 39007 163961 39041 163989
rect 39069 163961 48837 163989
rect 48865 163961 48899 163989
rect 48927 163961 48961 163989
rect 48989 163961 49023 163989
rect 49051 163961 54339 163989
rect 54367 163961 54401 163989
rect 54429 163961 64197 163989
rect 64225 163961 64259 163989
rect 64287 163961 64321 163989
rect 64349 163961 64383 163989
rect 64411 163961 69699 163989
rect 69727 163961 69761 163989
rect 69789 163961 79557 163989
rect 79585 163961 79619 163989
rect 79647 163961 79681 163989
rect 79709 163961 79743 163989
rect 79771 163961 85059 163989
rect 85087 163961 85121 163989
rect 85149 163961 94917 163989
rect 94945 163961 94979 163989
rect 95007 163961 95041 163989
rect 95069 163961 95103 163989
rect 95131 163961 100419 163989
rect 100447 163961 100481 163989
rect 100509 163961 110277 163989
rect 110305 163961 110339 163989
rect 110367 163961 110401 163989
rect 110429 163961 110463 163989
rect 110491 163961 115779 163989
rect 115807 163961 115841 163989
rect 115869 163961 125637 163989
rect 125665 163961 125699 163989
rect 125727 163961 125761 163989
rect 125789 163961 125823 163989
rect 125851 163961 131139 163989
rect 131167 163961 131201 163989
rect 131229 163961 140997 163989
rect 141025 163961 141059 163989
rect 141087 163961 141121 163989
rect 141149 163961 141183 163989
rect 141211 163961 146499 163989
rect 146527 163961 146561 163989
rect 146589 163961 156357 163989
rect 156385 163961 156419 163989
rect 156447 163961 156481 163989
rect 156509 163961 156543 163989
rect 156571 163961 161859 163989
rect 161887 163961 161921 163989
rect 161949 163961 171717 163989
rect 171745 163961 171779 163989
rect 171807 163961 171841 163989
rect 171869 163961 171903 163989
rect 171931 163961 177219 163989
rect 177247 163961 177281 163989
rect 177309 163961 187077 163989
rect 187105 163961 187139 163989
rect 187167 163961 187201 163989
rect 187229 163961 187263 163989
rect 187291 163961 192579 163989
rect 192607 163961 192641 163989
rect 192669 163961 202437 163989
rect 202465 163961 202499 163989
rect 202527 163961 202561 163989
rect 202589 163961 202623 163989
rect 202651 163961 207939 163989
rect 207967 163961 208001 163989
rect 208029 163961 217797 163989
rect 217825 163961 217859 163989
rect 217887 163961 217921 163989
rect 217949 163961 217983 163989
rect 218011 163961 223299 163989
rect 223327 163961 223361 163989
rect 223389 163961 233157 163989
rect 233185 163961 233219 163989
rect 233247 163961 233281 163989
rect 233309 163961 233343 163989
rect 233371 163961 238659 163989
rect 238687 163961 238721 163989
rect 238749 163961 248517 163989
rect 248545 163961 248579 163989
rect 248607 163961 248641 163989
rect 248669 163961 248703 163989
rect 248731 163961 254019 163989
rect 254047 163961 254081 163989
rect 254109 163961 263877 163989
rect 263905 163961 263939 163989
rect 263967 163961 264001 163989
rect 264029 163961 264063 163989
rect 264091 163961 269379 163989
rect 269407 163961 269441 163989
rect 269469 163961 279237 163989
rect 279265 163961 279299 163989
rect 279327 163961 279361 163989
rect 279389 163961 279423 163989
rect 279451 163961 284739 163989
rect 284767 163961 284801 163989
rect 284829 163961 294597 163989
rect 294625 163961 294659 163989
rect 294687 163961 294721 163989
rect 294749 163961 294783 163989
rect 294811 163961 298248 163989
rect 298276 163961 298310 163989
rect 298338 163961 298372 163989
rect 298400 163961 298434 163989
rect 298462 163961 298990 163989
rect -958 163913 298990 163961
rect -958 158175 298990 158223
rect -958 158147 -910 158175
rect -882 158147 -848 158175
rect -820 158147 -786 158175
rect -758 158147 -724 158175
rect -696 158147 4617 158175
rect 4645 158147 4679 158175
rect 4707 158147 4741 158175
rect 4769 158147 4803 158175
rect 4831 158147 15939 158175
rect 15967 158147 16001 158175
rect 16029 158147 19977 158175
rect 20005 158147 20039 158175
rect 20067 158147 20101 158175
rect 20129 158147 20163 158175
rect 20191 158147 31299 158175
rect 31327 158147 31361 158175
rect 31389 158147 35337 158175
rect 35365 158147 35399 158175
rect 35427 158147 35461 158175
rect 35489 158147 35523 158175
rect 35551 158147 46659 158175
rect 46687 158147 46721 158175
rect 46749 158147 50697 158175
rect 50725 158147 50759 158175
rect 50787 158147 50821 158175
rect 50849 158147 50883 158175
rect 50911 158147 62019 158175
rect 62047 158147 62081 158175
rect 62109 158147 66057 158175
rect 66085 158147 66119 158175
rect 66147 158147 66181 158175
rect 66209 158147 66243 158175
rect 66271 158147 77379 158175
rect 77407 158147 77441 158175
rect 77469 158147 81417 158175
rect 81445 158147 81479 158175
rect 81507 158147 81541 158175
rect 81569 158147 81603 158175
rect 81631 158147 92739 158175
rect 92767 158147 92801 158175
rect 92829 158147 96777 158175
rect 96805 158147 96839 158175
rect 96867 158147 96901 158175
rect 96929 158147 96963 158175
rect 96991 158147 108099 158175
rect 108127 158147 108161 158175
rect 108189 158147 112137 158175
rect 112165 158147 112199 158175
rect 112227 158147 112261 158175
rect 112289 158147 112323 158175
rect 112351 158147 123459 158175
rect 123487 158147 123521 158175
rect 123549 158147 127497 158175
rect 127525 158147 127559 158175
rect 127587 158147 127621 158175
rect 127649 158147 127683 158175
rect 127711 158147 138819 158175
rect 138847 158147 138881 158175
rect 138909 158147 142857 158175
rect 142885 158147 142919 158175
rect 142947 158147 142981 158175
rect 143009 158147 143043 158175
rect 143071 158147 154179 158175
rect 154207 158147 154241 158175
rect 154269 158147 158217 158175
rect 158245 158147 158279 158175
rect 158307 158147 158341 158175
rect 158369 158147 158403 158175
rect 158431 158147 169539 158175
rect 169567 158147 169601 158175
rect 169629 158147 173577 158175
rect 173605 158147 173639 158175
rect 173667 158147 173701 158175
rect 173729 158147 173763 158175
rect 173791 158147 184899 158175
rect 184927 158147 184961 158175
rect 184989 158147 188937 158175
rect 188965 158147 188999 158175
rect 189027 158147 189061 158175
rect 189089 158147 189123 158175
rect 189151 158147 200259 158175
rect 200287 158147 200321 158175
rect 200349 158147 204297 158175
rect 204325 158147 204359 158175
rect 204387 158147 204421 158175
rect 204449 158147 204483 158175
rect 204511 158147 215619 158175
rect 215647 158147 215681 158175
rect 215709 158147 219657 158175
rect 219685 158147 219719 158175
rect 219747 158147 219781 158175
rect 219809 158147 219843 158175
rect 219871 158147 230979 158175
rect 231007 158147 231041 158175
rect 231069 158147 235017 158175
rect 235045 158147 235079 158175
rect 235107 158147 235141 158175
rect 235169 158147 235203 158175
rect 235231 158147 246339 158175
rect 246367 158147 246401 158175
rect 246429 158147 250377 158175
rect 250405 158147 250439 158175
rect 250467 158147 250501 158175
rect 250529 158147 250563 158175
rect 250591 158147 261699 158175
rect 261727 158147 261761 158175
rect 261789 158147 265737 158175
rect 265765 158147 265799 158175
rect 265827 158147 265861 158175
rect 265889 158147 265923 158175
rect 265951 158147 277059 158175
rect 277087 158147 277121 158175
rect 277149 158147 281097 158175
rect 281125 158147 281159 158175
rect 281187 158147 281221 158175
rect 281249 158147 281283 158175
rect 281311 158147 296457 158175
rect 296485 158147 296519 158175
rect 296547 158147 296581 158175
rect 296609 158147 296643 158175
rect 296671 158147 298728 158175
rect 298756 158147 298790 158175
rect 298818 158147 298852 158175
rect 298880 158147 298914 158175
rect 298942 158147 298990 158175
rect -958 158113 298990 158147
rect -958 158085 -910 158113
rect -882 158085 -848 158113
rect -820 158085 -786 158113
rect -758 158085 -724 158113
rect -696 158085 4617 158113
rect 4645 158085 4679 158113
rect 4707 158085 4741 158113
rect 4769 158085 4803 158113
rect 4831 158085 15939 158113
rect 15967 158085 16001 158113
rect 16029 158085 19977 158113
rect 20005 158085 20039 158113
rect 20067 158085 20101 158113
rect 20129 158085 20163 158113
rect 20191 158085 31299 158113
rect 31327 158085 31361 158113
rect 31389 158085 35337 158113
rect 35365 158085 35399 158113
rect 35427 158085 35461 158113
rect 35489 158085 35523 158113
rect 35551 158085 46659 158113
rect 46687 158085 46721 158113
rect 46749 158085 50697 158113
rect 50725 158085 50759 158113
rect 50787 158085 50821 158113
rect 50849 158085 50883 158113
rect 50911 158085 62019 158113
rect 62047 158085 62081 158113
rect 62109 158085 66057 158113
rect 66085 158085 66119 158113
rect 66147 158085 66181 158113
rect 66209 158085 66243 158113
rect 66271 158085 77379 158113
rect 77407 158085 77441 158113
rect 77469 158085 81417 158113
rect 81445 158085 81479 158113
rect 81507 158085 81541 158113
rect 81569 158085 81603 158113
rect 81631 158085 92739 158113
rect 92767 158085 92801 158113
rect 92829 158085 96777 158113
rect 96805 158085 96839 158113
rect 96867 158085 96901 158113
rect 96929 158085 96963 158113
rect 96991 158085 108099 158113
rect 108127 158085 108161 158113
rect 108189 158085 112137 158113
rect 112165 158085 112199 158113
rect 112227 158085 112261 158113
rect 112289 158085 112323 158113
rect 112351 158085 123459 158113
rect 123487 158085 123521 158113
rect 123549 158085 127497 158113
rect 127525 158085 127559 158113
rect 127587 158085 127621 158113
rect 127649 158085 127683 158113
rect 127711 158085 138819 158113
rect 138847 158085 138881 158113
rect 138909 158085 142857 158113
rect 142885 158085 142919 158113
rect 142947 158085 142981 158113
rect 143009 158085 143043 158113
rect 143071 158085 154179 158113
rect 154207 158085 154241 158113
rect 154269 158085 158217 158113
rect 158245 158085 158279 158113
rect 158307 158085 158341 158113
rect 158369 158085 158403 158113
rect 158431 158085 169539 158113
rect 169567 158085 169601 158113
rect 169629 158085 173577 158113
rect 173605 158085 173639 158113
rect 173667 158085 173701 158113
rect 173729 158085 173763 158113
rect 173791 158085 184899 158113
rect 184927 158085 184961 158113
rect 184989 158085 188937 158113
rect 188965 158085 188999 158113
rect 189027 158085 189061 158113
rect 189089 158085 189123 158113
rect 189151 158085 200259 158113
rect 200287 158085 200321 158113
rect 200349 158085 204297 158113
rect 204325 158085 204359 158113
rect 204387 158085 204421 158113
rect 204449 158085 204483 158113
rect 204511 158085 215619 158113
rect 215647 158085 215681 158113
rect 215709 158085 219657 158113
rect 219685 158085 219719 158113
rect 219747 158085 219781 158113
rect 219809 158085 219843 158113
rect 219871 158085 230979 158113
rect 231007 158085 231041 158113
rect 231069 158085 235017 158113
rect 235045 158085 235079 158113
rect 235107 158085 235141 158113
rect 235169 158085 235203 158113
rect 235231 158085 246339 158113
rect 246367 158085 246401 158113
rect 246429 158085 250377 158113
rect 250405 158085 250439 158113
rect 250467 158085 250501 158113
rect 250529 158085 250563 158113
rect 250591 158085 261699 158113
rect 261727 158085 261761 158113
rect 261789 158085 265737 158113
rect 265765 158085 265799 158113
rect 265827 158085 265861 158113
rect 265889 158085 265923 158113
rect 265951 158085 277059 158113
rect 277087 158085 277121 158113
rect 277149 158085 281097 158113
rect 281125 158085 281159 158113
rect 281187 158085 281221 158113
rect 281249 158085 281283 158113
rect 281311 158085 296457 158113
rect 296485 158085 296519 158113
rect 296547 158085 296581 158113
rect 296609 158085 296643 158113
rect 296671 158085 298728 158113
rect 298756 158085 298790 158113
rect 298818 158085 298852 158113
rect 298880 158085 298914 158113
rect 298942 158085 298990 158113
rect -958 158051 298990 158085
rect -958 158023 -910 158051
rect -882 158023 -848 158051
rect -820 158023 -786 158051
rect -758 158023 -724 158051
rect -696 158023 4617 158051
rect 4645 158023 4679 158051
rect 4707 158023 4741 158051
rect 4769 158023 4803 158051
rect 4831 158023 15939 158051
rect 15967 158023 16001 158051
rect 16029 158023 19977 158051
rect 20005 158023 20039 158051
rect 20067 158023 20101 158051
rect 20129 158023 20163 158051
rect 20191 158023 31299 158051
rect 31327 158023 31361 158051
rect 31389 158023 35337 158051
rect 35365 158023 35399 158051
rect 35427 158023 35461 158051
rect 35489 158023 35523 158051
rect 35551 158023 46659 158051
rect 46687 158023 46721 158051
rect 46749 158023 50697 158051
rect 50725 158023 50759 158051
rect 50787 158023 50821 158051
rect 50849 158023 50883 158051
rect 50911 158023 62019 158051
rect 62047 158023 62081 158051
rect 62109 158023 66057 158051
rect 66085 158023 66119 158051
rect 66147 158023 66181 158051
rect 66209 158023 66243 158051
rect 66271 158023 77379 158051
rect 77407 158023 77441 158051
rect 77469 158023 81417 158051
rect 81445 158023 81479 158051
rect 81507 158023 81541 158051
rect 81569 158023 81603 158051
rect 81631 158023 92739 158051
rect 92767 158023 92801 158051
rect 92829 158023 96777 158051
rect 96805 158023 96839 158051
rect 96867 158023 96901 158051
rect 96929 158023 96963 158051
rect 96991 158023 108099 158051
rect 108127 158023 108161 158051
rect 108189 158023 112137 158051
rect 112165 158023 112199 158051
rect 112227 158023 112261 158051
rect 112289 158023 112323 158051
rect 112351 158023 123459 158051
rect 123487 158023 123521 158051
rect 123549 158023 127497 158051
rect 127525 158023 127559 158051
rect 127587 158023 127621 158051
rect 127649 158023 127683 158051
rect 127711 158023 138819 158051
rect 138847 158023 138881 158051
rect 138909 158023 142857 158051
rect 142885 158023 142919 158051
rect 142947 158023 142981 158051
rect 143009 158023 143043 158051
rect 143071 158023 154179 158051
rect 154207 158023 154241 158051
rect 154269 158023 158217 158051
rect 158245 158023 158279 158051
rect 158307 158023 158341 158051
rect 158369 158023 158403 158051
rect 158431 158023 169539 158051
rect 169567 158023 169601 158051
rect 169629 158023 173577 158051
rect 173605 158023 173639 158051
rect 173667 158023 173701 158051
rect 173729 158023 173763 158051
rect 173791 158023 184899 158051
rect 184927 158023 184961 158051
rect 184989 158023 188937 158051
rect 188965 158023 188999 158051
rect 189027 158023 189061 158051
rect 189089 158023 189123 158051
rect 189151 158023 200259 158051
rect 200287 158023 200321 158051
rect 200349 158023 204297 158051
rect 204325 158023 204359 158051
rect 204387 158023 204421 158051
rect 204449 158023 204483 158051
rect 204511 158023 215619 158051
rect 215647 158023 215681 158051
rect 215709 158023 219657 158051
rect 219685 158023 219719 158051
rect 219747 158023 219781 158051
rect 219809 158023 219843 158051
rect 219871 158023 230979 158051
rect 231007 158023 231041 158051
rect 231069 158023 235017 158051
rect 235045 158023 235079 158051
rect 235107 158023 235141 158051
rect 235169 158023 235203 158051
rect 235231 158023 246339 158051
rect 246367 158023 246401 158051
rect 246429 158023 250377 158051
rect 250405 158023 250439 158051
rect 250467 158023 250501 158051
rect 250529 158023 250563 158051
rect 250591 158023 261699 158051
rect 261727 158023 261761 158051
rect 261789 158023 265737 158051
rect 265765 158023 265799 158051
rect 265827 158023 265861 158051
rect 265889 158023 265923 158051
rect 265951 158023 277059 158051
rect 277087 158023 277121 158051
rect 277149 158023 281097 158051
rect 281125 158023 281159 158051
rect 281187 158023 281221 158051
rect 281249 158023 281283 158051
rect 281311 158023 296457 158051
rect 296485 158023 296519 158051
rect 296547 158023 296581 158051
rect 296609 158023 296643 158051
rect 296671 158023 298728 158051
rect 298756 158023 298790 158051
rect 298818 158023 298852 158051
rect 298880 158023 298914 158051
rect 298942 158023 298990 158051
rect -958 157989 298990 158023
rect -958 157961 -910 157989
rect -882 157961 -848 157989
rect -820 157961 -786 157989
rect -758 157961 -724 157989
rect -696 157961 4617 157989
rect 4645 157961 4679 157989
rect 4707 157961 4741 157989
rect 4769 157961 4803 157989
rect 4831 157961 15939 157989
rect 15967 157961 16001 157989
rect 16029 157961 19977 157989
rect 20005 157961 20039 157989
rect 20067 157961 20101 157989
rect 20129 157961 20163 157989
rect 20191 157961 31299 157989
rect 31327 157961 31361 157989
rect 31389 157961 35337 157989
rect 35365 157961 35399 157989
rect 35427 157961 35461 157989
rect 35489 157961 35523 157989
rect 35551 157961 46659 157989
rect 46687 157961 46721 157989
rect 46749 157961 50697 157989
rect 50725 157961 50759 157989
rect 50787 157961 50821 157989
rect 50849 157961 50883 157989
rect 50911 157961 62019 157989
rect 62047 157961 62081 157989
rect 62109 157961 66057 157989
rect 66085 157961 66119 157989
rect 66147 157961 66181 157989
rect 66209 157961 66243 157989
rect 66271 157961 77379 157989
rect 77407 157961 77441 157989
rect 77469 157961 81417 157989
rect 81445 157961 81479 157989
rect 81507 157961 81541 157989
rect 81569 157961 81603 157989
rect 81631 157961 92739 157989
rect 92767 157961 92801 157989
rect 92829 157961 96777 157989
rect 96805 157961 96839 157989
rect 96867 157961 96901 157989
rect 96929 157961 96963 157989
rect 96991 157961 108099 157989
rect 108127 157961 108161 157989
rect 108189 157961 112137 157989
rect 112165 157961 112199 157989
rect 112227 157961 112261 157989
rect 112289 157961 112323 157989
rect 112351 157961 123459 157989
rect 123487 157961 123521 157989
rect 123549 157961 127497 157989
rect 127525 157961 127559 157989
rect 127587 157961 127621 157989
rect 127649 157961 127683 157989
rect 127711 157961 138819 157989
rect 138847 157961 138881 157989
rect 138909 157961 142857 157989
rect 142885 157961 142919 157989
rect 142947 157961 142981 157989
rect 143009 157961 143043 157989
rect 143071 157961 154179 157989
rect 154207 157961 154241 157989
rect 154269 157961 158217 157989
rect 158245 157961 158279 157989
rect 158307 157961 158341 157989
rect 158369 157961 158403 157989
rect 158431 157961 169539 157989
rect 169567 157961 169601 157989
rect 169629 157961 173577 157989
rect 173605 157961 173639 157989
rect 173667 157961 173701 157989
rect 173729 157961 173763 157989
rect 173791 157961 184899 157989
rect 184927 157961 184961 157989
rect 184989 157961 188937 157989
rect 188965 157961 188999 157989
rect 189027 157961 189061 157989
rect 189089 157961 189123 157989
rect 189151 157961 200259 157989
rect 200287 157961 200321 157989
rect 200349 157961 204297 157989
rect 204325 157961 204359 157989
rect 204387 157961 204421 157989
rect 204449 157961 204483 157989
rect 204511 157961 215619 157989
rect 215647 157961 215681 157989
rect 215709 157961 219657 157989
rect 219685 157961 219719 157989
rect 219747 157961 219781 157989
rect 219809 157961 219843 157989
rect 219871 157961 230979 157989
rect 231007 157961 231041 157989
rect 231069 157961 235017 157989
rect 235045 157961 235079 157989
rect 235107 157961 235141 157989
rect 235169 157961 235203 157989
rect 235231 157961 246339 157989
rect 246367 157961 246401 157989
rect 246429 157961 250377 157989
rect 250405 157961 250439 157989
rect 250467 157961 250501 157989
rect 250529 157961 250563 157989
rect 250591 157961 261699 157989
rect 261727 157961 261761 157989
rect 261789 157961 265737 157989
rect 265765 157961 265799 157989
rect 265827 157961 265861 157989
rect 265889 157961 265923 157989
rect 265951 157961 277059 157989
rect 277087 157961 277121 157989
rect 277149 157961 281097 157989
rect 281125 157961 281159 157989
rect 281187 157961 281221 157989
rect 281249 157961 281283 157989
rect 281311 157961 296457 157989
rect 296485 157961 296519 157989
rect 296547 157961 296581 157989
rect 296609 157961 296643 157989
rect 296671 157961 298728 157989
rect 298756 157961 298790 157989
rect 298818 157961 298852 157989
rect 298880 157961 298914 157989
rect 298942 157961 298990 157989
rect -958 157913 298990 157961
rect -958 155175 298990 155223
rect -958 155147 -430 155175
rect -402 155147 -368 155175
rect -340 155147 -306 155175
rect -278 155147 -244 155175
rect -216 155147 2757 155175
rect 2785 155147 2819 155175
rect 2847 155147 2881 155175
rect 2909 155147 2943 155175
rect 2971 155147 8259 155175
rect 8287 155147 8321 155175
rect 8349 155147 18117 155175
rect 18145 155147 18179 155175
rect 18207 155147 18241 155175
rect 18269 155147 18303 155175
rect 18331 155147 23619 155175
rect 23647 155147 23681 155175
rect 23709 155147 33477 155175
rect 33505 155147 33539 155175
rect 33567 155147 33601 155175
rect 33629 155147 33663 155175
rect 33691 155147 38979 155175
rect 39007 155147 39041 155175
rect 39069 155147 48837 155175
rect 48865 155147 48899 155175
rect 48927 155147 48961 155175
rect 48989 155147 49023 155175
rect 49051 155147 54339 155175
rect 54367 155147 54401 155175
rect 54429 155147 64197 155175
rect 64225 155147 64259 155175
rect 64287 155147 64321 155175
rect 64349 155147 64383 155175
rect 64411 155147 69699 155175
rect 69727 155147 69761 155175
rect 69789 155147 79557 155175
rect 79585 155147 79619 155175
rect 79647 155147 79681 155175
rect 79709 155147 79743 155175
rect 79771 155147 85059 155175
rect 85087 155147 85121 155175
rect 85149 155147 94917 155175
rect 94945 155147 94979 155175
rect 95007 155147 95041 155175
rect 95069 155147 95103 155175
rect 95131 155147 100419 155175
rect 100447 155147 100481 155175
rect 100509 155147 110277 155175
rect 110305 155147 110339 155175
rect 110367 155147 110401 155175
rect 110429 155147 110463 155175
rect 110491 155147 115779 155175
rect 115807 155147 115841 155175
rect 115869 155147 125637 155175
rect 125665 155147 125699 155175
rect 125727 155147 125761 155175
rect 125789 155147 125823 155175
rect 125851 155147 131139 155175
rect 131167 155147 131201 155175
rect 131229 155147 140997 155175
rect 141025 155147 141059 155175
rect 141087 155147 141121 155175
rect 141149 155147 141183 155175
rect 141211 155147 146499 155175
rect 146527 155147 146561 155175
rect 146589 155147 156357 155175
rect 156385 155147 156419 155175
rect 156447 155147 156481 155175
rect 156509 155147 156543 155175
rect 156571 155147 161859 155175
rect 161887 155147 161921 155175
rect 161949 155147 171717 155175
rect 171745 155147 171779 155175
rect 171807 155147 171841 155175
rect 171869 155147 171903 155175
rect 171931 155147 177219 155175
rect 177247 155147 177281 155175
rect 177309 155147 187077 155175
rect 187105 155147 187139 155175
rect 187167 155147 187201 155175
rect 187229 155147 187263 155175
rect 187291 155147 192579 155175
rect 192607 155147 192641 155175
rect 192669 155147 202437 155175
rect 202465 155147 202499 155175
rect 202527 155147 202561 155175
rect 202589 155147 202623 155175
rect 202651 155147 207939 155175
rect 207967 155147 208001 155175
rect 208029 155147 217797 155175
rect 217825 155147 217859 155175
rect 217887 155147 217921 155175
rect 217949 155147 217983 155175
rect 218011 155147 223299 155175
rect 223327 155147 223361 155175
rect 223389 155147 233157 155175
rect 233185 155147 233219 155175
rect 233247 155147 233281 155175
rect 233309 155147 233343 155175
rect 233371 155147 238659 155175
rect 238687 155147 238721 155175
rect 238749 155147 248517 155175
rect 248545 155147 248579 155175
rect 248607 155147 248641 155175
rect 248669 155147 248703 155175
rect 248731 155147 254019 155175
rect 254047 155147 254081 155175
rect 254109 155147 263877 155175
rect 263905 155147 263939 155175
rect 263967 155147 264001 155175
rect 264029 155147 264063 155175
rect 264091 155147 269379 155175
rect 269407 155147 269441 155175
rect 269469 155147 279237 155175
rect 279265 155147 279299 155175
rect 279327 155147 279361 155175
rect 279389 155147 279423 155175
rect 279451 155147 284739 155175
rect 284767 155147 284801 155175
rect 284829 155147 294597 155175
rect 294625 155147 294659 155175
rect 294687 155147 294721 155175
rect 294749 155147 294783 155175
rect 294811 155147 298248 155175
rect 298276 155147 298310 155175
rect 298338 155147 298372 155175
rect 298400 155147 298434 155175
rect 298462 155147 298990 155175
rect -958 155113 298990 155147
rect -958 155085 -430 155113
rect -402 155085 -368 155113
rect -340 155085 -306 155113
rect -278 155085 -244 155113
rect -216 155085 2757 155113
rect 2785 155085 2819 155113
rect 2847 155085 2881 155113
rect 2909 155085 2943 155113
rect 2971 155085 8259 155113
rect 8287 155085 8321 155113
rect 8349 155085 18117 155113
rect 18145 155085 18179 155113
rect 18207 155085 18241 155113
rect 18269 155085 18303 155113
rect 18331 155085 23619 155113
rect 23647 155085 23681 155113
rect 23709 155085 33477 155113
rect 33505 155085 33539 155113
rect 33567 155085 33601 155113
rect 33629 155085 33663 155113
rect 33691 155085 38979 155113
rect 39007 155085 39041 155113
rect 39069 155085 48837 155113
rect 48865 155085 48899 155113
rect 48927 155085 48961 155113
rect 48989 155085 49023 155113
rect 49051 155085 54339 155113
rect 54367 155085 54401 155113
rect 54429 155085 64197 155113
rect 64225 155085 64259 155113
rect 64287 155085 64321 155113
rect 64349 155085 64383 155113
rect 64411 155085 69699 155113
rect 69727 155085 69761 155113
rect 69789 155085 79557 155113
rect 79585 155085 79619 155113
rect 79647 155085 79681 155113
rect 79709 155085 79743 155113
rect 79771 155085 85059 155113
rect 85087 155085 85121 155113
rect 85149 155085 94917 155113
rect 94945 155085 94979 155113
rect 95007 155085 95041 155113
rect 95069 155085 95103 155113
rect 95131 155085 100419 155113
rect 100447 155085 100481 155113
rect 100509 155085 110277 155113
rect 110305 155085 110339 155113
rect 110367 155085 110401 155113
rect 110429 155085 110463 155113
rect 110491 155085 115779 155113
rect 115807 155085 115841 155113
rect 115869 155085 125637 155113
rect 125665 155085 125699 155113
rect 125727 155085 125761 155113
rect 125789 155085 125823 155113
rect 125851 155085 131139 155113
rect 131167 155085 131201 155113
rect 131229 155085 140997 155113
rect 141025 155085 141059 155113
rect 141087 155085 141121 155113
rect 141149 155085 141183 155113
rect 141211 155085 146499 155113
rect 146527 155085 146561 155113
rect 146589 155085 156357 155113
rect 156385 155085 156419 155113
rect 156447 155085 156481 155113
rect 156509 155085 156543 155113
rect 156571 155085 161859 155113
rect 161887 155085 161921 155113
rect 161949 155085 171717 155113
rect 171745 155085 171779 155113
rect 171807 155085 171841 155113
rect 171869 155085 171903 155113
rect 171931 155085 177219 155113
rect 177247 155085 177281 155113
rect 177309 155085 187077 155113
rect 187105 155085 187139 155113
rect 187167 155085 187201 155113
rect 187229 155085 187263 155113
rect 187291 155085 192579 155113
rect 192607 155085 192641 155113
rect 192669 155085 202437 155113
rect 202465 155085 202499 155113
rect 202527 155085 202561 155113
rect 202589 155085 202623 155113
rect 202651 155085 207939 155113
rect 207967 155085 208001 155113
rect 208029 155085 217797 155113
rect 217825 155085 217859 155113
rect 217887 155085 217921 155113
rect 217949 155085 217983 155113
rect 218011 155085 223299 155113
rect 223327 155085 223361 155113
rect 223389 155085 233157 155113
rect 233185 155085 233219 155113
rect 233247 155085 233281 155113
rect 233309 155085 233343 155113
rect 233371 155085 238659 155113
rect 238687 155085 238721 155113
rect 238749 155085 248517 155113
rect 248545 155085 248579 155113
rect 248607 155085 248641 155113
rect 248669 155085 248703 155113
rect 248731 155085 254019 155113
rect 254047 155085 254081 155113
rect 254109 155085 263877 155113
rect 263905 155085 263939 155113
rect 263967 155085 264001 155113
rect 264029 155085 264063 155113
rect 264091 155085 269379 155113
rect 269407 155085 269441 155113
rect 269469 155085 279237 155113
rect 279265 155085 279299 155113
rect 279327 155085 279361 155113
rect 279389 155085 279423 155113
rect 279451 155085 284739 155113
rect 284767 155085 284801 155113
rect 284829 155085 294597 155113
rect 294625 155085 294659 155113
rect 294687 155085 294721 155113
rect 294749 155085 294783 155113
rect 294811 155085 298248 155113
rect 298276 155085 298310 155113
rect 298338 155085 298372 155113
rect 298400 155085 298434 155113
rect 298462 155085 298990 155113
rect -958 155051 298990 155085
rect -958 155023 -430 155051
rect -402 155023 -368 155051
rect -340 155023 -306 155051
rect -278 155023 -244 155051
rect -216 155023 2757 155051
rect 2785 155023 2819 155051
rect 2847 155023 2881 155051
rect 2909 155023 2943 155051
rect 2971 155023 8259 155051
rect 8287 155023 8321 155051
rect 8349 155023 18117 155051
rect 18145 155023 18179 155051
rect 18207 155023 18241 155051
rect 18269 155023 18303 155051
rect 18331 155023 23619 155051
rect 23647 155023 23681 155051
rect 23709 155023 33477 155051
rect 33505 155023 33539 155051
rect 33567 155023 33601 155051
rect 33629 155023 33663 155051
rect 33691 155023 38979 155051
rect 39007 155023 39041 155051
rect 39069 155023 48837 155051
rect 48865 155023 48899 155051
rect 48927 155023 48961 155051
rect 48989 155023 49023 155051
rect 49051 155023 54339 155051
rect 54367 155023 54401 155051
rect 54429 155023 64197 155051
rect 64225 155023 64259 155051
rect 64287 155023 64321 155051
rect 64349 155023 64383 155051
rect 64411 155023 69699 155051
rect 69727 155023 69761 155051
rect 69789 155023 79557 155051
rect 79585 155023 79619 155051
rect 79647 155023 79681 155051
rect 79709 155023 79743 155051
rect 79771 155023 85059 155051
rect 85087 155023 85121 155051
rect 85149 155023 94917 155051
rect 94945 155023 94979 155051
rect 95007 155023 95041 155051
rect 95069 155023 95103 155051
rect 95131 155023 100419 155051
rect 100447 155023 100481 155051
rect 100509 155023 110277 155051
rect 110305 155023 110339 155051
rect 110367 155023 110401 155051
rect 110429 155023 110463 155051
rect 110491 155023 115779 155051
rect 115807 155023 115841 155051
rect 115869 155023 125637 155051
rect 125665 155023 125699 155051
rect 125727 155023 125761 155051
rect 125789 155023 125823 155051
rect 125851 155023 131139 155051
rect 131167 155023 131201 155051
rect 131229 155023 140997 155051
rect 141025 155023 141059 155051
rect 141087 155023 141121 155051
rect 141149 155023 141183 155051
rect 141211 155023 146499 155051
rect 146527 155023 146561 155051
rect 146589 155023 156357 155051
rect 156385 155023 156419 155051
rect 156447 155023 156481 155051
rect 156509 155023 156543 155051
rect 156571 155023 161859 155051
rect 161887 155023 161921 155051
rect 161949 155023 171717 155051
rect 171745 155023 171779 155051
rect 171807 155023 171841 155051
rect 171869 155023 171903 155051
rect 171931 155023 177219 155051
rect 177247 155023 177281 155051
rect 177309 155023 187077 155051
rect 187105 155023 187139 155051
rect 187167 155023 187201 155051
rect 187229 155023 187263 155051
rect 187291 155023 192579 155051
rect 192607 155023 192641 155051
rect 192669 155023 202437 155051
rect 202465 155023 202499 155051
rect 202527 155023 202561 155051
rect 202589 155023 202623 155051
rect 202651 155023 207939 155051
rect 207967 155023 208001 155051
rect 208029 155023 217797 155051
rect 217825 155023 217859 155051
rect 217887 155023 217921 155051
rect 217949 155023 217983 155051
rect 218011 155023 223299 155051
rect 223327 155023 223361 155051
rect 223389 155023 233157 155051
rect 233185 155023 233219 155051
rect 233247 155023 233281 155051
rect 233309 155023 233343 155051
rect 233371 155023 238659 155051
rect 238687 155023 238721 155051
rect 238749 155023 248517 155051
rect 248545 155023 248579 155051
rect 248607 155023 248641 155051
rect 248669 155023 248703 155051
rect 248731 155023 254019 155051
rect 254047 155023 254081 155051
rect 254109 155023 263877 155051
rect 263905 155023 263939 155051
rect 263967 155023 264001 155051
rect 264029 155023 264063 155051
rect 264091 155023 269379 155051
rect 269407 155023 269441 155051
rect 269469 155023 279237 155051
rect 279265 155023 279299 155051
rect 279327 155023 279361 155051
rect 279389 155023 279423 155051
rect 279451 155023 284739 155051
rect 284767 155023 284801 155051
rect 284829 155023 294597 155051
rect 294625 155023 294659 155051
rect 294687 155023 294721 155051
rect 294749 155023 294783 155051
rect 294811 155023 298248 155051
rect 298276 155023 298310 155051
rect 298338 155023 298372 155051
rect 298400 155023 298434 155051
rect 298462 155023 298990 155051
rect -958 154989 298990 155023
rect -958 154961 -430 154989
rect -402 154961 -368 154989
rect -340 154961 -306 154989
rect -278 154961 -244 154989
rect -216 154961 2757 154989
rect 2785 154961 2819 154989
rect 2847 154961 2881 154989
rect 2909 154961 2943 154989
rect 2971 154961 8259 154989
rect 8287 154961 8321 154989
rect 8349 154961 18117 154989
rect 18145 154961 18179 154989
rect 18207 154961 18241 154989
rect 18269 154961 18303 154989
rect 18331 154961 23619 154989
rect 23647 154961 23681 154989
rect 23709 154961 33477 154989
rect 33505 154961 33539 154989
rect 33567 154961 33601 154989
rect 33629 154961 33663 154989
rect 33691 154961 38979 154989
rect 39007 154961 39041 154989
rect 39069 154961 48837 154989
rect 48865 154961 48899 154989
rect 48927 154961 48961 154989
rect 48989 154961 49023 154989
rect 49051 154961 54339 154989
rect 54367 154961 54401 154989
rect 54429 154961 64197 154989
rect 64225 154961 64259 154989
rect 64287 154961 64321 154989
rect 64349 154961 64383 154989
rect 64411 154961 69699 154989
rect 69727 154961 69761 154989
rect 69789 154961 79557 154989
rect 79585 154961 79619 154989
rect 79647 154961 79681 154989
rect 79709 154961 79743 154989
rect 79771 154961 85059 154989
rect 85087 154961 85121 154989
rect 85149 154961 94917 154989
rect 94945 154961 94979 154989
rect 95007 154961 95041 154989
rect 95069 154961 95103 154989
rect 95131 154961 100419 154989
rect 100447 154961 100481 154989
rect 100509 154961 110277 154989
rect 110305 154961 110339 154989
rect 110367 154961 110401 154989
rect 110429 154961 110463 154989
rect 110491 154961 115779 154989
rect 115807 154961 115841 154989
rect 115869 154961 125637 154989
rect 125665 154961 125699 154989
rect 125727 154961 125761 154989
rect 125789 154961 125823 154989
rect 125851 154961 131139 154989
rect 131167 154961 131201 154989
rect 131229 154961 140997 154989
rect 141025 154961 141059 154989
rect 141087 154961 141121 154989
rect 141149 154961 141183 154989
rect 141211 154961 146499 154989
rect 146527 154961 146561 154989
rect 146589 154961 156357 154989
rect 156385 154961 156419 154989
rect 156447 154961 156481 154989
rect 156509 154961 156543 154989
rect 156571 154961 161859 154989
rect 161887 154961 161921 154989
rect 161949 154961 171717 154989
rect 171745 154961 171779 154989
rect 171807 154961 171841 154989
rect 171869 154961 171903 154989
rect 171931 154961 177219 154989
rect 177247 154961 177281 154989
rect 177309 154961 187077 154989
rect 187105 154961 187139 154989
rect 187167 154961 187201 154989
rect 187229 154961 187263 154989
rect 187291 154961 192579 154989
rect 192607 154961 192641 154989
rect 192669 154961 202437 154989
rect 202465 154961 202499 154989
rect 202527 154961 202561 154989
rect 202589 154961 202623 154989
rect 202651 154961 207939 154989
rect 207967 154961 208001 154989
rect 208029 154961 217797 154989
rect 217825 154961 217859 154989
rect 217887 154961 217921 154989
rect 217949 154961 217983 154989
rect 218011 154961 223299 154989
rect 223327 154961 223361 154989
rect 223389 154961 233157 154989
rect 233185 154961 233219 154989
rect 233247 154961 233281 154989
rect 233309 154961 233343 154989
rect 233371 154961 238659 154989
rect 238687 154961 238721 154989
rect 238749 154961 248517 154989
rect 248545 154961 248579 154989
rect 248607 154961 248641 154989
rect 248669 154961 248703 154989
rect 248731 154961 254019 154989
rect 254047 154961 254081 154989
rect 254109 154961 263877 154989
rect 263905 154961 263939 154989
rect 263967 154961 264001 154989
rect 264029 154961 264063 154989
rect 264091 154961 269379 154989
rect 269407 154961 269441 154989
rect 269469 154961 279237 154989
rect 279265 154961 279299 154989
rect 279327 154961 279361 154989
rect 279389 154961 279423 154989
rect 279451 154961 284739 154989
rect 284767 154961 284801 154989
rect 284829 154961 294597 154989
rect 294625 154961 294659 154989
rect 294687 154961 294721 154989
rect 294749 154961 294783 154989
rect 294811 154961 298248 154989
rect 298276 154961 298310 154989
rect 298338 154961 298372 154989
rect 298400 154961 298434 154989
rect 298462 154961 298990 154989
rect -958 154913 298990 154961
rect -958 149175 298990 149223
rect -958 149147 -910 149175
rect -882 149147 -848 149175
rect -820 149147 -786 149175
rect -758 149147 -724 149175
rect -696 149147 4617 149175
rect 4645 149147 4679 149175
rect 4707 149147 4741 149175
rect 4769 149147 4803 149175
rect 4831 149147 15939 149175
rect 15967 149147 16001 149175
rect 16029 149147 19977 149175
rect 20005 149147 20039 149175
rect 20067 149147 20101 149175
rect 20129 149147 20163 149175
rect 20191 149147 31299 149175
rect 31327 149147 31361 149175
rect 31389 149147 35337 149175
rect 35365 149147 35399 149175
rect 35427 149147 35461 149175
rect 35489 149147 35523 149175
rect 35551 149147 46659 149175
rect 46687 149147 46721 149175
rect 46749 149147 50697 149175
rect 50725 149147 50759 149175
rect 50787 149147 50821 149175
rect 50849 149147 50883 149175
rect 50911 149147 62019 149175
rect 62047 149147 62081 149175
rect 62109 149147 66057 149175
rect 66085 149147 66119 149175
rect 66147 149147 66181 149175
rect 66209 149147 66243 149175
rect 66271 149147 77379 149175
rect 77407 149147 77441 149175
rect 77469 149147 81417 149175
rect 81445 149147 81479 149175
rect 81507 149147 81541 149175
rect 81569 149147 81603 149175
rect 81631 149147 92739 149175
rect 92767 149147 92801 149175
rect 92829 149147 96777 149175
rect 96805 149147 96839 149175
rect 96867 149147 96901 149175
rect 96929 149147 96963 149175
rect 96991 149147 108099 149175
rect 108127 149147 108161 149175
rect 108189 149147 112137 149175
rect 112165 149147 112199 149175
rect 112227 149147 112261 149175
rect 112289 149147 112323 149175
rect 112351 149147 123459 149175
rect 123487 149147 123521 149175
rect 123549 149147 127497 149175
rect 127525 149147 127559 149175
rect 127587 149147 127621 149175
rect 127649 149147 127683 149175
rect 127711 149147 138819 149175
rect 138847 149147 138881 149175
rect 138909 149147 142857 149175
rect 142885 149147 142919 149175
rect 142947 149147 142981 149175
rect 143009 149147 143043 149175
rect 143071 149147 154179 149175
rect 154207 149147 154241 149175
rect 154269 149147 158217 149175
rect 158245 149147 158279 149175
rect 158307 149147 158341 149175
rect 158369 149147 158403 149175
rect 158431 149147 169539 149175
rect 169567 149147 169601 149175
rect 169629 149147 173577 149175
rect 173605 149147 173639 149175
rect 173667 149147 173701 149175
rect 173729 149147 173763 149175
rect 173791 149147 184899 149175
rect 184927 149147 184961 149175
rect 184989 149147 188937 149175
rect 188965 149147 188999 149175
rect 189027 149147 189061 149175
rect 189089 149147 189123 149175
rect 189151 149147 200259 149175
rect 200287 149147 200321 149175
rect 200349 149147 204297 149175
rect 204325 149147 204359 149175
rect 204387 149147 204421 149175
rect 204449 149147 204483 149175
rect 204511 149147 215619 149175
rect 215647 149147 215681 149175
rect 215709 149147 219657 149175
rect 219685 149147 219719 149175
rect 219747 149147 219781 149175
rect 219809 149147 219843 149175
rect 219871 149147 230979 149175
rect 231007 149147 231041 149175
rect 231069 149147 235017 149175
rect 235045 149147 235079 149175
rect 235107 149147 235141 149175
rect 235169 149147 235203 149175
rect 235231 149147 246339 149175
rect 246367 149147 246401 149175
rect 246429 149147 250377 149175
rect 250405 149147 250439 149175
rect 250467 149147 250501 149175
rect 250529 149147 250563 149175
rect 250591 149147 261699 149175
rect 261727 149147 261761 149175
rect 261789 149147 265737 149175
rect 265765 149147 265799 149175
rect 265827 149147 265861 149175
rect 265889 149147 265923 149175
rect 265951 149147 277059 149175
rect 277087 149147 277121 149175
rect 277149 149147 281097 149175
rect 281125 149147 281159 149175
rect 281187 149147 281221 149175
rect 281249 149147 281283 149175
rect 281311 149147 296457 149175
rect 296485 149147 296519 149175
rect 296547 149147 296581 149175
rect 296609 149147 296643 149175
rect 296671 149147 298728 149175
rect 298756 149147 298790 149175
rect 298818 149147 298852 149175
rect 298880 149147 298914 149175
rect 298942 149147 298990 149175
rect -958 149113 298990 149147
rect -958 149085 -910 149113
rect -882 149085 -848 149113
rect -820 149085 -786 149113
rect -758 149085 -724 149113
rect -696 149085 4617 149113
rect 4645 149085 4679 149113
rect 4707 149085 4741 149113
rect 4769 149085 4803 149113
rect 4831 149085 15939 149113
rect 15967 149085 16001 149113
rect 16029 149085 19977 149113
rect 20005 149085 20039 149113
rect 20067 149085 20101 149113
rect 20129 149085 20163 149113
rect 20191 149085 31299 149113
rect 31327 149085 31361 149113
rect 31389 149085 35337 149113
rect 35365 149085 35399 149113
rect 35427 149085 35461 149113
rect 35489 149085 35523 149113
rect 35551 149085 46659 149113
rect 46687 149085 46721 149113
rect 46749 149085 50697 149113
rect 50725 149085 50759 149113
rect 50787 149085 50821 149113
rect 50849 149085 50883 149113
rect 50911 149085 62019 149113
rect 62047 149085 62081 149113
rect 62109 149085 66057 149113
rect 66085 149085 66119 149113
rect 66147 149085 66181 149113
rect 66209 149085 66243 149113
rect 66271 149085 77379 149113
rect 77407 149085 77441 149113
rect 77469 149085 81417 149113
rect 81445 149085 81479 149113
rect 81507 149085 81541 149113
rect 81569 149085 81603 149113
rect 81631 149085 92739 149113
rect 92767 149085 92801 149113
rect 92829 149085 96777 149113
rect 96805 149085 96839 149113
rect 96867 149085 96901 149113
rect 96929 149085 96963 149113
rect 96991 149085 108099 149113
rect 108127 149085 108161 149113
rect 108189 149085 112137 149113
rect 112165 149085 112199 149113
rect 112227 149085 112261 149113
rect 112289 149085 112323 149113
rect 112351 149085 123459 149113
rect 123487 149085 123521 149113
rect 123549 149085 127497 149113
rect 127525 149085 127559 149113
rect 127587 149085 127621 149113
rect 127649 149085 127683 149113
rect 127711 149085 138819 149113
rect 138847 149085 138881 149113
rect 138909 149085 142857 149113
rect 142885 149085 142919 149113
rect 142947 149085 142981 149113
rect 143009 149085 143043 149113
rect 143071 149085 154179 149113
rect 154207 149085 154241 149113
rect 154269 149085 158217 149113
rect 158245 149085 158279 149113
rect 158307 149085 158341 149113
rect 158369 149085 158403 149113
rect 158431 149085 169539 149113
rect 169567 149085 169601 149113
rect 169629 149085 173577 149113
rect 173605 149085 173639 149113
rect 173667 149085 173701 149113
rect 173729 149085 173763 149113
rect 173791 149085 184899 149113
rect 184927 149085 184961 149113
rect 184989 149085 188937 149113
rect 188965 149085 188999 149113
rect 189027 149085 189061 149113
rect 189089 149085 189123 149113
rect 189151 149085 200259 149113
rect 200287 149085 200321 149113
rect 200349 149085 204297 149113
rect 204325 149085 204359 149113
rect 204387 149085 204421 149113
rect 204449 149085 204483 149113
rect 204511 149085 215619 149113
rect 215647 149085 215681 149113
rect 215709 149085 219657 149113
rect 219685 149085 219719 149113
rect 219747 149085 219781 149113
rect 219809 149085 219843 149113
rect 219871 149085 230979 149113
rect 231007 149085 231041 149113
rect 231069 149085 235017 149113
rect 235045 149085 235079 149113
rect 235107 149085 235141 149113
rect 235169 149085 235203 149113
rect 235231 149085 246339 149113
rect 246367 149085 246401 149113
rect 246429 149085 250377 149113
rect 250405 149085 250439 149113
rect 250467 149085 250501 149113
rect 250529 149085 250563 149113
rect 250591 149085 261699 149113
rect 261727 149085 261761 149113
rect 261789 149085 265737 149113
rect 265765 149085 265799 149113
rect 265827 149085 265861 149113
rect 265889 149085 265923 149113
rect 265951 149085 277059 149113
rect 277087 149085 277121 149113
rect 277149 149085 281097 149113
rect 281125 149085 281159 149113
rect 281187 149085 281221 149113
rect 281249 149085 281283 149113
rect 281311 149085 296457 149113
rect 296485 149085 296519 149113
rect 296547 149085 296581 149113
rect 296609 149085 296643 149113
rect 296671 149085 298728 149113
rect 298756 149085 298790 149113
rect 298818 149085 298852 149113
rect 298880 149085 298914 149113
rect 298942 149085 298990 149113
rect -958 149051 298990 149085
rect -958 149023 -910 149051
rect -882 149023 -848 149051
rect -820 149023 -786 149051
rect -758 149023 -724 149051
rect -696 149023 4617 149051
rect 4645 149023 4679 149051
rect 4707 149023 4741 149051
rect 4769 149023 4803 149051
rect 4831 149023 15939 149051
rect 15967 149023 16001 149051
rect 16029 149023 19977 149051
rect 20005 149023 20039 149051
rect 20067 149023 20101 149051
rect 20129 149023 20163 149051
rect 20191 149023 31299 149051
rect 31327 149023 31361 149051
rect 31389 149023 35337 149051
rect 35365 149023 35399 149051
rect 35427 149023 35461 149051
rect 35489 149023 35523 149051
rect 35551 149023 46659 149051
rect 46687 149023 46721 149051
rect 46749 149023 50697 149051
rect 50725 149023 50759 149051
rect 50787 149023 50821 149051
rect 50849 149023 50883 149051
rect 50911 149023 62019 149051
rect 62047 149023 62081 149051
rect 62109 149023 66057 149051
rect 66085 149023 66119 149051
rect 66147 149023 66181 149051
rect 66209 149023 66243 149051
rect 66271 149023 77379 149051
rect 77407 149023 77441 149051
rect 77469 149023 81417 149051
rect 81445 149023 81479 149051
rect 81507 149023 81541 149051
rect 81569 149023 81603 149051
rect 81631 149023 92739 149051
rect 92767 149023 92801 149051
rect 92829 149023 96777 149051
rect 96805 149023 96839 149051
rect 96867 149023 96901 149051
rect 96929 149023 96963 149051
rect 96991 149023 108099 149051
rect 108127 149023 108161 149051
rect 108189 149023 112137 149051
rect 112165 149023 112199 149051
rect 112227 149023 112261 149051
rect 112289 149023 112323 149051
rect 112351 149023 123459 149051
rect 123487 149023 123521 149051
rect 123549 149023 127497 149051
rect 127525 149023 127559 149051
rect 127587 149023 127621 149051
rect 127649 149023 127683 149051
rect 127711 149023 138819 149051
rect 138847 149023 138881 149051
rect 138909 149023 142857 149051
rect 142885 149023 142919 149051
rect 142947 149023 142981 149051
rect 143009 149023 143043 149051
rect 143071 149023 154179 149051
rect 154207 149023 154241 149051
rect 154269 149023 158217 149051
rect 158245 149023 158279 149051
rect 158307 149023 158341 149051
rect 158369 149023 158403 149051
rect 158431 149023 169539 149051
rect 169567 149023 169601 149051
rect 169629 149023 173577 149051
rect 173605 149023 173639 149051
rect 173667 149023 173701 149051
rect 173729 149023 173763 149051
rect 173791 149023 184899 149051
rect 184927 149023 184961 149051
rect 184989 149023 188937 149051
rect 188965 149023 188999 149051
rect 189027 149023 189061 149051
rect 189089 149023 189123 149051
rect 189151 149023 200259 149051
rect 200287 149023 200321 149051
rect 200349 149023 204297 149051
rect 204325 149023 204359 149051
rect 204387 149023 204421 149051
rect 204449 149023 204483 149051
rect 204511 149023 215619 149051
rect 215647 149023 215681 149051
rect 215709 149023 219657 149051
rect 219685 149023 219719 149051
rect 219747 149023 219781 149051
rect 219809 149023 219843 149051
rect 219871 149023 230979 149051
rect 231007 149023 231041 149051
rect 231069 149023 235017 149051
rect 235045 149023 235079 149051
rect 235107 149023 235141 149051
rect 235169 149023 235203 149051
rect 235231 149023 246339 149051
rect 246367 149023 246401 149051
rect 246429 149023 250377 149051
rect 250405 149023 250439 149051
rect 250467 149023 250501 149051
rect 250529 149023 250563 149051
rect 250591 149023 261699 149051
rect 261727 149023 261761 149051
rect 261789 149023 265737 149051
rect 265765 149023 265799 149051
rect 265827 149023 265861 149051
rect 265889 149023 265923 149051
rect 265951 149023 277059 149051
rect 277087 149023 277121 149051
rect 277149 149023 281097 149051
rect 281125 149023 281159 149051
rect 281187 149023 281221 149051
rect 281249 149023 281283 149051
rect 281311 149023 296457 149051
rect 296485 149023 296519 149051
rect 296547 149023 296581 149051
rect 296609 149023 296643 149051
rect 296671 149023 298728 149051
rect 298756 149023 298790 149051
rect 298818 149023 298852 149051
rect 298880 149023 298914 149051
rect 298942 149023 298990 149051
rect -958 148989 298990 149023
rect -958 148961 -910 148989
rect -882 148961 -848 148989
rect -820 148961 -786 148989
rect -758 148961 -724 148989
rect -696 148961 4617 148989
rect 4645 148961 4679 148989
rect 4707 148961 4741 148989
rect 4769 148961 4803 148989
rect 4831 148961 15939 148989
rect 15967 148961 16001 148989
rect 16029 148961 19977 148989
rect 20005 148961 20039 148989
rect 20067 148961 20101 148989
rect 20129 148961 20163 148989
rect 20191 148961 31299 148989
rect 31327 148961 31361 148989
rect 31389 148961 35337 148989
rect 35365 148961 35399 148989
rect 35427 148961 35461 148989
rect 35489 148961 35523 148989
rect 35551 148961 46659 148989
rect 46687 148961 46721 148989
rect 46749 148961 50697 148989
rect 50725 148961 50759 148989
rect 50787 148961 50821 148989
rect 50849 148961 50883 148989
rect 50911 148961 62019 148989
rect 62047 148961 62081 148989
rect 62109 148961 66057 148989
rect 66085 148961 66119 148989
rect 66147 148961 66181 148989
rect 66209 148961 66243 148989
rect 66271 148961 77379 148989
rect 77407 148961 77441 148989
rect 77469 148961 81417 148989
rect 81445 148961 81479 148989
rect 81507 148961 81541 148989
rect 81569 148961 81603 148989
rect 81631 148961 92739 148989
rect 92767 148961 92801 148989
rect 92829 148961 96777 148989
rect 96805 148961 96839 148989
rect 96867 148961 96901 148989
rect 96929 148961 96963 148989
rect 96991 148961 108099 148989
rect 108127 148961 108161 148989
rect 108189 148961 112137 148989
rect 112165 148961 112199 148989
rect 112227 148961 112261 148989
rect 112289 148961 112323 148989
rect 112351 148961 123459 148989
rect 123487 148961 123521 148989
rect 123549 148961 127497 148989
rect 127525 148961 127559 148989
rect 127587 148961 127621 148989
rect 127649 148961 127683 148989
rect 127711 148961 138819 148989
rect 138847 148961 138881 148989
rect 138909 148961 142857 148989
rect 142885 148961 142919 148989
rect 142947 148961 142981 148989
rect 143009 148961 143043 148989
rect 143071 148961 154179 148989
rect 154207 148961 154241 148989
rect 154269 148961 158217 148989
rect 158245 148961 158279 148989
rect 158307 148961 158341 148989
rect 158369 148961 158403 148989
rect 158431 148961 169539 148989
rect 169567 148961 169601 148989
rect 169629 148961 173577 148989
rect 173605 148961 173639 148989
rect 173667 148961 173701 148989
rect 173729 148961 173763 148989
rect 173791 148961 184899 148989
rect 184927 148961 184961 148989
rect 184989 148961 188937 148989
rect 188965 148961 188999 148989
rect 189027 148961 189061 148989
rect 189089 148961 189123 148989
rect 189151 148961 200259 148989
rect 200287 148961 200321 148989
rect 200349 148961 204297 148989
rect 204325 148961 204359 148989
rect 204387 148961 204421 148989
rect 204449 148961 204483 148989
rect 204511 148961 215619 148989
rect 215647 148961 215681 148989
rect 215709 148961 219657 148989
rect 219685 148961 219719 148989
rect 219747 148961 219781 148989
rect 219809 148961 219843 148989
rect 219871 148961 230979 148989
rect 231007 148961 231041 148989
rect 231069 148961 235017 148989
rect 235045 148961 235079 148989
rect 235107 148961 235141 148989
rect 235169 148961 235203 148989
rect 235231 148961 246339 148989
rect 246367 148961 246401 148989
rect 246429 148961 250377 148989
rect 250405 148961 250439 148989
rect 250467 148961 250501 148989
rect 250529 148961 250563 148989
rect 250591 148961 261699 148989
rect 261727 148961 261761 148989
rect 261789 148961 265737 148989
rect 265765 148961 265799 148989
rect 265827 148961 265861 148989
rect 265889 148961 265923 148989
rect 265951 148961 277059 148989
rect 277087 148961 277121 148989
rect 277149 148961 281097 148989
rect 281125 148961 281159 148989
rect 281187 148961 281221 148989
rect 281249 148961 281283 148989
rect 281311 148961 296457 148989
rect 296485 148961 296519 148989
rect 296547 148961 296581 148989
rect 296609 148961 296643 148989
rect 296671 148961 298728 148989
rect 298756 148961 298790 148989
rect 298818 148961 298852 148989
rect 298880 148961 298914 148989
rect 298942 148961 298990 148989
rect -958 148913 298990 148961
rect -958 146175 298990 146223
rect -958 146147 -430 146175
rect -402 146147 -368 146175
rect -340 146147 -306 146175
rect -278 146147 -244 146175
rect -216 146147 2757 146175
rect 2785 146147 2819 146175
rect 2847 146147 2881 146175
rect 2909 146147 2943 146175
rect 2971 146147 8259 146175
rect 8287 146147 8321 146175
rect 8349 146147 18117 146175
rect 18145 146147 18179 146175
rect 18207 146147 18241 146175
rect 18269 146147 18303 146175
rect 18331 146147 23619 146175
rect 23647 146147 23681 146175
rect 23709 146147 33477 146175
rect 33505 146147 33539 146175
rect 33567 146147 33601 146175
rect 33629 146147 33663 146175
rect 33691 146147 38979 146175
rect 39007 146147 39041 146175
rect 39069 146147 48837 146175
rect 48865 146147 48899 146175
rect 48927 146147 48961 146175
rect 48989 146147 49023 146175
rect 49051 146147 54339 146175
rect 54367 146147 54401 146175
rect 54429 146147 64197 146175
rect 64225 146147 64259 146175
rect 64287 146147 64321 146175
rect 64349 146147 64383 146175
rect 64411 146147 69699 146175
rect 69727 146147 69761 146175
rect 69789 146147 79557 146175
rect 79585 146147 79619 146175
rect 79647 146147 79681 146175
rect 79709 146147 79743 146175
rect 79771 146147 85059 146175
rect 85087 146147 85121 146175
rect 85149 146147 94917 146175
rect 94945 146147 94979 146175
rect 95007 146147 95041 146175
rect 95069 146147 95103 146175
rect 95131 146147 100419 146175
rect 100447 146147 100481 146175
rect 100509 146147 110277 146175
rect 110305 146147 110339 146175
rect 110367 146147 110401 146175
rect 110429 146147 110463 146175
rect 110491 146147 115779 146175
rect 115807 146147 115841 146175
rect 115869 146147 125637 146175
rect 125665 146147 125699 146175
rect 125727 146147 125761 146175
rect 125789 146147 125823 146175
rect 125851 146147 131139 146175
rect 131167 146147 131201 146175
rect 131229 146147 140997 146175
rect 141025 146147 141059 146175
rect 141087 146147 141121 146175
rect 141149 146147 141183 146175
rect 141211 146147 146499 146175
rect 146527 146147 146561 146175
rect 146589 146147 156357 146175
rect 156385 146147 156419 146175
rect 156447 146147 156481 146175
rect 156509 146147 156543 146175
rect 156571 146147 161859 146175
rect 161887 146147 161921 146175
rect 161949 146147 171717 146175
rect 171745 146147 171779 146175
rect 171807 146147 171841 146175
rect 171869 146147 171903 146175
rect 171931 146147 177219 146175
rect 177247 146147 177281 146175
rect 177309 146147 187077 146175
rect 187105 146147 187139 146175
rect 187167 146147 187201 146175
rect 187229 146147 187263 146175
rect 187291 146147 192579 146175
rect 192607 146147 192641 146175
rect 192669 146147 202437 146175
rect 202465 146147 202499 146175
rect 202527 146147 202561 146175
rect 202589 146147 202623 146175
rect 202651 146147 207939 146175
rect 207967 146147 208001 146175
rect 208029 146147 217797 146175
rect 217825 146147 217859 146175
rect 217887 146147 217921 146175
rect 217949 146147 217983 146175
rect 218011 146147 223299 146175
rect 223327 146147 223361 146175
rect 223389 146147 233157 146175
rect 233185 146147 233219 146175
rect 233247 146147 233281 146175
rect 233309 146147 233343 146175
rect 233371 146147 238659 146175
rect 238687 146147 238721 146175
rect 238749 146147 248517 146175
rect 248545 146147 248579 146175
rect 248607 146147 248641 146175
rect 248669 146147 248703 146175
rect 248731 146147 254019 146175
rect 254047 146147 254081 146175
rect 254109 146147 263877 146175
rect 263905 146147 263939 146175
rect 263967 146147 264001 146175
rect 264029 146147 264063 146175
rect 264091 146147 269379 146175
rect 269407 146147 269441 146175
rect 269469 146147 279237 146175
rect 279265 146147 279299 146175
rect 279327 146147 279361 146175
rect 279389 146147 279423 146175
rect 279451 146147 284739 146175
rect 284767 146147 284801 146175
rect 284829 146147 294597 146175
rect 294625 146147 294659 146175
rect 294687 146147 294721 146175
rect 294749 146147 294783 146175
rect 294811 146147 298248 146175
rect 298276 146147 298310 146175
rect 298338 146147 298372 146175
rect 298400 146147 298434 146175
rect 298462 146147 298990 146175
rect -958 146113 298990 146147
rect -958 146085 -430 146113
rect -402 146085 -368 146113
rect -340 146085 -306 146113
rect -278 146085 -244 146113
rect -216 146085 2757 146113
rect 2785 146085 2819 146113
rect 2847 146085 2881 146113
rect 2909 146085 2943 146113
rect 2971 146085 8259 146113
rect 8287 146085 8321 146113
rect 8349 146085 18117 146113
rect 18145 146085 18179 146113
rect 18207 146085 18241 146113
rect 18269 146085 18303 146113
rect 18331 146085 23619 146113
rect 23647 146085 23681 146113
rect 23709 146085 33477 146113
rect 33505 146085 33539 146113
rect 33567 146085 33601 146113
rect 33629 146085 33663 146113
rect 33691 146085 38979 146113
rect 39007 146085 39041 146113
rect 39069 146085 48837 146113
rect 48865 146085 48899 146113
rect 48927 146085 48961 146113
rect 48989 146085 49023 146113
rect 49051 146085 54339 146113
rect 54367 146085 54401 146113
rect 54429 146085 64197 146113
rect 64225 146085 64259 146113
rect 64287 146085 64321 146113
rect 64349 146085 64383 146113
rect 64411 146085 69699 146113
rect 69727 146085 69761 146113
rect 69789 146085 79557 146113
rect 79585 146085 79619 146113
rect 79647 146085 79681 146113
rect 79709 146085 79743 146113
rect 79771 146085 85059 146113
rect 85087 146085 85121 146113
rect 85149 146085 94917 146113
rect 94945 146085 94979 146113
rect 95007 146085 95041 146113
rect 95069 146085 95103 146113
rect 95131 146085 100419 146113
rect 100447 146085 100481 146113
rect 100509 146085 110277 146113
rect 110305 146085 110339 146113
rect 110367 146085 110401 146113
rect 110429 146085 110463 146113
rect 110491 146085 115779 146113
rect 115807 146085 115841 146113
rect 115869 146085 125637 146113
rect 125665 146085 125699 146113
rect 125727 146085 125761 146113
rect 125789 146085 125823 146113
rect 125851 146085 131139 146113
rect 131167 146085 131201 146113
rect 131229 146085 140997 146113
rect 141025 146085 141059 146113
rect 141087 146085 141121 146113
rect 141149 146085 141183 146113
rect 141211 146085 146499 146113
rect 146527 146085 146561 146113
rect 146589 146085 156357 146113
rect 156385 146085 156419 146113
rect 156447 146085 156481 146113
rect 156509 146085 156543 146113
rect 156571 146085 161859 146113
rect 161887 146085 161921 146113
rect 161949 146085 171717 146113
rect 171745 146085 171779 146113
rect 171807 146085 171841 146113
rect 171869 146085 171903 146113
rect 171931 146085 177219 146113
rect 177247 146085 177281 146113
rect 177309 146085 187077 146113
rect 187105 146085 187139 146113
rect 187167 146085 187201 146113
rect 187229 146085 187263 146113
rect 187291 146085 192579 146113
rect 192607 146085 192641 146113
rect 192669 146085 202437 146113
rect 202465 146085 202499 146113
rect 202527 146085 202561 146113
rect 202589 146085 202623 146113
rect 202651 146085 207939 146113
rect 207967 146085 208001 146113
rect 208029 146085 217797 146113
rect 217825 146085 217859 146113
rect 217887 146085 217921 146113
rect 217949 146085 217983 146113
rect 218011 146085 223299 146113
rect 223327 146085 223361 146113
rect 223389 146085 233157 146113
rect 233185 146085 233219 146113
rect 233247 146085 233281 146113
rect 233309 146085 233343 146113
rect 233371 146085 238659 146113
rect 238687 146085 238721 146113
rect 238749 146085 248517 146113
rect 248545 146085 248579 146113
rect 248607 146085 248641 146113
rect 248669 146085 248703 146113
rect 248731 146085 254019 146113
rect 254047 146085 254081 146113
rect 254109 146085 263877 146113
rect 263905 146085 263939 146113
rect 263967 146085 264001 146113
rect 264029 146085 264063 146113
rect 264091 146085 269379 146113
rect 269407 146085 269441 146113
rect 269469 146085 279237 146113
rect 279265 146085 279299 146113
rect 279327 146085 279361 146113
rect 279389 146085 279423 146113
rect 279451 146085 284739 146113
rect 284767 146085 284801 146113
rect 284829 146085 294597 146113
rect 294625 146085 294659 146113
rect 294687 146085 294721 146113
rect 294749 146085 294783 146113
rect 294811 146085 298248 146113
rect 298276 146085 298310 146113
rect 298338 146085 298372 146113
rect 298400 146085 298434 146113
rect 298462 146085 298990 146113
rect -958 146051 298990 146085
rect -958 146023 -430 146051
rect -402 146023 -368 146051
rect -340 146023 -306 146051
rect -278 146023 -244 146051
rect -216 146023 2757 146051
rect 2785 146023 2819 146051
rect 2847 146023 2881 146051
rect 2909 146023 2943 146051
rect 2971 146023 8259 146051
rect 8287 146023 8321 146051
rect 8349 146023 18117 146051
rect 18145 146023 18179 146051
rect 18207 146023 18241 146051
rect 18269 146023 18303 146051
rect 18331 146023 23619 146051
rect 23647 146023 23681 146051
rect 23709 146023 33477 146051
rect 33505 146023 33539 146051
rect 33567 146023 33601 146051
rect 33629 146023 33663 146051
rect 33691 146023 38979 146051
rect 39007 146023 39041 146051
rect 39069 146023 48837 146051
rect 48865 146023 48899 146051
rect 48927 146023 48961 146051
rect 48989 146023 49023 146051
rect 49051 146023 54339 146051
rect 54367 146023 54401 146051
rect 54429 146023 64197 146051
rect 64225 146023 64259 146051
rect 64287 146023 64321 146051
rect 64349 146023 64383 146051
rect 64411 146023 69699 146051
rect 69727 146023 69761 146051
rect 69789 146023 79557 146051
rect 79585 146023 79619 146051
rect 79647 146023 79681 146051
rect 79709 146023 79743 146051
rect 79771 146023 85059 146051
rect 85087 146023 85121 146051
rect 85149 146023 94917 146051
rect 94945 146023 94979 146051
rect 95007 146023 95041 146051
rect 95069 146023 95103 146051
rect 95131 146023 100419 146051
rect 100447 146023 100481 146051
rect 100509 146023 110277 146051
rect 110305 146023 110339 146051
rect 110367 146023 110401 146051
rect 110429 146023 110463 146051
rect 110491 146023 115779 146051
rect 115807 146023 115841 146051
rect 115869 146023 125637 146051
rect 125665 146023 125699 146051
rect 125727 146023 125761 146051
rect 125789 146023 125823 146051
rect 125851 146023 131139 146051
rect 131167 146023 131201 146051
rect 131229 146023 140997 146051
rect 141025 146023 141059 146051
rect 141087 146023 141121 146051
rect 141149 146023 141183 146051
rect 141211 146023 146499 146051
rect 146527 146023 146561 146051
rect 146589 146023 156357 146051
rect 156385 146023 156419 146051
rect 156447 146023 156481 146051
rect 156509 146023 156543 146051
rect 156571 146023 161859 146051
rect 161887 146023 161921 146051
rect 161949 146023 171717 146051
rect 171745 146023 171779 146051
rect 171807 146023 171841 146051
rect 171869 146023 171903 146051
rect 171931 146023 177219 146051
rect 177247 146023 177281 146051
rect 177309 146023 187077 146051
rect 187105 146023 187139 146051
rect 187167 146023 187201 146051
rect 187229 146023 187263 146051
rect 187291 146023 192579 146051
rect 192607 146023 192641 146051
rect 192669 146023 202437 146051
rect 202465 146023 202499 146051
rect 202527 146023 202561 146051
rect 202589 146023 202623 146051
rect 202651 146023 207939 146051
rect 207967 146023 208001 146051
rect 208029 146023 217797 146051
rect 217825 146023 217859 146051
rect 217887 146023 217921 146051
rect 217949 146023 217983 146051
rect 218011 146023 223299 146051
rect 223327 146023 223361 146051
rect 223389 146023 233157 146051
rect 233185 146023 233219 146051
rect 233247 146023 233281 146051
rect 233309 146023 233343 146051
rect 233371 146023 238659 146051
rect 238687 146023 238721 146051
rect 238749 146023 248517 146051
rect 248545 146023 248579 146051
rect 248607 146023 248641 146051
rect 248669 146023 248703 146051
rect 248731 146023 254019 146051
rect 254047 146023 254081 146051
rect 254109 146023 263877 146051
rect 263905 146023 263939 146051
rect 263967 146023 264001 146051
rect 264029 146023 264063 146051
rect 264091 146023 269379 146051
rect 269407 146023 269441 146051
rect 269469 146023 279237 146051
rect 279265 146023 279299 146051
rect 279327 146023 279361 146051
rect 279389 146023 279423 146051
rect 279451 146023 284739 146051
rect 284767 146023 284801 146051
rect 284829 146023 294597 146051
rect 294625 146023 294659 146051
rect 294687 146023 294721 146051
rect 294749 146023 294783 146051
rect 294811 146023 298248 146051
rect 298276 146023 298310 146051
rect 298338 146023 298372 146051
rect 298400 146023 298434 146051
rect 298462 146023 298990 146051
rect -958 145989 298990 146023
rect -958 145961 -430 145989
rect -402 145961 -368 145989
rect -340 145961 -306 145989
rect -278 145961 -244 145989
rect -216 145961 2757 145989
rect 2785 145961 2819 145989
rect 2847 145961 2881 145989
rect 2909 145961 2943 145989
rect 2971 145961 8259 145989
rect 8287 145961 8321 145989
rect 8349 145961 18117 145989
rect 18145 145961 18179 145989
rect 18207 145961 18241 145989
rect 18269 145961 18303 145989
rect 18331 145961 23619 145989
rect 23647 145961 23681 145989
rect 23709 145961 33477 145989
rect 33505 145961 33539 145989
rect 33567 145961 33601 145989
rect 33629 145961 33663 145989
rect 33691 145961 38979 145989
rect 39007 145961 39041 145989
rect 39069 145961 48837 145989
rect 48865 145961 48899 145989
rect 48927 145961 48961 145989
rect 48989 145961 49023 145989
rect 49051 145961 54339 145989
rect 54367 145961 54401 145989
rect 54429 145961 64197 145989
rect 64225 145961 64259 145989
rect 64287 145961 64321 145989
rect 64349 145961 64383 145989
rect 64411 145961 69699 145989
rect 69727 145961 69761 145989
rect 69789 145961 79557 145989
rect 79585 145961 79619 145989
rect 79647 145961 79681 145989
rect 79709 145961 79743 145989
rect 79771 145961 85059 145989
rect 85087 145961 85121 145989
rect 85149 145961 94917 145989
rect 94945 145961 94979 145989
rect 95007 145961 95041 145989
rect 95069 145961 95103 145989
rect 95131 145961 100419 145989
rect 100447 145961 100481 145989
rect 100509 145961 110277 145989
rect 110305 145961 110339 145989
rect 110367 145961 110401 145989
rect 110429 145961 110463 145989
rect 110491 145961 115779 145989
rect 115807 145961 115841 145989
rect 115869 145961 125637 145989
rect 125665 145961 125699 145989
rect 125727 145961 125761 145989
rect 125789 145961 125823 145989
rect 125851 145961 131139 145989
rect 131167 145961 131201 145989
rect 131229 145961 140997 145989
rect 141025 145961 141059 145989
rect 141087 145961 141121 145989
rect 141149 145961 141183 145989
rect 141211 145961 146499 145989
rect 146527 145961 146561 145989
rect 146589 145961 156357 145989
rect 156385 145961 156419 145989
rect 156447 145961 156481 145989
rect 156509 145961 156543 145989
rect 156571 145961 161859 145989
rect 161887 145961 161921 145989
rect 161949 145961 171717 145989
rect 171745 145961 171779 145989
rect 171807 145961 171841 145989
rect 171869 145961 171903 145989
rect 171931 145961 177219 145989
rect 177247 145961 177281 145989
rect 177309 145961 187077 145989
rect 187105 145961 187139 145989
rect 187167 145961 187201 145989
rect 187229 145961 187263 145989
rect 187291 145961 192579 145989
rect 192607 145961 192641 145989
rect 192669 145961 202437 145989
rect 202465 145961 202499 145989
rect 202527 145961 202561 145989
rect 202589 145961 202623 145989
rect 202651 145961 207939 145989
rect 207967 145961 208001 145989
rect 208029 145961 217797 145989
rect 217825 145961 217859 145989
rect 217887 145961 217921 145989
rect 217949 145961 217983 145989
rect 218011 145961 223299 145989
rect 223327 145961 223361 145989
rect 223389 145961 233157 145989
rect 233185 145961 233219 145989
rect 233247 145961 233281 145989
rect 233309 145961 233343 145989
rect 233371 145961 238659 145989
rect 238687 145961 238721 145989
rect 238749 145961 248517 145989
rect 248545 145961 248579 145989
rect 248607 145961 248641 145989
rect 248669 145961 248703 145989
rect 248731 145961 254019 145989
rect 254047 145961 254081 145989
rect 254109 145961 263877 145989
rect 263905 145961 263939 145989
rect 263967 145961 264001 145989
rect 264029 145961 264063 145989
rect 264091 145961 269379 145989
rect 269407 145961 269441 145989
rect 269469 145961 279237 145989
rect 279265 145961 279299 145989
rect 279327 145961 279361 145989
rect 279389 145961 279423 145989
rect 279451 145961 284739 145989
rect 284767 145961 284801 145989
rect 284829 145961 294597 145989
rect 294625 145961 294659 145989
rect 294687 145961 294721 145989
rect 294749 145961 294783 145989
rect 294811 145961 298248 145989
rect 298276 145961 298310 145989
rect 298338 145961 298372 145989
rect 298400 145961 298434 145989
rect 298462 145961 298990 145989
rect -958 145913 298990 145961
rect -958 140175 298990 140223
rect -958 140147 -910 140175
rect -882 140147 -848 140175
rect -820 140147 -786 140175
rect -758 140147 -724 140175
rect -696 140147 4617 140175
rect 4645 140147 4679 140175
rect 4707 140147 4741 140175
rect 4769 140147 4803 140175
rect 4831 140147 15939 140175
rect 15967 140147 16001 140175
rect 16029 140147 19977 140175
rect 20005 140147 20039 140175
rect 20067 140147 20101 140175
rect 20129 140147 20163 140175
rect 20191 140147 31299 140175
rect 31327 140147 31361 140175
rect 31389 140147 35337 140175
rect 35365 140147 35399 140175
rect 35427 140147 35461 140175
rect 35489 140147 35523 140175
rect 35551 140147 46659 140175
rect 46687 140147 46721 140175
rect 46749 140147 50697 140175
rect 50725 140147 50759 140175
rect 50787 140147 50821 140175
rect 50849 140147 50883 140175
rect 50911 140147 62019 140175
rect 62047 140147 62081 140175
rect 62109 140147 66057 140175
rect 66085 140147 66119 140175
rect 66147 140147 66181 140175
rect 66209 140147 66243 140175
rect 66271 140147 77379 140175
rect 77407 140147 77441 140175
rect 77469 140147 81417 140175
rect 81445 140147 81479 140175
rect 81507 140147 81541 140175
rect 81569 140147 81603 140175
rect 81631 140147 92739 140175
rect 92767 140147 92801 140175
rect 92829 140147 96777 140175
rect 96805 140147 96839 140175
rect 96867 140147 96901 140175
rect 96929 140147 96963 140175
rect 96991 140147 108099 140175
rect 108127 140147 108161 140175
rect 108189 140147 112137 140175
rect 112165 140147 112199 140175
rect 112227 140147 112261 140175
rect 112289 140147 112323 140175
rect 112351 140147 123459 140175
rect 123487 140147 123521 140175
rect 123549 140147 127497 140175
rect 127525 140147 127559 140175
rect 127587 140147 127621 140175
rect 127649 140147 127683 140175
rect 127711 140147 138819 140175
rect 138847 140147 138881 140175
rect 138909 140147 142857 140175
rect 142885 140147 142919 140175
rect 142947 140147 142981 140175
rect 143009 140147 143043 140175
rect 143071 140147 154179 140175
rect 154207 140147 154241 140175
rect 154269 140147 158217 140175
rect 158245 140147 158279 140175
rect 158307 140147 158341 140175
rect 158369 140147 158403 140175
rect 158431 140147 169539 140175
rect 169567 140147 169601 140175
rect 169629 140147 173577 140175
rect 173605 140147 173639 140175
rect 173667 140147 173701 140175
rect 173729 140147 173763 140175
rect 173791 140147 184899 140175
rect 184927 140147 184961 140175
rect 184989 140147 188937 140175
rect 188965 140147 188999 140175
rect 189027 140147 189061 140175
rect 189089 140147 189123 140175
rect 189151 140147 200259 140175
rect 200287 140147 200321 140175
rect 200349 140147 204297 140175
rect 204325 140147 204359 140175
rect 204387 140147 204421 140175
rect 204449 140147 204483 140175
rect 204511 140147 215619 140175
rect 215647 140147 215681 140175
rect 215709 140147 219657 140175
rect 219685 140147 219719 140175
rect 219747 140147 219781 140175
rect 219809 140147 219843 140175
rect 219871 140147 230979 140175
rect 231007 140147 231041 140175
rect 231069 140147 235017 140175
rect 235045 140147 235079 140175
rect 235107 140147 235141 140175
rect 235169 140147 235203 140175
rect 235231 140147 246339 140175
rect 246367 140147 246401 140175
rect 246429 140147 250377 140175
rect 250405 140147 250439 140175
rect 250467 140147 250501 140175
rect 250529 140147 250563 140175
rect 250591 140147 261699 140175
rect 261727 140147 261761 140175
rect 261789 140147 265737 140175
rect 265765 140147 265799 140175
rect 265827 140147 265861 140175
rect 265889 140147 265923 140175
rect 265951 140147 277059 140175
rect 277087 140147 277121 140175
rect 277149 140147 281097 140175
rect 281125 140147 281159 140175
rect 281187 140147 281221 140175
rect 281249 140147 281283 140175
rect 281311 140147 296457 140175
rect 296485 140147 296519 140175
rect 296547 140147 296581 140175
rect 296609 140147 296643 140175
rect 296671 140147 298728 140175
rect 298756 140147 298790 140175
rect 298818 140147 298852 140175
rect 298880 140147 298914 140175
rect 298942 140147 298990 140175
rect -958 140113 298990 140147
rect -958 140085 -910 140113
rect -882 140085 -848 140113
rect -820 140085 -786 140113
rect -758 140085 -724 140113
rect -696 140085 4617 140113
rect 4645 140085 4679 140113
rect 4707 140085 4741 140113
rect 4769 140085 4803 140113
rect 4831 140085 15939 140113
rect 15967 140085 16001 140113
rect 16029 140085 19977 140113
rect 20005 140085 20039 140113
rect 20067 140085 20101 140113
rect 20129 140085 20163 140113
rect 20191 140085 31299 140113
rect 31327 140085 31361 140113
rect 31389 140085 35337 140113
rect 35365 140085 35399 140113
rect 35427 140085 35461 140113
rect 35489 140085 35523 140113
rect 35551 140085 46659 140113
rect 46687 140085 46721 140113
rect 46749 140085 50697 140113
rect 50725 140085 50759 140113
rect 50787 140085 50821 140113
rect 50849 140085 50883 140113
rect 50911 140085 62019 140113
rect 62047 140085 62081 140113
rect 62109 140085 66057 140113
rect 66085 140085 66119 140113
rect 66147 140085 66181 140113
rect 66209 140085 66243 140113
rect 66271 140085 77379 140113
rect 77407 140085 77441 140113
rect 77469 140085 81417 140113
rect 81445 140085 81479 140113
rect 81507 140085 81541 140113
rect 81569 140085 81603 140113
rect 81631 140085 92739 140113
rect 92767 140085 92801 140113
rect 92829 140085 96777 140113
rect 96805 140085 96839 140113
rect 96867 140085 96901 140113
rect 96929 140085 96963 140113
rect 96991 140085 108099 140113
rect 108127 140085 108161 140113
rect 108189 140085 112137 140113
rect 112165 140085 112199 140113
rect 112227 140085 112261 140113
rect 112289 140085 112323 140113
rect 112351 140085 123459 140113
rect 123487 140085 123521 140113
rect 123549 140085 127497 140113
rect 127525 140085 127559 140113
rect 127587 140085 127621 140113
rect 127649 140085 127683 140113
rect 127711 140085 138819 140113
rect 138847 140085 138881 140113
rect 138909 140085 142857 140113
rect 142885 140085 142919 140113
rect 142947 140085 142981 140113
rect 143009 140085 143043 140113
rect 143071 140085 154179 140113
rect 154207 140085 154241 140113
rect 154269 140085 158217 140113
rect 158245 140085 158279 140113
rect 158307 140085 158341 140113
rect 158369 140085 158403 140113
rect 158431 140085 169539 140113
rect 169567 140085 169601 140113
rect 169629 140085 173577 140113
rect 173605 140085 173639 140113
rect 173667 140085 173701 140113
rect 173729 140085 173763 140113
rect 173791 140085 184899 140113
rect 184927 140085 184961 140113
rect 184989 140085 188937 140113
rect 188965 140085 188999 140113
rect 189027 140085 189061 140113
rect 189089 140085 189123 140113
rect 189151 140085 200259 140113
rect 200287 140085 200321 140113
rect 200349 140085 204297 140113
rect 204325 140085 204359 140113
rect 204387 140085 204421 140113
rect 204449 140085 204483 140113
rect 204511 140085 215619 140113
rect 215647 140085 215681 140113
rect 215709 140085 219657 140113
rect 219685 140085 219719 140113
rect 219747 140085 219781 140113
rect 219809 140085 219843 140113
rect 219871 140085 230979 140113
rect 231007 140085 231041 140113
rect 231069 140085 235017 140113
rect 235045 140085 235079 140113
rect 235107 140085 235141 140113
rect 235169 140085 235203 140113
rect 235231 140085 246339 140113
rect 246367 140085 246401 140113
rect 246429 140085 250377 140113
rect 250405 140085 250439 140113
rect 250467 140085 250501 140113
rect 250529 140085 250563 140113
rect 250591 140085 261699 140113
rect 261727 140085 261761 140113
rect 261789 140085 265737 140113
rect 265765 140085 265799 140113
rect 265827 140085 265861 140113
rect 265889 140085 265923 140113
rect 265951 140085 277059 140113
rect 277087 140085 277121 140113
rect 277149 140085 281097 140113
rect 281125 140085 281159 140113
rect 281187 140085 281221 140113
rect 281249 140085 281283 140113
rect 281311 140085 296457 140113
rect 296485 140085 296519 140113
rect 296547 140085 296581 140113
rect 296609 140085 296643 140113
rect 296671 140085 298728 140113
rect 298756 140085 298790 140113
rect 298818 140085 298852 140113
rect 298880 140085 298914 140113
rect 298942 140085 298990 140113
rect -958 140051 298990 140085
rect -958 140023 -910 140051
rect -882 140023 -848 140051
rect -820 140023 -786 140051
rect -758 140023 -724 140051
rect -696 140023 4617 140051
rect 4645 140023 4679 140051
rect 4707 140023 4741 140051
rect 4769 140023 4803 140051
rect 4831 140023 15939 140051
rect 15967 140023 16001 140051
rect 16029 140023 19977 140051
rect 20005 140023 20039 140051
rect 20067 140023 20101 140051
rect 20129 140023 20163 140051
rect 20191 140023 31299 140051
rect 31327 140023 31361 140051
rect 31389 140023 35337 140051
rect 35365 140023 35399 140051
rect 35427 140023 35461 140051
rect 35489 140023 35523 140051
rect 35551 140023 46659 140051
rect 46687 140023 46721 140051
rect 46749 140023 50697 140051
rect 50725 140023 50759 140051
rect 50787 140023 50821 140051
rect 50849 140023 50883 140051
rect 50911 140023 62019 140051
rect 62047 140023 62081 140051
rect 62109 140023 66057 140051
rect 66085 140023 66119 140051
rect 66147 140023 66181 140051
rect 66209 140023 66243 140051
rect 66271 140023 77379 140051
rect 77407 140023 77441 140051
rect 77469 140023 81417 140051
rect 81445 140023 81479 140051
rect 81507 140023 81541 140051
rect 81569 140023 81603 140051
rect 81631 140023 92739 140051
rect 92767 140023 92801 140051
rect 92829 140023 96777 140051
rect 96805 140023 96839 140051
rect 96867 140023 96901 140051
rect 96929 140023 96963 140051
rect 96991 140023 108099 140051
rect 108127 140023 108161 140051
rect 108189 140023 112137 140051
rect 112165 140023 112199 140051
rect 112227 140023 112261 140051
rect 112289 140023 112323 140051
rect 112351 140023 123459 140051
rect 123487 140023 123521 140051
rect 123549 140023 127497 140051
rect 127525 140023 127559 140051
rect 127587 140023 127621 140051
rect 127649 140023 127683 140051
rect 127711 140023 138819 140051
rect 138847 140023 138881 140051
rect 138909 140023 142857 140051
rect 142885 140023 142919 140051
rect 142947 140023 142981 140051
rect 143009 140023 143043 140051
rect 143071 140023 154179 140051
rect 154207 140023 154241 140051
rect 154269 140023 158217 140051
rect 158245 140023 158279 140051
rect 158307 140023 158341 140051
rect 158369 140023 158403 140051
rect 158431 140023 169539 140051
rect 169567 140023 169601 140051
rect 169629 140023 173577 140051
rect 173605 140023 173639 140051
rect 173667 140023 173701 140051
rect 173729 140023 173763 140051
rect 173791 140023 184899 140051
rect 184927 140023 184961 140051
rect 184989 140023 188937 140051
rect 188965 140023 188999 140051
rect 189027 140023 189061 140051
rect 189089 140023 189123 140051
rect 189151 140023 200259 140051
rect 200287 140023 200321 140051
rect 200349 140023 204297 140051
rect 204325 140023 204359 140051
rect 204387 140023 204421 140051
rect 204449 140023 204483 140051
rect 204511 140023 215619 140051
rect 215647 140023 215681 140051
rect 215709 140023 219657 140051
rect 219685 140023 219719 140051
rect 219747 140023 219781 140051
rect 219809 140023 219843 140051
rect 219871 140023 230979 140051
rect 231007 140023 231041 140051
rect 231069 140023 235017 140051
rect 235045 140023 235079 140051
rect 235107 140023 235141 140051
rect 235169 140023 235203 140051
rect 235231 140023 246339 140051
rect 246367 140023 246401 140051
rect 246429 140023 250377 140051
rect 250405 140023 250439 140051
rect 250467 140023 250501 140051
rect 250529 140023 250563 140051
rect 250591 140023 261699 140051
rect 261727 140023 261761 140051
rect 261789 140023 265737 140051
rect 265765 140023 265799 140051
rect 265827 140023 265861 140051
rect 265889 140023 265923 140051
rect 265951 140023 277059 140051
rect 277087 140023 277121 140051
rect 277149 140023 281097 140051
rect 281125 140023 281159 140051
rect 281187 140023 281221 140051
rect 281249 140023 281283 140051
rect 281311 140023 296457 140051
rect 296485 140023 296519 140051
rect 296547 140023 296581 140051
rect 296609 140023 296643 140051
rect 296671 140023 298728 140051
rect 298756 140023 298790 140051
rect 298818 140023 298852 140051
rect 298880 140023 298914 140051
rect 298942 140023 298990 140051
rect -958 139989 298990 140023
rect -958 139961 -910 139989
rect -882 139961 -848 139989
rect -820 139961 -786 139989
rect -758 139961 -724 139989
rect -696 139961 4617 139989
rect 4645 139961 4679 139989
rect 4707 139961 4741 139989
rect 4769 139961 4803 139989
rect 4831 139961 15939 139989
rect 15967 139961 16001 139989
rect 16029 139961 19977 139989
rect 20005 139961 20039 139989
rect 20067 139961 20101 139989
rect 20129 139961 20163 139989
rect 20191 139961 31299 139989
rect 31327 139961 31361 139989
rect 31389 139961 35337 139989
rect 35365 139961 35399 139989
rect 35427 139961 35461 139989
rect 35489 139961 35523 139989
rect 35551 139961 46659 139989
rect 46687 139961 46721 139989
rect 46749 139961 50697 139989
rect 50725 139961 50759 139989
rect 50787 139961 50821 139989
rect 50849 139961 50883 139989
rect 50911 139961 62019 139989
rect 62047 139961 62081 139989
rect 62109 139961 66057 139989
rect 66085 139961 66119 139989
rect 66147 139961 66181 139989
rect 66209 139961 66243 139989
rect 66271 139961 77379 139989
rect 77407 139961 77441 139989
rect 77469 139961 81417 139989
rect 81445 139961 81479 139989
rect 81507 139961 81541 139989
rect 81569 139961 81603 139989
rect 81631 139961 92739 139989
rect 92767 139961 92801 139989
rect 92829 139961 96777 139989
rect 96805 139961 96839 139989
rect 96867 139961 96901 139989
rect 96929 139961 96963 139989
rect 96991 139961 108099 139989
rect 108127 139961 108161 139989
rect 108189 139961 112137 139989
rect 112165 139961 112199 139989
rect 112227 139961 112261 139989
rect 112289 139961 112323 139989
rect 112351 139961 123459 139989
rect 123487 139961 123521 139989
rect 123549 139961 127497 139989
rect 127525 139961 127559 139989
rect 127587 139961 127621 139989
rect 127649 139961 127683 139989
rect 127711 139961 138819 139989
rect 138847 139961 138881 139989
rect 138909 139961 142857 139989
rect 142885 139961 142919 139989
rect 142947 139961 142981 139989
rect 143009 139961 143043 139989
rect 143071 139961 154179 139989
rect 154207 139961 154241 139989
rect 154269 139961 158217 139989
rect 158245 139961 158279 139989
rect 158307 139961 158341 139989
rect 158369 139961 158403 139989
rect 158431 139961 169539 139989
rect 169567 139961 169601 139989
rect 169629 139961 173577 139989
rect 173605 139961 173639 139989
rect 173667 139961 173701 139989
rect 173729 139961 173763 139989
rect 173791 139961 184899 139989
rect 184927 139961 184961 139989
rect 184989 139961 188937 139989
rect 188965 139961 188999 139989
rect 189027 139961 189061 139989
rect 189089 139961 189123 139989
rect 189151 139961 200259 139989
rect 200287 139961 200321 139989
rect 200349 139961 204297 139989
rect 204325 139961 204359 139989
rect 204387 139961 204421 139989
rect 204449 139961 204483 139989
rect 204511 139961 215619 139989
rect 215647 139961 215681 139989
rect 215709 139961 219657 139989
rect 219685 139961 219719 139989
rect 219747 139961 219781 139989
rect 219809 139961 219843 139989
rect 219871 139961 230979 139989
rect 231007 139961 231041 139989
rect 231069 139961 235017 139989
rect 235045 139961 235079 139989
rect 235107 139961 235141 139989
rect 235169 139961 235203 139989
rect 235231 139961 246339 139989
rect 246367 139961 246401 139989
rect 246429 139961 250377 139989
rect 250405 139961 250439 139989
rect 250467 139961 250501 139989
rect 250529 139961 250563 139989
rect 250591 139961 261699 139989
rect 261727 139961 261761 139989
rect 261789 139961 265737 139989
rect 265765 139961 265799 139989
rect 265827 139961 265861 139989
rect 265889 139961 265923 139989
rect 265951 139961 277059 139989
rect 277087 139961 277121 139989
rect 277149 139961 281097 139989
rect 281125 139961 281159 139989
rect 281187 139961 281221 139989
rect 281249 139961 281283 139989
rect 281311 139961 296457 139989
rect 296485 139961 296519 139989
rect 296547 139961 296581 139989
rect 296609 139961 296643 139989
rect 296671 139961 298728 139989
rect 298756 139961 298790 139989
rect 298818 139961 298852 139989
rect 298880 139961 298914 139989
rect 298942 139961 298990 139989
rect -958 139913 298990 139961
rect -958 137175 298990 137223
rect -958 137147 -430 137175
rect -402 137147 -368 137175
rect -340 137147 -306 137175
rect -278 137147 -244 137175
rect -216 137147 2757 137175
rect 2785 137147 2819 137175
rect 2847 137147 2881 137175
rect 2909 137147 2943 137175
rect 2971 137147 8259 137175
rect 8287 137147 8321 137175
rect 8349 137147 18117 137175
rect 18145 137147 18179 137175
rect 18207 137147 18241 137175
rect 18269 137147 18303 137175
rect 18331 137147 23619 137175
rect 23647 137147 23681 137175
rect 23709 137147 33477 137175
rect 33505 137147 33539 137175
rect 33567 137147 33601 137175
rect 33629 137147 33663 137175
rect 33691 137147 38979 137175
rect 39007 137147 39041 137175
rect 39069 137147 48837 137175
rect 48865 137147 48899 137175
rect 48927 137147 48961 137175
rect 48989 137147 49023 137175
rect 49051 137147 54339 137175
rect 54367 137147 54401 137175
rect 54429 137147 64197 137175
rect 64225 137147 64259 137175
rect 64287 137147 64321 137175
rect 64349 137147 64383 137175
rect 64411 137147 69699 137175
rect 69727 137147 69761 137175
rect 69789 137147 79557 137175
rect 79585 137147 79619 137175
rect 79647 137147 79681 137175
rect 79709 137147 79743 137175
rect 79771 137147 85059 137175
rect 85087 137147 85121 137175
rect 85149 137147 94917 137175
rect 94945 137147 94979 137175
rect 95007 137147 95041 137175
rect 95069 137147 95103 137175
rect 95131 137147 100419 137175
rect 100447 137147 100481 137175
rect 100509 137147 110277 137175
rect 110305 137147 110339 137175
rect 110367 137147 110401 137175
rect 110429 137147 110463 137175
rect 110491 137147 115779 137175
rect 115807 137147 115841 137175
rect 115869 137147 125637 137175
rect 125665 137147 125699 137175
rect 125727 137147 125761 137175
rect 125789 137147 125823 137175
rect 125851 137147 131139 137175
rect 131167 137147 131201 137175
rect 131229 137147 140997 137175
rect 141025 137147 141059 137175
rect 141087 137147 141121 137175
rect 141149 137147 141183 137175
rect 141211 137147 146499 137175
rect 146527 137147 146561 137175
rect 146589 137147 156357 137175
rect 156385 137147 156419 137175
rect 156447 137147 156481 137175
rect 156509 137147 156543 137175
rect 156571 137147 161859 137175
rect 161887 137147 161921 137175
rect 161949 137147 171717 137175
rect 171745 137147 171779 137175
rect 171807 137147 171841 137175
rect 171869 137147 171903 137175
rect 171931 137147 177219 137175
rect 177247 137147 177281 137175
rect 177309 137147 187077 137175
rect 187105 137147 187139 137175
rect 187167 137147 187201 137175
rect 187229 137147 187263 137175
rect 187291 137147 192579 137175
rect 192607 137147 192641 137175
rect 192669 137147 202437 137175
rect 202465 137147 202499 137175
rect 202527 137147 202561 137175
rect 202589 137147 202623 137175
rect 202651 137147 207939 137175
rect 207967 137147 208001 137175
rect 208029 137147 217797 137175
rect 217825 137147 217859 137175
rect 217887 137147 217921 137175
rect 217949 137147 217983 137175
rect 218011 137147 223299 137175
rect 223327 137147 223361 137175
rect 223389 137147 233157 137175
rect 233185 137147 233219 137175
rect 233247 137147 233281 137175
rect 233309 137147 233343 137175
rect 233371 137147 238659 137175
rect 238687 137147 238721 137175
rect 238749 137147 248517 137175
rect 248545 137147 248579 137175
rect 248607 137147 248641 137175
rect 248669 137147 248703 137175
rect 248731 137147 254019 137175
rect 254047 137147 254081 137175
rect 254109 137147 263877 137175
rect 263905 137147 263939 137175
rect 263967 137147 264001 137175
rect 264029 137147 264063 137175
rect 264091 137147 269379 137175
rect 269407 137147 269441 137175
rect 269469 137147 279237 137175
rect 279265 137147 279299 137175
rect 279327 137147 279361 137175
rect 279389 137147 279423 137175
rect 279451 137147 284739 137175
rect 284767 137147 284801 137175
rect 284829 137147 294597 137175
rect 294625 137147 294659 137175
rect 294687 137147 294721 137175
rect 294749 137147 294783 137175
rect 294811 137147 298248 137175
rect 298276 137147 298310 137175
rect 298338 137147 298372 137175
rect 298400 137147 298434 137175
rect 298462 137147 298990 137175
rect -958 137113 298990 137147
rect -958 137085 -430 137113
rect -402 137085 -368 137113
rect -340 137085 -306 137113
rect -278 137085 -244 137113
rect -216 137085 2757 137113
rect 2785 137085 2819 137113
rect 2847 137085 2881 137113
rect 2909 137085 2943 137113
rect 2971 137085 8259 137113
rect 8287 137085 8321 137113
rect 8349 137085 18117 137113
rect 18145 137085 18179 137113
rect 18207 137085 18241 137113
rect 18269 137085 18303 137113
rect 18331 137085 23619 137113
rect 23647 137085 23681 137113
rect 23709 137085 33477 137113
rect 33505 137085 33539 137113
rect 33567 137085 33601 137113
rect 33629 137085 33663 137113
rect 33691 137085 38979 137113
rect 39007 137085 39041 137113
rect 39069 137085 48837 137113
rect 48865 137085 48899 137113
rect 48927 137085 48961 137113
rect 48989 137085 49023 137113
rect 49051 137085 54339 137113
rect 54367 137085 54401 137113
rect 54429 137085 64197 137113
rect 64225 137085 64259 137113
rect 64287 137085 64321 137113
rect 64349 137085 64383 137113
rect 64411 137085 69699 137113
rect 69727 137085 69761 137113
rect 69789 137085 79557 137113
rect 79585 137085 79619 137113
rect 79647 137085 79681 137113
rect 79709 137085 79743 137113
rect 79771 137085 85059 137113
rect 85087 137085 85121 137113
rect 85149 137085 94917 137113
rect 94945 137085 94979 137113
rect 95007 137085 95041 137113
rect 95069 137085 95103 137113
rect 95131 137085 100419 137113
rect 100447 137085 100481 137113
rect 100509 137085 110277 137113
rect 110305 137085 110339 137113
rect 110367 137085 110401 137113
rect 110429 137085 110463 137113
rect 110491 137085 115779 137113
rect 115807 137085 115841 137113
rect 115869 137085 125637 137113
rect 125665 137085 125699 137113
rect 125727 137085 125761 137113
rect 125789 137085 125823 137113
rect 125851 137085 131139 137113
rect 131167 137085 131201 137113
rect 131229 137085 140997 137113
rect 141025 137085 141059 137113
rect 141087 137085 141121 137113
rect 141149 137085 141183 137113
rect 141211 137085 146499 137113
rect 146527 137085 146561 137113
rect 146589 137085 156357 137113
rect 156385 137085 156419 137113
rect 156447 137085 156481 137113
rect 156509 137085 156543 137113
rect 156571 137085 161859 137113
rect 161887 137085 161921 137113
rect 161949 137085 171717 137113
rect 171745 137085 171779 137113
rect 171807 137085 171841 137113
rect 171869 137085 171903 137113
rect 171931 137085 177219 137113
rect 177247 137085 177281 137113
rect 177309 137085 187077 137113
rect 187105 137085 187139 137113
rect 187167 137085 187201 137113
rect 187229 137085 187263 137113
rect 187291 137085 192579 137113
rect 192607 137085 192641 137113
rect 192669 137085 202437 137113
rect 202465 137085 202499 137113
rect 202527 137085 202561 137113
rect 202589 137085 202623 137113
rect 202651 137085 207939 137113
rect 207967 137085 208001 137113
rect 208029 137085 217797 137113
rect 217825 137085 217859 137113
rect 217887 137085 217921 137113
rect 217949 137085 217983 137113
rect 218011 137085 223299 137113
rect 223327 137085 223361 137113
rect 223389 137085 233157 137113
rect 233185 137085 233219 137113
rect 233247 137085 233281 137113
rect 233309 137085 233343 137113
rect 233371 137085 238659 137113
rect 238687 137085 238721 137113
rect 238749 137085 248517 137113
rect 248545 137085 248579 137113
rect 248607 137085 248641 137113
rect 248669 137085 248703 137113
rect 248731 137085 254019 137113
rect 254047 137085 254081 137113
rect 254109 137085 263877 137113
rect 263905 137085 263939 137113
rect 263967 137085 264001 137113
rect 264029 137085 264063 137113
rect 264091 137085 269379 137113
rect 269407 137085 269441 137113
rect 269469 137085 279237 137113
rect 279265 137085 279299 137113
rect 279327 137085 279361 137113
rect 279389 137085 279423 137113
rect 279451 137085 284739 137113
rect 284767 137085 284801 137113
rect 284829 137085 294597 137113
rect 294625 137085 294659 137113
rect 294687 137085 294721 137113
rect 294749 137085 294783 137113
rect 294811 137085 298248 137113
rect 298276 137085 298310 137113
rect 298338 137085 298372 137113
rect 298400 137085 298434 137113
rect 298462 137085 298990 137113
rect -958 137051 298990 137085
rect -958 137023 -430 137051
rect -402 137023 -368 137051
rect -340 137023 -306 137051
rect -278 137023 -244 137051
rect -216 137023 2757 137051
rect 2785 137023 2819 137051
rect 2847 137023 2881 137051
rect 2909 137023 2943 137051
rect 2971 137023 8259 137051
rect 8287 137023 8321 137051
rect 8349 137023 18117 137051
rect 18145 137023 18179 137051
rect 18207 137023 18241 137051
rect 18269 137023 18303 137051
rect 18331 137023 23619 137051
rect 23647 137023 23681 137051
rect 23709 137023 33477 137051
rect 33505 137023 33539 137051
rect 33567 137023 33601 137051
rect 33629 137023 33663 137051
rect 33691 137023 38979 137051
rect 39007 137023 39041 137051
rect 39069 137023 48837 137051
rect 48865 137023 48899 137051
rect 48927 137023 48961 137051
rect 48989 137023 49023 137051
rect 49051 137023 54339 137051
rect 54367 137023 54401 137051
rect 54429 137023 64197 137051
rect 64225 137023 64259 137051
rect 64287 137023 64321 137051
rect 64349 137023 64383 137051
rect 64411 137023 69699 137051
rect 69727 137023 69761 137051
rect 69789 137023 79557 137051
rect 79585 137023 79619 137051
rect 79647 137023 79681 137051
rect 79709 137023 79743 137051
rect 79771 137023 85059 137051
rect 85087 137023 85121 137051
rect 85149 137023 94917 137051
rect 94945 137023 94979 137051
rect 95007 137023 95041 137051
rect 95069 137023 95103 137051
rect 95131 137023 100419 137051
rect 100447 137023 100481 137051
rect 100509 137023 110277 137051
rect 110305 137023 110339 137051
rect 110367 137023 110401 137051
rect 110429 137023 110463 137051
rect 110491 137023 115779 137051
rect 115807 137023 115841 137051
rect 115869 137023 125637 137051
rect 125665 137023 125699 137051
rect 125727 137023 125761 137051
rect 125789 137023 125823 137051
rect 125851 137023 131139 137051
rect 131167 137023 131201 137051
rect 131229 137023 140997 137051
rect 141025 137023 141059 137051
rect 141087 137023 141121 137051
rect 141149 137023 141183 137051
rect 141211 137023 146499 137051
rect 146527 137023 146561 137051
rect 146589 137023 156357 137051
rect 156385 137023 156419 137051
rect 156447 137023 156481 137051
rect 156509 137023 156543 137051
rect 156571 137023 161859 137051
rect 161887 137023 161921 137051
rect 161949 137023 171717 137051
rect 171745 137023 171779 137051
rect 171807 137023 171841 137051
rect 171869 137023 171903 137051
rect 171931 137023 177219 137051
rect 177247 137023 177281 137051
rect 177309 137023 187077 137051
rect 187105 137023 187139 137051
rect 187167 137023 187201 137051
rect 187229 137023 187263 137051
rect 187291 137023 192579 137051
rect 192607 137023 192641 137051
rect 192669 137023 202437 137051
rect 202465 137023 202499 137051
rect 202527 137023 202561 137051
rect 202589 137023 202623 137051
rect 202651 137023 207939 137051
rect 207967 137023 208001 137051
rect 208029 137023 217797 137051
rect 217825 137023 217859 137051
rect 217887 137023 217921 137051
rect 217949 137023 217983 137051
rect 218011 137023 223299 137051
rect 223327 137023 223361 137051
rect 223389 137023 233157 137051
rect 233185 137023 233219 137051
rect 233247 137023 233281 137051
rect 233309 137023 233343 137051
rect 233371 137023 238659 137051
rect 238687 137023 238721 137051
rect 238749 137023 248517 137051
rect 248545 137023 248579 137051
rect 248607 137023 248641 137051
rect 248669 137023 248703 137051
rect 248731 137023 254019 137051
rect 254047 137023 254081 137051
rect 254109 137023 263877 137051
rect 263905 137023 263939 137051
rect 263967 137023 264001 137051
rect 264029 137023 264063 137051
rect 264091 137023 269379 137051
rect 269407 137023 269441 137051
rect 269469 137023 279237 137051
rect 279265 137023 279299 137051
rect 279327 137023 279361 137051
rect 279389 137023 279423 137051
rect 279451 137023 284739 137051
rect 284767 137023 284801 137051
rect 284829 137023 294597 137051
rect 294625 137023 294659 137051
rect 294687 137023 294721 137051
rect 294749 137023 294783 137051
rect 294811 137023 298248 137051
rect 298276 137023 298310 137051
rect 298338 137023 298372 137051
rect 298400 137023 298434 137051
rect 298462 137023 298990 137051
rect -958 136989 298990 137023
rect -958 136961 -430 136989
rect -402 136961 -368 136989
rect -340 136961 -306 136989
rect -278 136961 -244 136989
rect -216 136961 2757 136989
rect 2785 136961 2819 136989
rect 2847 136961 2881 136989
rect 2909 136961 2943 136989
rect 2971 136961 8259 136989
rect 8287 136961 8321 136989
rect 8349 136961 18117 136989
rect 18145 136961 18179 136989
rect 18207 136961 18241 136989
rect 18269 136961 18303 136989
rect 18331 136961 23619 136989
rect 23647 136961 23681 136989
rect 23709 136961 33477 136989
rect 33505 136961 33539 136989
rect 33567 136961 33601 136989
rect 33629 136961 33663 136989
rect 33691 136961 38979 136989
rect 39007 136961 39041 136989
rect 39069 136961 48837 136989
rect 48865 136961 48899 136989
rect 48927 136961 48961 136989
rect 48989 136961 49023 136989
rect 49051 136961 54339 136989
rect 54367 136961 54401 136989
rect 54429 136961 64197 136989
rect 64225 136961 64259 136989
rect 64287 136961 64321 136989
rect 64349 136961 64383 136989
rect 64411 136961 69699 136989
rect 69727 136961 69761 136989
rect 69789 136961 79557 136989
rect 79585 136961 79619 136989
rect 79647 136961 79681 136989
rect 79709 136961 79743 136989
rect 79771 136961 85059 136989
rect 85087 136961 85121 136989
rect 85149 136961 94917 136989
rect 94945 136961 94979 136989
rect 95007 136961 95041 136989
rect 95069 136961 95103 136989
rect 95131 136961 100419 136989
rect 100447 136961 100481 136989
rect 100509 136961 110277 136989
rect 110305 136961 110339 136989
rect 110367 136961 110401 136989
rect 110429 136961 110463 136989
rect 110491 136961 115779 136989
rect 115807 136961 115841 136989
rect 115869 136961 125637 136989
rect 125665 136961 125699 136989
rect 125727 136961 125761 136989
rect 125789 136961 125823 136989
rect 125851 136961 131139 136989
rect 131167 136961 131201 136989
rect 131229 136961 140997 136989
rect 141025 136961 141059 136989
rect 141087 136961 141121 136989
rect 141149 136961 141183 136989
rect 141211 136961 146499 136989
rect 146527 136961 146561 136989
rect 146589 136961 156357 136989
rect 156385 136961 156419 136989
rect 156447 136961 156481 136989
rect 156509 136961 156543 136989
rect 156571 136961 161859 136989
rect 161887 136961 161921 136989
rect 161949 136961 171717 136989
rect 171745 136961 171779 136989
rect 171807 136961 171841 136989
rect 171869 136961 171903 136989
rect 171931 136961 177219 136989
rect 177247 136961 177281 136989
rect 177309 136961 187077 136989
rect 187105 136961 187139 136989
rect 187167 136961 187201 136989
rect 187229 136961 187263 136989
rect 187291 136961 192579 136989
rect 192607 136961 192641 136989
rect 192669 136961 202437 136989
rect 202465 136961 202499 136989
rect 202527 136961 202561 136989
rect 202589 136961 202623 136989
rect 202651 136961 207939 136989
rect 207967 136961 208001 136989
rect 208029 136961 217797 136989
rect 217825 136961 217859 136989
rect 217887 136961 217921 136989
rect 217949 136961 217983 136989
rect 218011 136961 223299 136989
rect 223327 136961 223361 136989
rect 223389 136961 233157 136989
rect 233185 136961 233219 136989
rect 233247 136961 233281 136989
rect 233309 136961 233343 136989
rect 233371 136961 238659 136989
rect 238687 136961 238721 136989
rect 238749 136961 248517 136989
rect 248545 136961 248579 136989
rect 248607 136961 248641 136989
rect 248669 136961 248703 136989
rect 248731 136961 254019 136989
rect 254047 136961 254081 136989
rect 254109 136961 263877 136989
rect 263905 136961 263939 136989
rect 263967 136961 264001 136989
rect 264029 136961 264063 136989
rect 264091 136961 269379 136989
rect 269407 136961 269441 136989
rect 269469 136961 279237 136989
rect 279265 136961 279299 136989
rect 279327 136961 279361 136989
rect 279389 136961 279423 136989
rect 279451 136961 284739 136989
rect 284767 136961 284801 136989
rect 284829 136961 294597 136989
rect 294625 136961 294659 136989
rect 294687 136961 294721 136989
rect 294749 136961 294783 136989
rect 294811 136961 298248 136989
rect 298276 136961 298310 136989
rect 298338 136961 298372 136989
rect 298400 136961 298434 136989
rect 298462 136961 298990 136989
rect -958 136913 298990 136961
rect -958 131175 298990 131223
rect -958 131147 -910 131175
rect -882 131147 -848 131175
rect -820 131147 -786 131175
rect -758 131147 -724 131175
rect -696 131147 4617 131175
rect 4645 131147 4679 131175
rect 4707 131147 4741 131175
rect 4769 131147 4803 131175
rect 4831 131147 15939 131175
rect 15967 131147 16001 131175
rect 16029 131147 19977 131175
rect 20005 131147 20039 131175
rect 20067 131147 20101 131175
rect 20129 131147 20163 131175
rect 20191 131147 31299 131175
rect 31327 131147 31361 131175
rect 31389 131147 35337 131175
rect 35365 131147 35399 131175
rect 35427 131147 35461 131175
rect 35489 131147 35523 131175
rect 35551 131147 46659 131175
rect 46687 131147 46721 131175
rect 46749 131147 50697 131175
rect 50725 131147 50759 131175
rect 50787 131147 50821 131175
rect 50849 131147 50883 131175
rect 50911 131147 62019 131175
rect 62047 131147 62081 131175
rect 62109 131147 66057 131175
rect 66085 131147 66119 131175
rect 66147 131147 66181 131175
rect 66209 131147 66243 131175
rect 66271 131147 77379 131175
rect 77407 131147 77441 131175
rect 77469 131147 81417 131175
rect 81445 131147 81479 131175
rect 81507 131147 81541 131175
rect 81569 131147 81603 131175
rect 81631 131147 92739 131175
rect 92767 131147 92801 131175
rect 92829 131147 96777 131175
rect 96805 131147 96839 131175
rect 96867 131147 96901 131175
rect 96929 131147 96963 131175
rect 96991 131147 108099 131175
rect 108127 131147 108161 131175
rect 108189 131147 112137 131175
rect 112165 131147 112199 131175
rect 112227 131147 112261 131175
rect 112289 131147 112323 131175
rect 112351 131147 123459 131175
rect 123487 131147 123521 131175
rect 123549 131147 127497 131175
rect 127525 131147 127559 131175
rect 127587 131147 127621 131175
rect 127649 131147 127683 131175
rect 127711 131147 138819 131175
rect 138847 131147 138881 131175
rect 138909 131147 142857 131175
rect 142885 131147 142919 131175
rect 142947 131147 142981 131175
rect 143009 131147 143043 131175
rect 143071 131147 154179 131175
rect 154207 131147 154241 131175
rect 154269 131147 158217 131175
rect 158245 131147 158279 131175
rect 158307 131147 158341 131175
rect 158369 131147 158403 131175
rect 158431 131147 169539 131175
rect 169567 131147 169601 131175
rect 169629 131147 173577 131175
rect 173605 131147 173639 131175
rect 173667 131147 173701 131175
rect 173729 131147 173763 131175
rect 173791 131147 184899 131175
rect 184927 131147 184961 131175
rect 184989 131147 188937 131175
rect 188965 131147 188999 131175
rect 189027 131147 189061 131175
rect 189089 131147 189123 131175
rect 189151 131147 200259 131175
rect 200287 131147 200321 131175
rect 200349 131147 204297 131175
rect 204325 131147 204359 131175
rect 204387 131147 204421 131175
rect 204449 131147 204483 131175
rect 204511 131147 215619 131175
rect 215647 131147 215681 131175
rect 215709 131147 219657 131175
rect 219685 131147 219719 131175
rect 219747 131147 219781 131175
rect 219809 131147 219843 131175
rect 219871 131147 230979 131175
rect 231007 131147 231041 131175
rect 231069 131147 235017 131175
rect 235045 131147 235079 131175
rect 235107 131147 235141 131175
rect 235169 131147 235203 131175
rect 235231 131147 246339 131175
rect 246367 131147 246401 131175
rect 246429 131147 250377 131175
rect 250405 131147 250439 131175
rect 250467 131147 250501 131175
rect 250529 131147 250563 131175
rect 250591 131147 261699 131175
rect 261727 131147 261761 131175
rect 261789 131147 265737 131175
rect 265765 131147 265799 131175
rect 265827 131147 265861 131175
rect 265889 131147 265923 131175
rect 265951 131147 277059 131175
rect 277087 131147 277121 131175
rect 277149 131147 281097 131175
rect 281125 131147 281159 131175
rect 281187 131147 281221 131175
rect 281249 131147 281283 131175
rect 281311 131147 296457 131175
rect 296485 131147 296519 131175
rect 296547 131147 296581 131175
rect 296609 131147 296643 131175
rect 296671 131147 298728 131175
rect 298756 131147 298790 131175
rect 298818 131147 298852 131175
rect 298880 131147 298914 131175
rect 298942 131147 298990 131175
rect -958 131113 298990 131147
rect -958 131085 -910 131113
rect -882 131085 -848 131113
rect -820 131085 -786 131113
rect -758 131085 -724 131113
rect -696 131085 4617 131113
rect 4645 131085 4679 131113
rect 4707 131085 4741 131113
rect 4769 131085 4803 131113
rect 4831 131085 15939 131113
rect 15967 131085 16001 131113
rect 16029 131085 19977 131113
rect 20005 131085 20039 131113
rect 20067 131085 20101 131113
rect 20129 131085 20163 131113
rect 20191 131085 31299 131113
rect 31327 131085 31361 131113
rect 31389 131085 35337 131113
rect 35365 131085 35399 131113
rect 35427 131085 35461 131113
rect 35489 131085 35523 131113
rect 35551 131085 46659 131113
rect 46687 131085 46721 131113
rect 46749 131085 50697 131113
rect 50725 131085 50759 131113
rect 50787 131085 50821 131113
rect 50849 131085 50883 131113
rect 50911 131085 62019 131113
rect 62047 131085 62081 131113
rect 62109 131085 66057 131113
rect 66085 131085 66119 131113
rect 66147 131085 66181 131113
rect 66209 131085 66243 131113
rect 66271 131085 77379 131113
rect 77407 131085 77441 131113
rect 77469 131085 81417 131113
rect 81445 131085 81479 131113
rect 81507 131085 81541 131113
rect 81569 131085 81603 131113
rect 81631 131085 92739 131113
rect 92767 131085 92801 131113
rect 92829 131085 96777 131113
rect 96805 131085 96839 131113
rect 96867 131085 96901 131113
rect 96929 131085 96963 131113
rect 96991 131085 108099 131113
rect 108127 131085 108161 131113
rect 108189 131085 112137 131113
rect 112165 131085 112199 131113
rect 112227 131085 112261 131113
rect 112289 131085 112323 131113
rect 112351 131085 123459 131113
rect 123487 131085 123521 131113
rect 123549 131085 127497 131113
rect 127525 131085 127559 131113
rect 127587 131085 127621 131113
rect 127649 131085 127683 131113
rect 127711 131085 138819 131113
rect 138847 131085 138881 131113
rect 138909 131085 142857 131113
rect 142885 131085 142919 131113
rect 142947 131085 142981 131113
rect 143009 131085 143043 131113
rect 143071 131085 154179 131113
rect 154207 131085 154241 131113
rect 154269 131085 158217 131113
rect 158245 131085 158279 131113
rect 158307 131085 158341 131113
rect 158369 131085 158403 131113
rect 158431 131085 169539 131113
rect 169567 131085 169601 131113
rect 169629 131085 173577 131113
rect 173605 131085 173639 131113
rect 173667 131085 173701 131113
rect 173729 131085 173763 131113
rect 173791 131085 184899 131113
rect 184927 131085 184961 131113
rect 184989 131085 188937 131113
rect 188965 131085 188999 131113
rect 189027 131085 189061 131113
rect 189089 131085 189123 131113
rect 189151 131085 200259 131113
rect 200287 131085 200321 131113
rect 200349 131085 204297 131113
rect 204325 131085 204359 131113
rect 204387 131085 204421 131113
rect 204449 131085 204483 131113
rect 204511 131085 215619 131113
rect 215647 131085 215681 131113
rect 215709 131085 219657 131113
rect 219685 131085 219719 131113
rect 219747 131085 219781 131113
rect 219809 131085 219843 131113
rect 219871 131085 230979 131113
rect 231007 131085 231041 131113
rect 231069 131085 235017 131113
rect 235045 131085 235079 131113
rect 235107 131085 235141 131113
rect 235169 131085 235203 131113
rect 235231 131085 246339 131113
rect 246367 131085 246401 131113
rect 246429 131085 250377 131113
rect 250405 131085 250439 131113
rect 250467 131085 250501 131113
rect 250529 131085 250563 131113
rect 250591 131085 261699 131113
rect 261727 131085 261761 131113
rect 261789 131085 265737 131113
rect 265765 131085 265799 131113
rect 265827 131085 265861 131113
rect 265889 131085 265923 131113
rect 265951 131085 277059 131113
rect 277087 131085 277121 131113
rect 277149 131085 281097 131113
rect 281125 131085 281159 131113
rect 281187 131085 281221 131113
rect 281249 131085 281283 131113
rect 281311 131085 296457 131113
rect 296485 131085 296519 131113
rect 296547 131085 296581 131113
rect 296609 131085 296643 131113
rect 296671 131085 298728 131113
rect 298756 131085 298790 131113
rect 298818 131085 298852 131113
rect 298880 131085 298914 131113
rect 298942 131085 298990 131113
rect -958 131051 298990 131085
rect -958 131023 -910 131051
rect -882 131023 -848 131051
rect -820 131023 -786 131051
rect -758 131023 -724 131051
rect -696 131023 4617 131051
rect 4645 131023 4679 131051
rect 4707 131023 4741 131051
rect 4769 131023 4803 131051
rect 4831 131023 15939 131051
rect 15967 131023 16001 131051
rect 16029 131023 19977 131051
rect 20005 131023 20039 131051
rect 20067 131023 20101 131051
rect 20129 131023 20163 131051
rect 20191 131023 31299 131051
rect 31327 131023 31361 131051
rect 31389 131023 35337 131051
rect 35365 131023 35399 131051
rect 35427 131023 35461 131051
rect 35489 131023 35523 131051
rect 35551 131023 46659 131051
rect 46687 131023 46721 131051
rect 46749 131023 50697 131051
rect 50725 131023 50759 131051
rect 50787 131023 50821 131051
rect 50849 131023 50883 131051
rect 50911 131023 62019 131051
rect 62047 131023 62081 131051
rect 62109 131023 66057 131051
rect 66085 131023 66119 131051
rect 66147 131023 66181 131051
rect 66209 131023 66243 131051
rect 66271 131023 77379 131051
rect 77407 131023 77441 131051
rect 77469 131023 81417 131051
rect 81445 131023 81479 131051
rect 81507 131023 81541 131051
rect 81569 131023 81603 131051
rect 81631 131023 92739 131051
rect 92767 131023 92801 131051
rect 92829 131023 96777 131051
rect 96805 131023 96839 131051
rect 96867 131023 96901 131051
rect 96929 131023 96963 131051
rect 96991 131023 108099 131051
rect 108127 131023 108161 131051
rect 108189 131023 112137 131051
rect 112165 131023 112199 131051
rect 112227 131023 112261 131051
rect 112289 131023 112323 131051
rect 112351 131023 123459 131051
rect 123487 131023 123521 131051
rect 123549 131023 127497 131051
rect 127525 131023 127559 131051
rect 127587 131023 127621 131051
rect 127649 131023 127683 131051
rect 127711 131023 138819 131051
rect 138847 131023 138881 131051
rect 138909 131023 142857 131051
rect 142885 131023 142919 131051
rect 142947 131023 142981 131051
rect 143009 131023 143043 131051
rect 143071 131023 154179 131051
rect 154207 131023 154241 131051
rect 154269 131023 158217 131051
rect 158245 131023 158279 131051
rect 158307 131023 158341 131051
rect 158369 131023 158403 131051
rect 158431 131023 169539 131051
rect 169567 131023 169601 131051
rect 169629 131023 173577 131051
rect 173605 131023 173639 131051
rect 173667 131023 173701 131051
rect 173729 131023 173763 131051
rect 173791 131023 184899 131051
rect 184927 131023 184961 131051
rect 184989 131023 188937 131051
rect 188965 131023 188999 131051
rect 189027 131023 189061 131051
rect 189089 131023 189123 131051
rect 189151 131023 200259 131051
rect 200287 131023 200321 131051
rect 200349 131023 204297 131051
rect 204325 131023 204359 131051
rect 204387 131023 204421 131051
rect 204449 131023 204483 131051
rect 204511 131023 215619 131051
rect 215647 131023 215681 131051
rect 215709 131023 219657 131051
rect 219685 131023 219719 131051
rect 219747 131023 219781 131051
rect 219809 131023 219843 131051
rect 219871 131023 230979 131051
rect 231007 131023 231041 131051
rect 231069 131023 235017 131051
rect 235045 131023 235079 131051
rect 235107 131023 235141 131051
rect 235169 131023 235203 131051
rect 235231 131023 246339 131051
rect 246367 131023 246401 131051
rect 246429 131023 250377 131051
rect 250405 131023 250439 131051
rect 250467 131023 250501 131051
rect 250529 131023 250563 131051
rect 250591 131023 261699 131051
rect 261727 131023 261761 131051
rect 261789 131023 265737 131051
rect 265765 131023 265799 131051
rect 265827 131023 265861 131051
rect 265889 131023 265923 131051
rect 265951 131023 277059 131051
rect 277087 131023 277121 131051
rect 277149 131023 281097 131051
rect 281125 131023 281159 131051
rect 281187 131023 281221 131051
rect 281249 131023 281283 131051
rect 281311 131023 296457 131051
rect 296485 131023 296519 131051
rect 296547 131023 296581 131051
rect 296609 131023 296643 131051
rect 296671 131023 298728 131051
rect 298756 131023 298790 131051
rect 298818 131023 298852 131051
rect 298880 131023 298914 131051
rect 298942 131023 298990 131051
rect -958 130989 298990 131023
rect -958 130961 -910 130989
rect -882 130961 -848 130989
rect -820 130961 -786 130989
rect -758 130961 -724 130989
rect -696 130961 4617 130989
rect 4645 130961 4679 130989
rect 4707 130961 4741 130989
rect 4769 130961 4803 130989
rect 4831 130961 15939 130989
rect 15967 130961 16001 130989
rect 16029 130961 19977 130989
rect 20005 130961 20039 130989
rect 20067 130961 20101 130989
rect 20129 130961 20163 130989
rect 20191 130961 31299 130989
rect 31327 130961 31361 130989
rect 31389 130961 35337 130989
rect 35365 130961 35399 130989
rect 35427 130961 35461 130989
rect 35489 130961 35523 130989
rect 35551 130961 46659 130989
rect 46687 130961 46721 130989
rect 46749 130961 50697 130989
rect 50725 130961 50759 130989
rect 50787 130961 50821 130989
rect 50849 130961 50883 130989
rect 50911 130961 62019 130989
rect 62047 130961 62081 130989
rect 62109 130961 66057 130989
rect 66085 130961 66119 130989
rect 66147 130961 66181 130989
rect 66209 130961 66243 130989
rect 66271 130961 77379 130989
rect 77407 130961 77441 130989
rect 77469 130961 81417 130989
rect 81445 130961 81479 130989
rect 81507 130961 81541 130989
rect 81569 130961 81603 130989
rect 81631 130961 92739 130989
rect 92767 130961 92801 130989
rect 92829 130961 96777 130989
rect 96805 130961 96839 130989
rect 96867 130961 96901 130989
rect 96929 130961 96963 130989
rect 96991 130961 108099 130989
rect 108127 130961 108161 130989
rect 108189 130961 112137 130989
rect 112165 130961 112199 130989
rect 112227 130961 112261 130989
rect 112289 130961 112323 130989
rect 112351 130961 123459 130989
rect 123487 130961 123521 130989
rect 123549 130961 127497 130989
rect 127525 130961 127559 130989
rect 127587 130961 127621 130989
rect 127649 130961 127683 130989
rect 127711 130961 138819 130989
rect 138847 130961 138881 130989
rect 138909 130961 142857 130989
rect 142885 130961 142919 130989
rect 142947 130961 142981 130989
rect 143009 130961 143043 130989
rect 143071 130961 154179 130989
rect 154207 130961 154241 130989
rect 154269 130961 158217 130989
rect 158245 130961 158279 130989
rect 158307 130961 158341 130989
rect 158369 130961 158403 130989
rect 158431 130961 169539 130989
rect 169567 130961 169601 130989
rect 169629 130961 173577 130989
rect 173605 130961 173639 130989
rect 173667 130961 173701 130989
rect 173729 130961 173763 130989
rect 173791 130961 184899 130989
rect 184927 130961 184961 130989
rect 184989 130961 188937 130989
rect 188965 130961 188999 130989
rect 189027 130961 189061 130989
rect 189089 130961 189123 130989
rect 189151 130961 200259 130989
rect 200287 130961 200321 130989
rect 200349 130961 204297 130989
rect 204325 130961 204359 130989
rect 204387 130961 204421 130989
rect 204449 130961 204483 130989
rect 204511 130961 215619 130989
rect 215647 130961 215681 130989
rect 215709 130961 219657 130989
rect 219685 130961 219719 130989
rect 219747 130961 219781 130989
rect 219809 130961 219843 130989
rect 219871 130961 230979 130989
rect 231007 130961 231041 130989
rect 231069 130961 235017 130989
rect 235045 130961 235079 130989
rect 235107 130961 235141 130989
rect 235169 130961 235203 130989
rect 235231 130961 246339 130989
rect 246367 130961 246401 130989
rect 246429 130961 250377 130989
rect 250405 130961 250439 130989
rect 250467 130961 250501 130989
rect 250529 130961 250563 130989
rect 250591 130961 261699 130989
rect 261727 130961 261761 130989
rect 261789 130961 265737 130989
rect 265765 130961 265799 130989
rect 265827 130961 265861 130989
rect 265889 130961 265923 130989
rect 265951 130961 277059 130989
rect 277087 130961 277121 130989
rect 277149 130961 281097 130989
rect 281125 130961 281159 130989
rect 281187 130961 281221 130989
rect 281249 130961 281283 130989
rect 281311 130961 296457 130989
rect 296485 130961 296519 130989
rect 296547 130961 296581 130989
rect 296609 130961 296643 130989
rect 296671 130961 298728 130989
rect 298756 130961 298790 130989
rect 298818 130961 298852 130989
rect 298880 130961 298914 130989
rect 298942 130961 298990 130989
rect -958 130913 298990 130961
rect -958 128175 298990 128223
rect -958 128147 -430 128175
rect -402 128147 -368 128175
rect -340 128147 -306 128175
rect -278 128147 -244 128175
rect -216 128147 2757 128175
rect 2785 128147 2819 128175
rect 2847 128147 2881 128175
rect 2909 128147 2943 128175
rect 2971 128147 8259 128175
rect 8287 128147 8321 128175
rect 8349 128147 18117 128175
rect 18145 128147 18179 128175
rect 18207 128147 18241 128175
rect 18269 128147 18303 128175
rect 18331 128147 23619 128175
rect 23647 128147 23681 128175
rect 23709 128147 33477 128175
rect 33505 128147 33539 128175
rect 33567 128147 33601 128175
rect 33629 128147 33663 128175
rect 33691 128147 38979 128175
rect 39007 128147 39041 128175
rect 39069 128147 48837 128175
rect 48865 128147 48899 128175
rect 48927 128147 48961 128175
rect 48989 128147 49023 128175
rect 49051 128147 54339 128175
rect 54367 128147 54401 128175
rect 54429 128147 64197 128175
rect 64225 128147 64259 128175
rect 64287 128147 64321 128175
rect 64349 128147 64383 128175
rect 64411 128147 69699 128175
rect 69727 128147 69761 128175
rect 69789 128147 79557 128175
rect 79585 128147 79619 128175
rect 79647 128147 79681 128175
rect 79709 128147 79743 128175
rect 79771 128147 85059 128175
rect 85087 128147 85121 128175
rect 85149 128147 94917 128175
rect 94945 128147 94979 128175
rect 95007 128147 95041 128175
rect 95069 128147 95103 128175
rect 95131 128147 100419 128175
rect 100447 128147 100481 128175
rect 100509 128147 110277 128175
rect 110305 128147 110339 128175
rect 110367 128147 110401 128175
rect 110429 128147 110463 128175
rect 110491 128147 115779 128175
rect 115807 128147 115841 128175
rect 115869 128147 125637 128175
rect 125665 128147 125699 128175
rect 125727 128147 125761 128175
rect 125789 128147 125823 128175
rect 125851 128147 131139 128175
rect 131167 128147 131201 128175
rect 131229 128147 140997 128175
rect 141025 128147 141059 128175
rect 141087 128147 141121 128175
rect 141149 128147 141183 128175
rect 141211 128147 146499 128175
rect 146527 128147 146561 128175
rect 146589 128147 156357 128175
rect 156385 128147 156419 128175
rect 156447 128147 156481 128175
rect 156509 128147 156543 128175
rect 156571 128147 161859 128175
rect 161887 128147 161921 128175
rect 161949 128147 171717 128175
rect 171745 128147 171779 128175
rect 171807 128147 171841 128175
rect 171869 128147 171903 128175
rect 171931 128147 177219 128175
rect 177247 128147 177281 128175
rect 177309 128147 187077 128175
rect 187105 128147 187139 128175
rect 187167 128147 187201 128175
rect 187229 128147 187263 128175
rect 187291 128147 192579 128175
rect 192607 128147 192641 128175
rect 192669 128147 202437 128175
rect 202465 128147 202499 128175
rect 202527 128147 202561 128175
rect 202589 128147 202623 128175
rect 202651 128147 207939 128175
rect 207967 128147 208001 128175
rect 208029 128147 217797 128175
rect 217825 128147 217859 128175
rect 217887 128147 217921 128175
rect 217949 128147 217983 128175
rect 218011 128147 223299 128175
rect 223327 128147 223361 128175
rect 223389 128147 233157 128175
rect 233185 128147 233219 128175
rect 233247 128147 233281 128175
rect 233309 128147 233343 128175
rect 233371 128147 238659 128175
rect 238687 128147 238721 128175
rect 238749 128147 248517 128175
rect 248545 128147 248579 128175
rect 248607 128147 248641 128175
rect 248669 128147 248703 128175
rect 248731 128147 254019 128175
rect 254047 128147 254081 128175
rect 254109 128147 263877 128175
rect 263905 128147 263939 128175
rect 263967 128147 264001 128175
rect 264029 128147 264063 128175
rect 264091 128147 269379 128175
rect 269407 128147 269441 128175
rect 269469 128147 279237 128175
rect 279265 128147 279299 128175
rect 279327 128147 279361 128175
rect 279389 128147 279423 128175
rect 279451 128147 284739 128175
rect 284767 128147 284801 128175
rect 284829 128147 294597 128175
rect 294625 128147 294659 128175
rect 294687 128147 294721 128175
rect 294749 128147 294783 128175
rect 294811 128147 298248 128175
rect 298276 128147 298310 128175
rect 298338 128147 298372 128175
rect 298400 128147 298434 128175
rect 298462 128147 298990 128175
rect -958 128113 298990 128147
rect -958 128085 -430 128113
rect -402 128085 -368 128113
rect -340 128085 -306 128113
rect -278 128085 -244 128113
rect -216 128085 2757 128113
rect 2785 128085 2819 128113
rect 2847 128085 2881 128113
rect 2909 128085 2943 128113
rect 2971 128085 8259 128113
rect 8287 128085 8321 128113
rect 8349 128085 18117 128113
rect 18145 128085 18179 128113
rect 18207 128085 18241 128113
rect 18269 128085 18303 128113
rect 18331 128085 23619 128113
rect 23647 128085 23681 128113
rect 23709 128085 33477 128113
rect 33505 128085 33539 128113
rect 33567 128085 33601 128113
rect 33629 128085 33663 128113
rect 33691 128085 38979 128113
rect 39007 128085 39041 128113
rect 39069 128085 48837 128113
rect 48865 128085 48899 128113
rect 48927 128085 48961 128113
rect 48989 128085 49023 128113
rect 49051 128085 54339 128113
rect 54367 128085 54401 128113
rect 54429 128085 64197 128113
rect 64225 128085 64259 128113
rect 64287 128085 64321 128113
rect 64349 128085 64383 128113
rect 64411 128085 69699 128113
rect 69727 128085 69761 128113
rect 69789 128085 79557 128113
rect 79585 128085 79619 128113
rect 79647 128085 79681 128113
rect 79709 128085 79743 128113
rect 79771 128085 85059 128113
rect 85087 128085 85121 128113
rect 85149 128085 94917 128113
rect 94945 128085 94979 128113
rect 95007 128085 95041 128113
rect 95069 128085 95103 128113
rect 95131 128085 100419 128113
rect 100447 128085 100481 128113
rect 100509 128085 110277 128113
rect 110305 128085 110339 128113
rect 110367 128085 110401 128113
rect 110429 128085 110463 128113
rect 110491 128085 115779 128113
rect 115807 128085 115841 128113
rect 115869 128085 125637 128113
rect 125665 128085 125699 128113
rect 125727 128085 125761 128113
rect 125789 128085 125823 128113
rect 125851 128085 131139 128113
rect 131167 128085 131201 128113
rect 131229 128085 140997 128113
rect 141025 128085 141059 128113
rect 141087 128085 141121 128113
rect 141149 128085 141183 128113
rect 141211 128085 146499 128113
rect 146527 128085 146561 128113
rect 146589 128085 156357 128113
rect 156385 128085 156419 128113
rect 156447 128085 156481 128113
rect 156509 128085 156543 128113
rect 156571 128085 161859 128113
rect 161887 128085 161921 128113
rect 161949 128085 171717 128113
rect 171745 128085 171779 128113
rect 171807 128085 171841 128113
rect 171869 128085 171903 128113
rect 171931 128085 177219 128113
rect 177247 128085 177281 128113
rect 177309 128085 187077 128113
rect 187105 128085 187139 128113
rect 187167 128085 187201 128113
rect 187229 128085 187263 128113
rect 187291 128085 192579 128113
rect 192607 128085 192641 128113
rect 192669 128085 202437 128113
rect 202465 128085 202499 128113
rect 202527 128085 202561 128113
rect 202589 128085 202623 128113
rect 202651 128085 207939 128113
rect 207967 128085 208001 128113
rect 208029 128085 217797 128113
rect 217825 128085 217859 128113
rect 217887 128085 217921 128113
rect 217949 128085 217983 128113
rect 218011 128085 223299 128113
rect 223327 128085 223361 128113
rect 223389 128085 233157 128113
rect 233185 128085 233219 128113
rect 233247 128085 233281 128113
rect 233309 128085 233343 128113
rect 233371 128085 238659 128113
rect 238687 128085 238721 128113
rect 238749 128085 248517 128113
rect 248545 128085 248579 128113
rect 248607 128085 248641 128113
rect 248669 128085 248703 128113
rect 248731 128085 254019 128113
rect 254047 128085 254081 128113
rect 254109 128085 263877 128113
rect 263905 128085 263939 128113
rect 263967 128085 264001 128113
rect 264029 128085 264063 128113
rect 264091 128085 269379 128113
rect 269407 128085 269441 128113
rect 269469 128085 279237 128113
rect 279265 128085 279299 128113
rect 279327 128085 279361 128113
rect 279389 128085 279423 128113
rect 279451 128085 284739 128113
rect 284767 128085 284801 128113
rect 284829 128085 294597 128113
rect 294625 128085 294659 128113
rect 294687 128085 294721 128113
rect 294749 128085 294783 128113
rect 294811 128085 298248 128113
rect 298276 128085 298310 128113
rect 298338 128085 298372 128113
rect 298400 128085 298434 128113
rect 298462 128085 298990 128113
rect -958 128051 298990 128085
rect -958 128023 -430 128051
rect -402 128023 -368 128051
rect -340 128023 -306 128051
rect -278 128023 -244 128051
rect -216 128023 2757 128051
rect 2785 128023 2819 128051
rect 2847 128023 2881 128051
rect 2909 128023 2943 128051
rect 2971 128023 8259 128051
rect 8287 128023 8321 128051
rect 8349 128023 18117 128051
rect 18145 128023 18179 128051
rect 18207 128023 18241 128051
rect 18269 128023 18303 128051
rect 18331 128023 23619 128051
rect 23647 128023 23681 128051
rect 23709 128023 33477 128051
rect 33505 128023 33539 128051
rect 33567 128023 33601 128051
rect 33629 128023 33663 128051
rect 33691 128023 38979 128051
rect 39007 128023 39041 128051
rect 39069 128023 48837 128051
rect 48865 128023 48899 128051
rect 48927 128023 48961 128051
rect 48989 128023 49023 128051
rect 49051 128023 54339 128051
rect 54367 128023 54401 128051
rect 54429 128023 64197 128051
rect 64225 128023 64259 128051
rect 64287 128023 64321 128051
rect 64349 128023 64383 128051
rect 64411 128023 69699 128051
rect 69727 128023 69761 128051
rect 69789 128023 79557 128051
rect 79585 128023 79619 128051
rect 79647 128023 79681 128051
rect 79709 128023 79743 128051
rect 79771 128023 85059 128051
rect 85087 128023 85121 128051
rect 85149 128023 94917 128051
rect 94945 128023 94979 128051
rect 95007 128023 95041 128051
rect 95069 128023 95103 128051
rect 95131 128023 100419 128051
rect 100447 128023 100481 128051
rect 100509 128023 110277 128051
rect 110305 128023 110339 128051
rect 110367 128023 110401 128051
rect 110429 128023 110463 128051
rect 110491 128023 115779 128051
rect 115807 128023 115841 128051
rect 115869 128023 125637 128051
rect 125665 128023 125699 128051
rect 125727 128023 125761 128051
rect 125789 128023 125823 128051
rect 125851 128023 131139 128051
rect 131167 128023 131201 128051
rect 131229 128023 140997 128051
rect 141025 128023 141059 128051
rect 141087 128023 141121 128051
rect 141149 128023 141183 128051
rect 141211 128023 146499 128051
rect 146527 128023 146561 128051
rect 146589 128023 156357 128051
rect 156385 128023 156419 128051
rect 156447 128023 156481 128051
rect 156509 128023 156543 128051
rect 156571 128023 161859 128051
rect 161887 128023 161921 128051
rect 161949 128023 171717 128051
rect 171745 128023 171779 128051
rect 171807 128023 171841 128051
rect 171869 128023 171903 128051
rect 171931 128023 177219 128051
rect 177247 128023 177281 128051
rect 177309 128023 187077 128051
rect 187105 128023 187139 128051
rect 187167 128023 187201 128051
rect 187229 128023 187263 128051
rect 187291 128023 192579 128051
rect 192607 128023 192641 128051
rect 192669 128023 202437 128051
rect 202465 128023 202499 128051
rect 202527 128023 202561 128051
rect 202589 128023 202623 128051
rect 202651 128023 207939 128051
rect 207967 128023 208001 128051
rect 208029 128023 217797 128051
rect 217825 128023 217859 128051
rect 217887 128023 217921 128051
rect 217949 128023 217983 128051
rect 218011 128023 223299 128051
rect 223327 128023 223361 128051
rect 223389 128023 233157 128051
rect 233185 128023 233219 128051
rect 233247 128023 233281 128051
rect 233309 128023 233343 128051
rect 233371 128023 238659 128051
rect 238687 128023 238721 128051
rect 238749 128023 248517 128051
rect 248545 128023 248579 128051
rect 248607 128023 248641 128051
rect 248669 128023 248703 128051
rect 248731 128023 254019 128051
rect 254047 128023 254081 128051
rect 254109 128023 263877 128051
rect 263905 128023 263939 128051
rect 263967 128023 264001 128051
rect 264029 128023 264063 128051
rect 264091 128023 269379 128051
rect 269407 128023 269441 128051
rect 269469 128023 279237 128051
rect 279265 128023 279299 128051
rect 279327 128023 279361 128051
rect 279389 128023 279423 128051
rect 279451 128023 284739 128051
rect 284767 128023 284801 128051
rect 284829 128023 294597 128051
rect 294625 128023 294659 128051
rect 294687 128023 294721 128051
rect 294749 128023 294783 128051
rect 294811 128023 298248 128051
rect 298276 128023 298310 128051
rect 298338 128023 298372 128051
rect 298400 128023 298434 128051
rect 298462 128023 298990 128051
rect -958 127989 298990 128023
rect -958 127961 -430 127989
rect -402 127961 -368 127989
rect -340 127961 -306 127989
rect -278 127961 -244 127989
rect -216 127961 2757 127989
rect 2785 127961 2819 127989
rect 2847 127961 2881 127989
rect 2909 127961 2943 127989
rect 2971 127961 8259 127989
rect 8287 127961 8321 127989
rect 8349 127961 18117 127989
rect 18145 127961 18179 127989
rect 18207 127961 18241 127989
rect 18269 127961 18303 127989
rect 18331 127961 23619 127989
rect 23647 127961 23681 127989
rect 23709 127961 33477 127989
rect 33505 127961 33539 127989
rect 33567 127961 33601 127989
rect 33629 127961 33663 127989
rect 33691 127961 38979 127989
rect 39007 127961 39041 127989
rect 39069 127961 48837 127989
rect 48865 127961 48899 127989
rect 48927 127961 48961 127989
rect 48989 127961 49023 127989
rect 49051 127961 54339 127989
rect 54367 127961 54401 127989
rect 54429 127961 64197 127989
rect 64225 127961 64259 127989
rect 64287 127961 64321 127989
rect 64349 127961 64383 127989
rect 64411 127961 69699 127989
rect 69727 127961 69761 127989
rect 69789 127961 79557 127989
rect 79585 127961 79619 127989
rect 79647 127961 79681 127989
rect 79709 127961 79743 127989
rect 79771 127961 85059 127989
rect 85087 127961 85121 127989
rect 85149 127961 94917 127989
rect 94945 127961 94979 127989
rect 95007 127961 95041 127989
rect 95069 127961 95103 127989
rect 95131 127961 100419 127989
rect 100447 127961 100481 127989
rect 100509 127961 110277 127989
rect 110305 127961 110339 127989
rect 110367 127961 110401 127989
rect 110429 127961 110463 127989
rect 110491 127961 115779 127989
rect 115807 127961 115841 127989
rect 115869 127961 125637 127989
rect 125665 127961 125699 127989
rect 125727 127961 125761 127989
rect 125789 127961 125823 127989
rect 125851 127961 131139 127989
rect 131167 127961 131201 127989
rect 131229 127961 140997 127989
rect 141025 127961 141059 127989
rect 141087 127961 141121 127989
rect 141149 127961 141183 127989
rect 141211 127961 146499 127989
rect 146527 127961 146561 127989
rect 146589 127961 156357 127989
rect 156385 127961 156419 127989
rect 156447 127961 156481 127989
rect 156509 127961 156543 127989
rect 156571 127961 161859 127989
rect 161887 127961 161921 127989
rect 161949 127961 171717 127989
rect 171745 127961 171779 127989
rect 171807 127961 171841 127989
rect 171869 127961 171903 127989
rect 171931 127961 177219 127989
rect 177247 127961 177281 127989
rect 177309 127961 187077 127989
rect 187105 127961 187139 127989
rect 187167 127961 187201 127989
rect 187229 127961 187263 127989
rect 187291 127961 192579 127989
rect 192607 127961 192641 127989
rect 192669 127961 202437 127989
rect 202465 127961 202499 127989
rect 202527 127961 202561 127989
rect 202589 127961 202623 127989
rect 202651 127961 207939 127989
rect 207967 127961 208001 127989
rect 208029 127961 217797 127989
rect 217825 127961 217859 127989
rect 217887 127961 217921 127989
rect 217949 127961 217983 127989
rect 218011 127961 223299 127989
rect 223327 127961 223361 127989
rect 223389 127961 233157 127989
rect 233185 127961 233219 127989
rect 233247 127961 233281 127989
rect 233309 127961 233343 127989
rect 233371 127961 238659 127989
rect 238687 127961 238721 127989
rect 238749 127961 248517 127989
rect 248545 127961 248579 127989
rect 248607 127961 248641 127989
rect 248669 127961 248703 127989
rect 248731 127961 254019 127989
rect 254047 127961 254081 127989
rect 254109 127961 263877 127989
rect 263905 127961 263939 127989
rect 263967 127961 264001 127989
rect 264029 127961 264063 127989
rect 264091 127961 269379 127989
rect 269407 127961 269441 127989
rect 269469 127961 279237 127989
rect 279265 127961 279299 127989
rect 279327 127961 279361 127989
rect 279389 127961 279423 127989
rect 279451 127961 284739 127989
rect 284767 127961 284801 127989
rect 284829 127961 294597 127989
rect 294625 127961 294659 127989
rect 294687 127961 294721 127989
rect 294749 127961 294783 127989
rect 294811 127961 298248 127989
rect 298276 127961 298310 127989
rect 298338 127961 298372 127989
rect 298400 127961 298434 127989
rect 298462 127961 298990 127989
rect -958 127913 298990 127961
rect -958 122175 298990 122223
rect -958 122147 -910 122175
rect -882 122147 -848 122175
rect -820 122147 -786 122175
rect -758 122147 -724 122175
rect -696 122147 4617 122175
rect 4645 122147 4679 122175
rect 4707 122147 4741 122175
rect 4769 122147 4803 122175
rect 4831 122147 15939 122175
rect 15967 122147 16001 122175
rect 16029 122147 19977 122175
rect 20005 122147 20039 122175
rect 20067 122147 20101 122175
rect 20129 122147 20163 122175
rect 20191 122147 31299 122175
rect 31327 122147 31361 122175
rect 31389 122147 35337 122175
rect 35365 122147 35399 122175
rect 35427 122147 35461 122175
rect 35489 122147 35523 122175
rect 35551 122147 46659 122175
rect 46687 122147 46721 122175
rect 46749 122147 50697 122175
rect 50725 122147 50759 122175
rect 50787 122147 50821 122175
rect 50849 122147 50883 122175
rect 50911 122147 62019 122175
rect 62047 122147 62081 122175
rect 62109 122147 66057 122175
rect 66085 122147 66119 122175
rect 66147 122147 66181 122175
rect 66209 122147 66243 122175
rect 66271 122147 77379 122175
rect 77407 122147 77441 122175
rect 77469 122147 81417 122175
rect 81445 122147 81479 122175
rect 81507 122147 81541 122175
rect 81569 122147 81603 122175
rect 81631 122147 92739 122175
rect 92767 122147 92801 122175
rect 92829 122147 96777 122175
rect 96805 122147 96839 122175
rect 96867 122147 96901 122175
rect 96929 122147 96963 122175
rect 96991 122147 108099 122175
rect 108127 122147 108161 122175
rect 108189 122147 112137 122175
rect 112165 122147 112199 122175
rect 112227 122147 112261 122175
rect 112289 122147 112323 122175
rect 112351 122147 123459 122175
rect 123487 122147 123521 122175
rect 123549 122147 127497 122175
rect 127525 122147 127559 122175
rect 127587 122147 127621 122175
rect 127649 122147 127683 122175
rect 127711 122147 138819 122175
rect 138847 122147 138881 122175
rect 138909 122147 142857 122175
rect 142885 122147 142919 122175
rect 142947 122147 142981 122175
rect 143009 122147 143043 122175
rect 143071 122147 154179 122175
rect 154207 122147 154241 122175
rect 154269 122147 158217 122175
rect 158245 122147 158279 122175
rect 158307 122147 158341 122175
rect 158369 122147 158403 122175
rect 158431 122147 169539 122175
rect 169567 122147 169601 122175
rect 169629 122147 173577 122175
rect 173605 122147 173639 122175
rect 173667 122147 173701 122175
rect 173729 122147 173763 122175
rect 173791 122147 184899 122175
rect 184927 122147 184961 122175
rect 184989 122147 188937 122175
rect 188965 122147 188999 122175
rect 189027 122147 189061 122175
rect 189089 122147 189123 122175
rect 189151 122147 200259 122175
rect 200287 122147 200321 122175
rect 200349 122147 204297 122175
rect 204325 122147 204359 122175
rect 204387 122147 204421 122175
rect 204449 122147 204483 122175
rect 204511 122147 215619 122175
rect 215647 122147 215681 122175
rect 215709 122147 219657 122175
rect 219685 122147 219719 122175
rect 219747 122147 219781 122175
rect 219809 122147 219843 122175
rect 219871 122147 230979 122175
rect 231007 122147 231041 122175
rect 231069 122147 235017 122175
rect 235045 122147 235079 122175
rect 235107 122147 235141 122175
rect 235169 122147 235203 122175
rect 235231 122147 246339 122175
rect 246367 122147 246401 122175
rect 246429 122147 250377 122175
rect 250405 122147 250439 122175
rect 250467 122147 250501 122175
rect 250529 122147 250563 122175
rect 250591 122147 261699 122175
rect 261727 122147 261761 122175
rect 261789 122147 265737 122175
rect 265765 122147 265799 122175
rect 265827 122147 265861 122175
rect 265889 122147 265923 122175
rect 265951 122147 277059 122175
rect 277087 122147 277121 122175
rect 277149 122147 281097 122175
rect 281125 122147 281159 122175
rect 281187 122147 281221 122175
rect 281249 122147 281283 122175
rect 281311 122147 296457 122175
rect 296485 122147 296519 122175
rect 296547 122147 296581 122175
rect 296609 122147 296643 122175
rect 296671 122147 298728 122175
rect 298756 122147 298790 122175
rect 298818 122147 298852 122175
rect 298880 122147 298914 122175
rect 298942 122147 298990 122175
rect -958 122113 298990 122147
rect -958 122085 -910 122113
rect -882 122085 -848 122113
rect -820 122085 -786 122113
rect -758 122085 -724 122113
rect -696 122085 4617 122113
rect 4645 122085 4679 122113
rect 4707 122085 4741 122113
rect 4769 122085 4803 122113
rect 4831 122085 15939 122113
rect 15967 122085 16001 122113
rect 16029 122085 19977 122113
rect 20005 122085 20039 122113
rect 20067 122085 20101 122113
rect 20129 122085 20163 122113
rect 20191 122085 31299 122113
rect 31327 122085 31361 122113
rect 31389 122085 35337 122113
rect 35365 122085 35399 122113
rect 35427 122085 35461 122113
rect 35489 122085 35523 122113
rect 35551 122085 46659 122113
rect 46687 122085 46721 122113
rect 46749 122085 50697 122113
rect 50725 122085 50759 122113
rect 50787 122085 50821 122113
rect 50849 122085 50883 122113
rect 50911 122085 62019 122113
rect 62047 122085 62081 122113
rect 62109 122085 66057 122113
rect 66085 122085 66119 122113
rect 66147 122085 66181 122113
rect 66209 122085 66243 122113
rect 66271 122085 77379 122113
rect 77407 122085 77441 122113
rect 77469 122085 81417 122113
rect 81445 122085 81479 122113
rect 81507 122085 81541 122113
rect 81569 122085 81603 122113
rect 81631 122085 92739 122113
rect 92767 122085 92801 122113
rect 92829 122085 96777 122113
rect 96805 122085 96839 122113
rect 96867 122085 96901 122113
rect 96929 122085 96963 122113
rect 96991 122085 108099 122113
rect 108127 122085 108161 122113
rect 108189 122085 112137 122113
rect 112165 122085 112199 122113
rect 112227 122085 112261 122113
rect 112289 122085 112323 122113
rect 112351 122085 123459 122113
rect 123487 122085 123521 122113
rect 123549 122085 127497 122113
rect 127525 122085 127559 122113
rect 127587 122085 127621 122113
rect 127649 122085 127683 122113
rect 127711 122085 138819 122113
rect 138847 122085 138881 122113
rect 138909 122085 142857 122113
rect 142885 122085 142919 122113
rect 142947 122085 142981 122113
rect 143009 122085 143043 122113
rect 143071 122085 154179 122113
rect 154207 122085 154241 122113
rect 154269 122085 158217 122113
rect 158245 122085 158279 122113
rect 158307 122085 158341 122113
rect 158369 122085 158403 122113
rect 158431 122085 169539 122113
rect 169567 122085 169601 122113
rect 169629 122085 173577 122113
rect 173605 122085 173639 122113
rect 173667 122085 173701 122113
rect 173729 122085 173763 122113
rect 173791 122085 184899 122113
rect 184927 122085 184961 122113
rect 184989 122085 188937 122113
rect 188965 122085 188999 122113
rect 189027 122085 189061 122113
rect 189089 122085 189123 122113
rect 189151 122085 200259 122113
rect 200287 122085 200321 122113
rect 200349 122085 204297 122113
rect 204325 122085 204359 122113
rect 204387 122085 204421 122113
rect 204449 122085 204483 122113
rect 204511 122085 215619 122113
rect 215647 122085 215681 122113
rect 215709 122085 219657 122113
rect 219685 122085 219719 122113
rect 219747 122085 219781 122113
rect 219809 122085 219843 122113
rect 219871 122085 230979 122113
rect 231007 122085 231041 122113
rect 231069 122085 235017 122113
rect 235045 122085 235079 122113
rect 235107 122085 235141 122113
rect 235169 122085 235203 122113
rect 235231 122085 246339 122113
rect 246367 122085 246401 122113
rect 246429 122085 250377 122113
rect 250405 122085 250439 122113
rect 250467 122085 250501 122113
rect 250529 122085 250563 122113
rect 250591 122085 261699 122113
rect 261727 122085 261761 122113
rect 261789 122085 265737 122113
rect 265765 122085 265799 122113
rect 265827 122085 265861 122113
rect 265889 122085 265923 122113
rect 265951 122085 277059 122113
rect 277087 122085 277121 122113
rect 277149 122085 281097 122113
rect 281125 122085 281159 122113
rect 281187 122085 281221 122113
rect 281249 122085 281283 122113
rect 281311 122085 296457 122113
rect 296485 122085 296519 122113
rect 296547 122085 296581 122113
rect 296609 122085 296643 122113
rect 296671 122085 298728 122113
rect 298756 122085 298790 122113
rect 298818 122085 298852 122113
rect 298880 122085 298914 122113
rect 298942 122085 298990 122113
rect -958 122051 298990 122085
rect -958 122023 -910 122051
rect -882 122023 -848 122051
rect -820 122023 -786 122051
rect -758 122023 -724 122051
rect -696 122023 4617 122051
rect 4645 122023 4679 122051
rect 4707 122023 4741 122051
rect 4769 122023 4803 122051
rect 4831 122023 15939 122051
rect 15967 122023 16001 122051
rect 16029 122023 19977 122051
rect 20005 122023 20039 122051
rect 20067 122023 20101 122051
rect 20129 122023 20163 122051
rect 20191 122023 31299 122051
rect 31327 122023 31361 122051
rect 31389 122023 35337 122051
rect 35365 122023 35399 122051
rect 35427 122023 35461 122051
rect 35489 122023 35523 122051
rect 35551 122023 46659 122051
rect 46687 122023 46721 122051
rect 46749 122023 50697 122051
rect 50725 122023 50759 122051
rect 50787 122023 50821 122051
rect 50849 122023 50883 122051
rect 50911 122023 62019 122051
rect 62047 122023 62081 122051
rect 62109 122023 66057 122051
rect 66085 122023 66119 122051
rect 66147 122023 66181 122051
rect 66209 122023 66243 122051
rect 66271 122023 77379 122051
rect 77407 122023 77441 122051
rect 77469 122023 81417 122051
rect 81445 122023 81479 122051
rect 81507 122023 81541 122051
rect 81569 122023 81603 122051
rect 81631 122023 92739 122051
rect 92767 122023 92801 122051
rect 92829 122023 96777 122051
rect 96805 122023 96839 122051
rect 96867 122023 96901 122051
rect 96929 122023 96963 122051
rect 96991 122023 108099 122051
rect 108127 122023 108161 122051
rect 108189 122023 112137 122051
rect 112165 122023 112199 122051
rect 112227 122023 112261 122051
rect 112289 122023 112323 122051
rect 112351 122023 123459 122051
rect 123487 122023 123521 122051
rect 123549 122023 127497 122051
rect 127525 122023 127559 122051
rect 127587 122023 127621 122051
rect 127649 122023 127683 122051
rect 127711 122023 138819 122051
rect 138847 122023 138881 122051
rect 138909 122023 142857 122051
rect 142885 122023 142919 122051
rect 142947 122023 142981 122051
rect 143009 122023 143043 122051
rect 143071 122023 154179 122051
rect 154207 122023 154241 122051
rect 154269 122023 158217 122051
rect 158245 122023 158279 122051
rect 158307 122023 158341 122051
rect 158369 122023 158403 122051
rect 158431 122023 169539 122051
rect 169567 122023 169601 122051
rect 169629 122023 173577 122051
rect 173605 122023 173639 122051
rect 173667 122023 173701 122051
rect 173729 122023 173763 122051
rect 173791 122023 184899 122051
rect 184927 122023 184961 122051
rect 184989 122023 188937 122051
rect 188965 122023 188999 122051
rect 189027 122023 189061 122051
rect 189089 122023 189123 122051
rect 189151 122023 200259 122051
rect 200287 122023 200321 122051
rect 200349 122023 204297 122051
rect 204325 122023 204359 122051
rect 204387 122023 204421 122051
rect 204449 122023 204483 122051
rect 204511 122023 215619 122051
rect 215647 122023 215681 122051
rect 215709 122023 219657 122051
rect 219685 122023 219719 122051
rect 219747 122023 219781 122051
rect 219809 122023 219843 122051
rect 219871 122023 230979 122051
rect 231007 122023 231041 122051
rect 231069 122023 235017 122051
rect 235045 122023 235079 122051
rect 235107 122023 235141 122051
rect 235169 122023 235203 122051
rect 235231 122023 246339 122051
rect 246367 122023 246401 122051
rect 246429 122023 250377 122051
rect 250405 122023 250439 122051
rect 250467 122023 250501 122051
rect 250529 122023 250563 122051
rect 250591 122023 261699 122051
rect 261727 122023 261761 122051
rect 261789 122023 265737 122051
rect 265765 122023 265799 122051
rect 265827 122023 265861 122051
rect 265889 122023 265923 122051
rect 265951 122023 277059 122051
rect 277087 122023 277121 122051
rect 277149 122023 281097 122051
rect 281125 122023 281159 122051
rect 281187 122023 281221 122051
rect 281249 122023 281283 122051
rect 281311 122023 296457 122051
rect 296485 122023 296519 122051
rect 296547 122023 296581 122051
rect 296609 122023 296643 122051
rect 296671 122023 298728 122051
rect 298756 122023 298790 122051
rect 298818 122023 298852 122051
rect 298880 122023 298914 122051
rect 298942 122023 298990 122051
rect -958 121989 298990 122023
rect -958 121961 -910 121989
rect -882 121961 -848 121989
rect -820 121961 -786 121989
rect -758 121961 -724 121989
rect -696 121961 4617 121989
rect 4645 121961 4679 121989
rect 4707 121961 4741 121989
rect 4769 121961 4803 121989
rect 4831 121961 15939 121989
rect 15967 121961 16001 121989
rect 16029 121961 19977 121989
rect 20005 121961 20039 121989
rect 20067 121961 20101 121989
rect 20129 121961 20163 121989
rect 20191 121961 31299 121989
rect 31327 121961 31361 121989
rect 31389 121961 35337 121989
rect 35365 121961 35399 121989
rect 35427 121961 35461 121989
rect 35489 121961 35523 121989
rect 35551 121961 46659 121989
rect 46687 121961 46721 121989
rect 46749 121961 50697 121989
rect 50725 121961 50759 121989
rect 50787 121961 50821 121989
rect 50849 121961 50883 121989
rect 50911 121961 62019 121989
rect 62047 121961 62081 121989
rect 62109 121961 66057 121989
rect 66085 121961 66119 121989
rect 66147 121961 66181 121989
rect 66209 121961 66243 121989
rect 66271 121961 77379 121989
rect 77407 121961 77441 121989
rect 77469 121961 81417 121989
rect 81445 121961 81479 121989
rect 81507 121961 81541 121989
rect 81569 121961 81603 121989
rect 81631 121961 92739 121989
rect 92767 121961 92801 121989
rect 92829 121961 96777 121989
rect 96805 121961 96839 121989
rect 96867 121961 96901 121989
rect 96929 121961 96963 121989
rect 96991 121961 108099 121989
rect 108127 121961 108161 121989
rect 108189 121961 112137 121989
rect 112165 121961 112199 121989
rect 112227 121961 112261 121989
rect 112289 121961 112323 121989
rect 112351 121961 123459 121989
rect 123487 121961 123521 121989
rect 123549 121961 127497 121989
rect 127525 121961 127559 121989
rect 127587 121961 127621 121989
rect 127649 121961 127683 121989
rect 127711 121961 138819 121989
rect 138847 121961 138881 121989
rect 138909 121961 142857 121989
rect 142885 121961 142919 121989
rect 142947 121961 142981 121989
rect 143009 121961 143043 121989
rect 143071 121961 154179 121989
rect 154207 121961 154241 121989
rect 154269 121961 158217 121989
rect 158245 121961 158279 121989
rect 158307 121961 158341 121989
rect 158369 121961 158403 121989
rect 158431 121961 169539 121989
rect 169567 121961 169601 121989
rect 169629 121961 173577 121989
rect 173605 121961 173639 121989
rect 173667 121961 173701 121989
rect 173729 121961 173763 121989
rect 173791 121961 184899 121989
rect 184927 121961 184961 121989
rect 184989 121961 188937 121989
rect 188965 121961 188999 121989
rect 189027 121961 189061 121989
rect 189089 121961 189123 121989
rect 189151 121961 200259 121989
rect 200287 121961 200321 121989
rect 200349 121961 204297 121989
rect 204325 121961 204359 121989
rect 204387 121961 204421 121989
rect 204449 121961 204483 121989
rect 204511 121961 215619 121989
rect 215647 121961 215681 121989
rect 215709 121961 219657 121989
rect 219685 121961 219719 121989
rect 219747 121961 219781 121989
rect 219809 121961 219843 121989
rect 219871 121961 230979 121989
rect 231007 121961 231041 121989
rect 231069 121961 235017 121989
rect 235045 121961 235079 121989
rect 235107 121961 235141 121989
rect 235169 121961 235203 121989
rect 235231 121961 246339 121989
rect 246367 121961 246401 121989
rect 246429 121961 250377 121989
rect 250405 121961 250439 121989
rect 250467 121961 250501 121989
rect 250529 121961 250563 121989
rect 250591 121961 261699 121989
rect 261727 121961 261761 121989
rect 261789 121961 265737 121989
rect 265765 121961 265799 121989
rect 265827 121961 265861 121989
rect 265889 121961 265923 121989
rect 265951 121961 277059 121989
rect 277087 121961 277121 121989
rect 277149 121961 281097 121989
rect 281125 121961 281159 121989
rect 281187 121961 281221 121989
rect 281249 121961 281283 121989
rect 281311 121961 296457 121989
rect 296485 121961 296519 121989
rect 296547 121961 296581 121989
rect 296609 121961 296643 121989
rect 296671 121961 298728 121989
rect 298756 121961 298790 121989
rect 298818 121961 298852 121989
rect 298880 121961 298914 121989
rect 298942 121961 298990 121989
rect -958 121913 298990 121961
rect -958 119175 298990 119223
rect -958 119147 -430 119175
rect -402 119147 -368 119175
rect -340 119147 -306 119175
rect -278 119147 -244 119175
rect -216 119147 2757 119175
rect 2785 119147 2819 119175
rect 2847 119147 2881 119175
rect 2909 119147 2943 119175
rect 2971 119147 8259 119175
rect 8287 119147 8321 119175
rect 8349 119147 18117 119175
rect 18145 119147 18179 119175
rect 18207 119147 18241 119175
rect 18269 119147 18303 119175
rect 18331 119147 23619 119175
rect 23647 119147 23681 119175
rect 23709 119147 33477 119175
rect 33505 119147 33539 119175
rect 33567 119147 33601 119175
rect 33629 119147 33663 119175
rect 33691 119147 38979 119175
rect 39007 119147 39041 119175
rect 39069 119147 48837 119175
rect 48865 119147 48899 119175
rect 48927 119147 48961 119175
rect 48989 119147 49023 119175
rect 49051 119147 54339 119175
rect 54367 119147 54401 119175
rect 54429 119147 64197 119175
rect 64225 119147 64259 119175
rect 64287 119147 64321 119175
rect 64349 119147 64383 119175
rect 64411 119147 69699 119175
rect 69727 119147 69761 119175
rect 69789 119147 79557 119175
rect 79585 119147 79619 119175
rect 79647 119147 79681 119175
rect 79709 119147 79743 119175
rect 79771 119147 85059 119175
rect 85087 119147 85121 119175
rect 85149 119147 94917 119175
rect 94945 119147 94979 119175
rect 95007 119147 95041 119175
rect 95069 119147 95103 119175
rect 95131 119147 100419 119175
rect 100447 119147 100481 119175
rect 100509 119147 110277 119175
rect 110305 119147 110339 119175
rect 110367 119147 110401 119175
rect 110429 119147 110463 119175
rect 110491 119147 115779 119175
rect 115807 119147 115841 119175
rect 115869 119147 125637 119175
rect 125665 119147 125699 119175
rect 125727 119147 125761 119175
rect 125789 119147 125823 119175
rect 125851 119147 131139 119175
rect 131167 119147 131201 119175
rect 131229 119147 140997 119175
rect 141025 119147 141059 119175
rect 141087 119147 141121 119175
rect 141149 119147 141183 119175
rect 141211 119147 146499 119175
rect 146527 119147 146561 119175
rect 146589 119147 156357 119175
rect 156385 119147 156419 119175
rect 156447 119147 156481 119175
rect 156509 119147 156543 119175
rect 156571 119147 161859 119175
rect 161887 119147 161921 119175
rect 161949 119147 171717 119175
rect 171745 119147 171779 119175
rect 171807 119147 171841 119175
rect 171869 119147 171903 119175
rect 171931 119147 177219 119175
rect 177247 119147 177281 119175
rect 177309 119147 187077 119175
rect 187105 119147 187139 119175
rect 187167 119147 187201 119175
rect 187229 119147 187263 119175
rect 187291 119147 192579 119175
rect 192607 119147 192641 119175
rect 192669 119147 202437 119175
rect 202465 119147 202499 119175
rect 202527 119147 202561 119175
rect 202589 119147 202623 119175
rect 202651 119147 207939 119175
rect 207967 119147 208001 119175
rect 208029 119147 217797 119175
rect 217825 119147 217859 119175
rect 217887 119147 217921 119175
rect 217949 119147 217983 119175
rect 218011 119147 223299 119175
rect 223327 119147 223361 119175
rect 223389 119147 233157 119175
rect 233185 119147 233219 119175
rect 233247 119147 233281 119175
rect 233309 119147 233343 119175
rect 233371 119147 238659 119175
rect 238687 119147 238721 119175
rect 238749 119147 248517 119175
rect 248545 119147 248579 119175
rect 248607 119147 248641 119175
rect 248669 119147 248703 119175
rect 248731 119147 254019 119175
rect 254047 119147 254081 119175
rect 254109 119147 263877 119175
rect 263905 119147 263939 119175
rect 263967 119147 264001 119175
rect 264029 119147 264063 119175
rect 264091 119147 269379 119175
rect 269407 119147 269441 119175
rect 269469 119147 279237 119175
rect 279265 119147 279299 119175
rect 279327 119147 279361 119175
rect 279389 119147 279423 119175
rect 279451 119147 284739 119175
rect 284767 119147 284801 119175
rect 284829 119147 294597 119175
rect 294625 119147 294659 119175
rect 294687 119147 294721 119175
rect 294749 119147 294783 119175
rect 294811 119147 298248 119175
rect 298276 119147 298310 119175
rect 298338 119147 298372 119175
rect 298400 119147 298434 119175
rect 298462 119147 298990 119175
rect -958 119113 298990 119147
rect -958 119085 -430 119113
rect -402 119085 -368 119113
rect -340 119085 -306 119113
rect -278 119085 -244 119113
rect -216 119085 2757 119113
rect 2785 119085 2819 119113
rect 2847 119085 2881 119113
rect 2909 119085 2943 119113
rect 2971 119085 8259 119113
rect 8287 119085 8321 119113
rect 8349 119085 18117 119113
rect 18145 119085 18179 119113
rect 18207 119085 18241 119113
rect 18269 119085 18303 119113
rect 18331 119085 23619 119113
rect 23647 119085 23681 119113
rect 23709 119085 33477 119113
rect 33505 119085 33539 119113
rect 33567 119085 33601 119113
rect 33629 119085 33663 119113
rect 33691 119085 38979 119113
rect 39007 119085 39041 119113
rect 39069 119085 48837 119113
rect 48865 119085 48899 119113
rect 48927 119085 48961 119113
rect 48989 119085 49023 119113
rect 49051 119085 54339 119113
rect 54367 119085 54401 119113
rect 54429 119085 64197 119113
rect 64225 119085 64259 119113
rect 64287 119085 64321 119113
rect 64349 119085 64383 119113
rect 64411 119085 69699 119113
rect 69727 119085 69761 119113
rect 69789 119085 79557 119113
rect 79585 119085 79619 119113
rect 79647 119085 79681 119113
rect 79709 119085 79743 119113
rect 79771 119085 85059 119113
rect 85087 119085 85121 119113
rect 85149 119085 94917 119113
rect 94945 119085 94979 119113
rect 95007 119085 95041 119113
rect 95069 119085 95103 119113
rect 95131 119085 100419 119113
rect 100447 119085 100481 119113
rect 100509 119085 110277 119113
rect 110305 119085 110339 119113
rect 110367 119085 110401 119113
rect 110429 119085 110463 119113
rect 110491 119085 115779 119113
rect 115807 119085 115841 119113
rect 115869 119085 125637 119113
rect 125665 119085 125699 119113
rect 125727 119085 125761 119113
rect 125789 119085 125823 119113
rect 125851 119085 131139 119113
rect 131167 119085 131201 119113
rect 131229 119085 140997 119113
rect 141025 119085 141059 119113
rect 141087 119085 141121 119113
rect 141149 119085 141183 119113
rect 141211 119085 146499 119113
rect 146527 119085 146561 119113
rect 146589 119085 156357 119113
rect 156385 119085 156419 119113
rect 156447 119085 156481 119113
rect 156509 119085 156543 119113
rect 156571 119085 161859 119113
rect 161887 119085 161921 119113
rect 161949 119085 171717 119113
rect 171745 119085 171779 119113
rect 171807 119085 171841 119113
rect 171869 119085 171903 119113
rect 171931 119085 177219 119113
rect 177247 119085 177281 119113
rect 177309 119085 187077 119113
rect 187105 119085 187139 119113
rect 187167 119085 187201 119113
rect 187229 119085 187263 119113
rect 187291 119085 192579 119113
rect 192607 119085 192641 119113
rect 192669 119085 202437 119113
rect 202465 119085 202499 119113
rect 202527 119085 202561 119113
rect 202589 119085 202623 119113
rect 202651 119085 207939 119113
rect 207967 119085 208001 119113
rect 208029 119085 217797 119113
rect 217825 119085 217859 119113
rect 217887 119085 217921 119113
rect 217949 119085 217983 119113
rect 218011 119085 223299 119113
rect 223327 119085 223361 119113
rect 223389 119085 233157 119113
rect 233185 119085 233219 119113
rect 233247 119085 233281 119113
rect 233309 119085 233343 119113
rect 233371 119085 238659 119113
rect 238687 119085 238721 119113
rect 238749 119085 248517 119113
rect 248545 119085 248579 119113
rect 248607 119085 248641 119113
rect 248669 119085 248703 119113
rect 248731 119085 254019 119113
rect 254047 119085 254081 119113
rect 254109 119085 263877 119113
rect 263905 119085 263939 119113
rect 263967 119085 264001 119113
rect 264029 119085 264063 119113
rect 264091 119085 269379 119113
rect 269407 119085 269441 119113
rect 269469 119085 279237 119113
rect 279265 119085 279299 119113
rect 279327 119085 279361 119113
rect 279389 119085 279423 119113
rect 279451 119085 284739 119113
rect 284767 119085 284801 119113
rect 284829 119085 294597 119113
rect 294625 119085 294659 119113
rect 294687 119085 294721 119113
rect 294749 119085 294783 119113
rect 294811 119085 298248 119113
rect 298276 119085 298310 119113
rect 298338 119085 298372 119113
rect 298400 119085 298434 119113
rect 298462 119085 298990 119113
rect -958 119051 298990 119085
rect -958 119023 -430 119051
rect -402 119023 -368 119051
rect -340 119023 -306 119051
rect -278 119023 -244 119051
rect -216 119023 2757 119051
rect 2785 119023 2819 119051
rect 2847 119023 2881 119051
rect 2909 119023 2943 119051
rect 2971 119023 8259 119051
rect 8287 119023 8321 119051
rect 8349 119023 18117 119051
rect 18145 119023 18179 119051
rect 18207 119023 18241 119051
rect 18269 119023 18303 119051
rect 18331 119023 23619 119051
rect 23647 119023 23681 119051
rect 23709 119023 33477 119051
rect 33505 119023 33539 119051
rect 33567 119023 33601 119051
rect 33629 119023 33663 119051
rect 33691 119023 38979 119051
rect 39007 119023 39041 119051
rect 39069 119023 48837 119051
rect 48865 119023 48899 119051
rect 48927 119023 48961 119051
rect 48989 119023 49023 119051
rect 49051 119023 54339 119051
rect 54367 119023 54401 119051
rect 54429 119023 64197 119051
rect 64225 119023 64259 119051
rect 64287 119023 64321 119051
rect 64349 119023 64383 119051
rect 64411 119023 69699 119051
rect 69727 119023 69761 119051
rect 69789 119023 79557 119051
rect 79585 119023 79619 119051
rect 79647 119023 79681 119051
rect 79709 119023 79743 119051
rect 79771 119023 85059 119051
rect 85087 119023 85121 119051
rect 85149 119023 94917 119051
rect 94945 119023 94979 119051
rect 95007 119023 95041 119051
rect 95069 119023 95103 119051
rect 95131 119023 100419 119051
rect 100447 119023 100481 119051
rect 100509 119023 110277 119051
rect 110305 119023 110339 119051
rect 110367 119023 110401 119051
rect 110429 119023 110463 119051
rect 110491 119023 115779 119051
rect 115807 119023 115841 119051
rect 115869 119023 125637 119051
rect 125665 119023 125699 119051
rect 125727 119023 125761 119051
rect 125789 119023 125823 119051
rect 125851 119023 131139 119051
rect 131167 119023 131201 119051
rect 131229 119023 140997 119051
rect 141025 119023 141059 119051
rect 141087 119023 141121 119051
rect 141149 119023 141183 119051
rect 141211 119023 146499 119051
rect 146527 119023 146561 119051
rect 146589 119023 156357 119051
rect 156385 119023 156419 119051
rect 156447 119023 156481 119051
rect 156509 119023 156543 119051
rect 156571 119023 161859 119051
rect 161887 119023 161921 119051
rect 161949 119023 171717 119051
rect 171745 119023 171779 119051
rect 171807 119023 171841 119051
rect 171869 119023 171903 119051
rect 171931 119023 177219 119051
rect 177247 119023 177281 119051
rect 177309 119023 187077 119051
rect 187105 119023 187139 119051
rect 187167 119023 187201 119051
rect 187229 119023 187263 119051
rect 187291 119023 192579 119051
rect 192607 119023 192641 119051
rect 192669 119023 202437 119051
rect 202465 119023 202499 119051
rect 202527 119023 202561 119051
rect 202589 119023 202623 119051
rect 202651 119023 207939 119051
rect 207967 119023 208001 119051
rect 208029 119023 217797 119051
rect 217825 119023 217859 119051
rect 217887 119023 217921 119051
rect 217949 119023 217983 119051
rect 218011 119023 223299 119051
rect 223327 119023 223361 119051
rect 223389 119023 233157 119051
rect 233185 119023 233219 119051
rect 233247 119023 233281 119051
rect 233309 119023 233343 119051
rect 233371 119023 238659 119051
rect 238687 119023 238721 119051
rect 238749 119023 248517 119051
rect 248545 119023 248579 119051
rect 248607 119023 248641 119051
rect 248669 119023 248703 119051
rect 248731 119023 254019 119051
rect 254047 119023 254081 119051
rect 254109 119023 263877 119051
rect 263905 119023 263939 119051
rect 263967 119023 264001 119051
rect 264029 119023 264063 119051
rect 264091 119023 269379 119051
rect 269407 119023 269441 119051
rect 269469 119023 279237 119051
rect 279265 119023 279299 119051
rect 279327 119023 279361 119051
rect 279389 119023 279423 119051
rect 279451 119023 284739 119051
rect 284767 119023 284801 119051
rect 284829 119023 294597 119051
rect 294625 119023 294659 119051
rect 294687 119023 294721 119051
rect 294749 119023 294783 119051
rect 294811 119023 298248 119051
rect 298276 119023 298310 119051
rect 298338 119023 298372 119051
rect 298400 119023 298434 119051
rect 298462 119023 298990 119051
rect -958 118989 298990 119023
rect -958 118961 -430 118989
rect -402 118961 -368 118989
rect -340 118961 -306 118989
rect -278 118961 -244 118989
rect -216 118961 2757 118989
rect 2785 118961 2819 118989
rect 2847 118961 2881 118989
rect 2909 118961 2943 118989
rect 2971 118961 8259 118989
rect 8287 118961 8321 118989
rect 8349 118961 18117 118989
rect 18145 118961 18179 118989
rect 18207 118961 18241 118989
rect 18269 118961 18303 118989
rect 18331 118961 23619 118989
rect 23647 118961 23681 118989
rect 23709 118961 33477 118989
rect 33505 118961 33539 118989
rect 33567 118961 33601 118989
rect 33629 118961 33663 118989
rect 33691 118961 38979 118989
rect 39007 118961 39041 118989
rect 39069 118961 48837 118989
rect 48865 118961 48899 118989
rect 48927 118961 48961 118989
rect 48989 118961 49023 118989
rect 49051 118961 54339 118989
rect 54367 118961 54401 118989
rect 54429 118961 64197 118989
rect 64225 118961 64259 118989
rect 64287 118961 64321 118989
rect 64349 118961 64383 118989
rect 64411 118961 69699 118989
rect 69727 118961 69761 118989
rect 69789 118961 79557 118989
rect 79585 118961 79619 118989
rect 79647 118961 79681 118989
rect 79709 118961 79743 118989
rect 79771 118961 85059 118989
rect 85087 118961 85121 118989
rect 85149 118961 94917 118989
rect 94945 118961 94979 118989
rect 95007 118961 95041 118989
rect 95069 118961 95103 118989
rect 95131 118961 100419 118989
rect 100447 118961 100481 118989
rect 100509 118961 110277 118989
rect 110305 118961 110339 118989
rect 110367 118961 110401 118989
rect 110429 118961 110463 118989
rect 110491 118961 115779 118989
rect 115807 118961 115841 118989
rect 115869 118961 125637 118989
rect 125665 118961 125699 118989
rect 125727 118961 125761 118989
rect 125789 118961 125823 118989
rect 125851 118961 131139 118989
rect 131167 118961 131201 118989
rect 131229 118961 140997 118989
rect 141025 118961 141059 118989
rect 141087 118961 141121 118989
rect 141149 118961 141183 118989
rect 141211 118961 146499 118989
rect 146527 118961 146561 118989
rect 146589 118961 156357 118989
rect 156385 118961 156419 118989
rect 156447 118961 156481 118989
rect 156509 118961 156543 118989
rect 156571 118961 161859 118989
rect 161887 118961 161921 118989
rect 161949 118961 171717 118989
rect 171745 118961 171779 118989
rect 171807 118961 171841 118989
rect 171869 118961 171903 118989
rect 171931 118961 177219 118989
rect 177247 118961 177281 118989
rect 177309 118961 187077 118989
rect 187105 118961 187139 118989
rect 187167 118961 187201 118989
rect 187229 118961 187263 118989
rect 187291 118961 192579 118989
rect 192607 118961 192641 118989
rect 192669 118961 202437 118989
rect 202465 118961 202499 118989
rect 202527 118961 202561 118989
rect 202589 118961 202623 118989
rect 202651 118961 207939 118989
rect 207967 118961 208001 118989
rect 208029 118961 217797 118989
rect 217825 118961 217859 118989
rect 217887 118961 217921 118989
rect 217949 118961 217983 118989
rect 218011 118961 223299 118989
rect 223327 118961 223361 118989
rect 223389 118961 233157 118989
rect 233185 118961 233219 118989
rect 233247 118961 233281 118989
rect 233309 118961 233343 118989
rect 233371 118961 238659 118989
rect 238687 118961 238721 118989
rect 238749 118961 248517 118989
rect 248545 118961 248579 118989
rect 248607 118961 248641 118989
rect 248669 118961 248703 118989
rect 248731 118961 254019 118989
rect 254047 118961 254081 118989
rect 254109 118961 263877 118989
rect 263905 118961 263939 118989
rect 263967 118961 264001 118989
rect 264029 118961 264063 118989
rect 264091 118961 269379 118989
rect 269407 118961 269441 118989
rect 269469 118961 279237 118989
rect 279265 118961 279299 118989
rect 279327 118961 279361 118989
rect 279389 118961 279423 118989
rect 279451 118961 284739 118989
rect 284767 118961 284801 118989
rect 284829 118961 294597 118989
rect 294625 118961 294659 118989
rect 294687 118961 294721 118989
rect 294749 118961 294783 118989
rect 294811 118961 298248 118989
rect 298276 118961 298310 118989
rect 298338 118961 298372 118989
rect 298400 118961 298434 118989
rect 298462 118961 298990 118989
rect -958 118913 298990 118961
rect -958 113175 298990 113223
rect -958 113147 -910 113175
rect -882 113147 -848 113175
rect -820 113147 -786 113175
rect -758 113147 -724 113175
rect -696 113147 4617 113175
rect 4645 113147 4679 113175
rect 4707 113147 4741 113175
rect 4769 113147 4803 113175
rect 4831 113147 15939 113175
rect 15967 113147 16001 113175
rect 16029 113147 19977 113175
rect 20005 113147 20039 113175
rect 20067 113147 20101 113175
rect 20129 113147 20163 113175
rect 20191 113147 31299 113175
rect 31327 113147 31361 113175
rect 31389 113147 35337 113175
rect 35365 113147 35399 113175
rect 35427 113147 35461 113175
rect 35489 113147 35523 113175
rect 35551 113147 46659 113175
rect 46687 113147 46721 113175
rect 46749 113147 50697 113175
rect 50725 113147 50759 113175
rect 50787 113147 50821 113175
rect 50849 113147 50883 113175
rect 50911 113147 62019 113175
rect 62047 113147 62081 113175
rect 62109 113147 66057 113175
rect 66085 113147 66119 113175
rect 66147 113147 66181 113175
rect 66209 113147 66243 113175
rect 66271 113147 77379 113175
rect 77407 113147 77441 113175
rect 77469 113147 81417 113175
rect 81445 113147 81479 113175
rect 81507 113147 81541 113175
rect 81569 113147 81603 113175
rect 81631 113147 92739 113175
rect 92767 113147 92801 113175
rect 92829 113147 96777 113175
rect 96805 113147 96839 113175
rect 96867 113147 96901 113175
rect 96929 113147 96963 113175
rect 96991 113147 108099 113175
rect 108127 113147 108161 113175
rect 108189 113147 112137 113175
rect 112165 113147 112199 113175
rect 112227 113147 112261 113175
rect 112289 113147 112323 113175
rect 112351 113147 123459 113175
rect 123487 113147 123521 113175
rect 123549 113147 127497 113175
rect 127525 113147 127559 113175
rect 127587 113147 127621 113175
rect 127649 113147 127683 113175
rect 127711 113147 138819 113175
rect 138847 113147 138881 113175
rect 138909 113147 142857 113175
rect 142885 113147 142919 113175
rect 142947 113147 142981 113175
rect 143009 113147 143043 113175
rect 143071 113147 154179 113175
rect 154207 113147 154241 113175
rect 154269 113147 158217 113175
rect 158245 113147 158279 113175
rect 158307 113147 158341 113175
rect 158369 113147 158403 113175
rect 158431 113147 169539 113175
rect 169567 113147 169601 113175
rect 169629 113147 173577 113175
rect 173605 113147 173639 113175
rect 173667 113147 173701 113175
rect 173729 113147 173763 113175
rect 173791 113147 184899 113175
rect 184927 113147 184961 113175
rect 184989 113147 188937 113175
rect 188965 113147 188999 113175
rect 189027 113147 189061 113175
rect 189089 113147 189123 113175
rect 189151 113147 200259 113175
rect 200287 113147 200321 113175
rect 200349 113147 204297 113175
rect 204325 113147 204359 113175
rect 204387 113147 204421 113175
rect 204449 113147 204483 113175
rect 204511 113147 215619 113175
rect 215647 113147 215681 113175
rect 215709 113147 219657 113175
rect 219685 113147 219719 113175
rect 219747 113147 219781 113175
rect 219809 113147 219843 113175
rect 219871 113147 230979 113175
rect 231007 113147 231041 113175
rect 231069 113147 235017 113175
rect 235045 113147 235079 113175
rect 235107 113147 235141 113175
rect 235169 113147 235203 113175
rect 235231 113147 246339 113175
rect 246367 113147 246401 113175
rect 246429 113147 250377 113175
rect 250405 113147 250439 113175
rect 250467 113147 250501 113175
rect 250529 113147 250563 113175
rect 250591 113147 261699 113175
rect 261727 113147 261761 113175
rect 261789 113147 265737 113175
rect 265765 113147 265799 113175
rect 265827 113147 265861 113175
rect 265889 113147 265923 113175
rect 265951 113147 277059 113175
rect 277087 113147 277121 113175
rect 277149 113147 281097 113175
rect 281125 113147 281159 113175
rect 281187 113147 281221 113175
rect 281249 113147 281283 113175
rect 281311 113147 296457 113175
rect 296485 113147 296519 113175
rect 296547 113147 296581 113175
rect 296609 113147 296643 113175
rect 296671 113147 298728 113175
rect 298756 113147 298790 113175
rect 298818 113147 298852 113175
rect 298880 113147 298914 113175
rect 298942 113147 298990 113175
rect -958 113113 298990 113147
rect -958 113085 -910 113113
rect -882 113085 -848 113113
rect -820 113085 -786 113113
rect -758 113085 -724 113113
rect -696 113085 4617 113113
rect 4645 113085 4679 113113
rect 4707 113085 4741 113113
rect 4769 113085 4803 113113
rect 4831 113085 15939 113113
rect 15967 113085 16001 113113
rect 16029 113085 19977 113113
rect 20005 113085 20039 113113
rect 20067 113085 20101 113113
rect 20129 113085 20163 113113
rect 20191 113085 31299 113113
rect 31327 113085 31361 113113
rect 31389 113085 35337 113113
rect 35365 113085 35399 113113
rect 35427 113085 35461 113113
rect 35489 113085 35523 113113
rect 35551 113085 46659 113113
rect 46687 113085 46721 113113
rect 46749 113085 50697 113113
rect 50725 113085 50759 113113
rect 50787 113085 50821 113113
rect 50849 113085 50883 113113
rect 50911 113085 62019 113113
rect 62047 113085 62081 113113
rect 62109 113085 66057 113113
rect 66085 113085 66119 113113
rect 66147 113085 66181 113113
rect 66209 113085 66243 113113
rect 66271 113085 77379 113113
rect 77407 113085 77441 113113
rect 77469 113085 81417 113113
rect 81445 113085 81479 113113
rect 81507 113085 81541 113113
rect 81569 113085 81603 113113
rect 81631 113085 92739 113113
rect 92767 113085 92801 113113
rect 92829 113085 96777 113113
rect 96805 113085 96839 113113
rect 96867 113085 96901 113113
rect 96929 113085 96963 113113
rect 96991 113085 108099 113113
rect 108127 113085 108161 113113
rect 108189 113085 112137 113113
rect 112165 113085 112199 113113
rect 112227 113085 112261 113113
rect 112289 113085 112323 113113
rect 112351 113085 123459 113113
rect 123487 113085 123521 113113
rect 123549 113085 127497 113113
rect 127525 113085 127559 113113
rect 127587 113085 127621 113113
rect 127649 113085 127683 113113
rect 127711 113085 138819 113113
rect 138847 113085 138881 113113
rect 138909 113085 142857 113113
rect 142885 113085 142919 113113
rect 142947 113085 142981 113113
rect 143009 113085 143043 113113
rect 143071 113085 154179 113113
rect 154207 113085 154241 113113
rect 154269 113085 158217 113113
rect 158245 113085 158279 113113
rect 158307 113085 158341 113113
rect 158369 113085 158403 113113
rect 158431 113085 169539 113113
rect 169567 113085 169601 113113
rect 169629 113085 173577 113113
rect 173605 113085 173639 113113
rect 173667 113085 173701 113113
rect 173729 113085 173763 113113
rect 173791 113085 184899 113113
rect 184927 113085 184961 113113
rect 184989 113085 188937 113113
rect 188965 113085 188999 113113
rect 189027 113085 189061 113113
rect 189089 113085 189123 113113
rect 189151 113085 200259 113113
rect 200287 113085 200321 113113
rect 200349 113085 204297 113113
rect 204325 113085 204359 113113
rect 204387 113085 204421 113113
rect 204449 113085 204483 113113
rect 204511 113085 215619 113113
rect 215647 113085 215681 113113
rect 215709 113085 219657 113113
rect 219685 113085 219719 113113
rect 219747 113085 219781 113113
rect 219809 113085 219843 113113
rect 219871 113085 230979 113113
rect 231007 113085 231041 113113
rect 231069 113085 235017 113113
rect 235045 113085 235079 113113
rect 235107 113085 235141 113113
rect 235169 113085 235203 113113
rect 235231 113085 246339 113113
rect 246367 113085 246401 113113
rect 246429 113085 250377 113113
rect 250405 113085 250439 113113
rect 250467 113085 250501 113113
rect 250529 113085 250563 113113
rect 250591 113085 261699 113113
rect 261727 113085 261761 113113
rect 261789 113085 265737 113113
rect 265765 113085 265799 113113
rect 265827 113085 265861 113113
rect 265889 113085 265923 113113
rect 265951 113085 277059 113113
rect 277087 113085 277121 113113
rect 277149 113085 281097 113113
rect 281125 113085 281159 113113
rect 281187 113085 281221 113113
rect 281249 113085 281283 113113
rect 281311 113085 296457 113113
rect 296485 113085 296519 113113
rect 296547 113085 296581 113113
rect 296609 113085 296643 113113
rect 296671 113085 298728 113113
rect 298756 113085 298790 113113
rect 298818 113085 298852 113113
rect 298880 113085 298914 113113
rect 298942 113085 298990 113113
rect -958 113051 298990 113085
rect -958 113023 -910 113051
rect -882 113023 -848 113051
rect -820 113023 -786 113051
rect -758 113023 -724 113051
rect -696 113023 4617 113051
rect 4645 113023 4679 113051
rect 4707 113023 4741 113051
rect 4769 113023 4803 113051
rect 4831 113023 15939 113051
rect 15967 113023 16001 113051
rect 16029 113023 19977 113051
rect 20005 113023 20039 113051
rect 20067 113023 20101 113051
rect 20129 113023 20163 113051
rect 20191 113023 31299 113051
rect 31327 113023 31361 113051
rect 31389 113023 35337 113051
rect 35365 113023 35399 113051
rect 35427 113023 35461 113051
rect 35489 113023 35523 113051
rect 35551 113023 46659 113051
rect 46687 113023 46721 113051
rect 46749 113023 50697 113051
rect 50725 113023 50759 113051
rect 50787 113023 50821 113051
rect 50849 113023 50883 113051
rect 50911 113023 62019 113051
rect 62047 113023 62081 113051
rect 62109 113023 66057 113051
rect 66085 113023 66119 113051
rect 66147 113023 66181 113051
rect 66209 113023 66243 113051
rect 66271 113023 77379 113051
rect 77407 113023 77441 113051
rect 77469 113023 81417 113051
rect 81445 113023 81479 113051
rect 81507 113023 81541 113051
rect 81569 113023 81603 113051
rect 81631 113023 92739 113051
rect 92767 113023 92801 113051
rect 92829 113023 96777 113051
rect 96805 113023 96839 113051
rect 96867 113023 96901 113051
rect 96929 113023 96963 113051
rect 96991 113023 108099 113051
rect 108127 113023 108161 113051
rect 108189 113023 112137 113051
rect 112165 113023 112199 113051
rect 112227 113023 112261 113051
rect 112289 113023 112323 113051
rect 112351 113023 123459 113051
rect 123487 113023 123521 113051
rect 123549 113023 127497 113051
rect 127525 113023 127559 113051
rect 127587 113023 127621 113051
rect 127649 113023 127683 113051
rect 127711 113023 138819 113051
rect 138847 113023 138881 113051
rect 138909 113023 142857 113051
rect 142885 113023 142919 113051
rect 142947 113023 142981 113051
rect 143009 113023 143043 113051
rect 143071 113023 154179 113051
rect 154207 113023 154241 113051
rect 154269 113023 158217 113051
rect 158245 113023 158279 113051
rect 158307 113023 158341 113051
rect 158369 113023 158403 113051
rect 158431 113023 169539 113051
rect 169567 113023 169601 113051
rect 169629 113023 173577 113051
rect 173605 113023 173639 113051
rect 173667 113023 173701 113051
rect 173729 113023 173763 113051
rect 173791 113023 184899 113051
rect 184927 113023 184961 113051
rect 184989 113023 188937 113051
rect 188965 113023 188999 113051
rect 189027 113023 189061 113051
rect 189089 113023 189123 113051
rect 189151 113023 200259 113051
rect 200287 113023 200321 113051
rect 200349 113023 204297 113051
rect 204325 113023 204359 113051
rect 204387 113023 204421 113051
rect 204449 113023 204483 113051
rect 204511 113023 215619 113051
rect 215647 113023 215681 113051
rect 215709 113023 219657 113051
rect 219685 113023 219719 113051
rect 219747 113023 219781 113051
rect 219809 113023 219843 113051
rect 219871 113023 230979 113051
rect 231007 113023 231041 113051
rect 231069 113023 235017 113051
rect 235045 113023 235079 113051
rect 235107 113023 235141 113051
rect 235169 113023 235203 113051
rect 235231 113023 246339 113051
rect 246367 113023 246401 113051
rect 246429 113023 250377 113051
rect 250405 113023 250439 113051
rect 250467 113023 250501 113051
rect 250529 113023 250563 113051
rect 250591 113023 261699 113051
rect 261727 113023 261761 113051
rect 261789 113023 265737 113051
rect 265765 113023 265799 113051
rect 265827 113023 265861 113051
rect 265889 113023 265923 113051
rect 265951 113023 277059 113051
rect 277087 113023 277121 113051
rect 277149 113023 281097 113051
rect 281125 113023 281159 113051
rect 281187 113023 281221 113051
rect 281249 113023 281283 113051
rect 281311 113023 296457 113051
rect 296485 113023 296519 113051
rect 296547 113023 296581 113051
rect 296609 113023 296643 113051
rect 296671 113023 298728 113051
rect 298756 113023 298790 113051
rect 298818 113023 298852 113051
rect 298880 113023 298914 113051
rect 298942 113023 298990 113051
rect -958 112989 298990 113023
rect -958 112961 -910 112989
rect -882 112961 -848 112989
rect -820 112961 -786 112989
rect -758 112961 -724 112989
rect -696 112961 4617 112989
rect 4645 112961 4679 112989
rect 4707 112961 4741 112989
rect 4769 112961 4803 112989
rect 4831 112961 15939 112989
rect 15967 112961 16001 112989
rect 16029 112961 19977 112989
rect 20005 112961 20039 112989
rect 20067 112961 20101 112989
rect 20129 112961 20163 112989
rect 20191 112961 31299 112989
rect 31327 112961 31361 112989
rect 31389 112961 35337 112989
rect 35365 112961 35399 112989
rect 35427 112961 35461 112989
rect 35489 112961 35523 112989
rect 35551 112961 46659 112989
rect 46687 112961 46721 112989
rect 46749 112961 50697 112989
rect 50725 112961 50759 112989
rect 50787 112961 50821 112989
rect 50849 112961 50883 112989
rect 50911 112961 62019 112989
rect 62047 112961 62081 112989
rect 62109 112961 66057 112989
rect 66085 112961 66119 112989
rect 66147 112961 66181 112989
rect 66209 112961 66243 112989
rect 66271 112961 77379 112989
rect 77407 112961 77441 112989
rect 77469 112961 81417 112989
rect 81445 112961 81479 112989
rect 81507 112961 81541 112989
rect 81569 112961 81603 112989
rect 81631 112961 92739 112989
rect 92767 112961 92801 112989
rect 92829 112961 96777 112989
rect 96805 112961 96839 112989
rect 96867 112961 96901 112989
rect 96929 112961 96963 112989
rect 96991 112961 108099 112989
rect 108127 112961 108161 112989
rect 108189 112961 112137 112989
rect 112165 112961 112199 112989
rect 112227 112961 112261 112989
rect 112289 112961 112323 112989
rect 112351 112961 123459 112989
rect 123487 112961 123521 112989
rect 123549 112961 127497 112989
rect 127525 112961 127559 112989
rect 127587 112961 127621 112989
rect 127649 112961 127683 112989
rect 127711 112961 138819 112989
rect 138847 112961 138881 112989
rect 138909 112961 142857 112989
rect 142885 112961 142919 112989
rect 142947 112961 142981 112989
rect 143009 112961 143043 112989
rect 143071 112961 154179 112989
rect 154207 112961 154241 112989
rect 154269 112961 158217 112989
rect 158245 112961 158279 112989
rect 158307 112961 158341 112989
rect 158369 112961 158403 112989
rect 158431 112961 169539 112989
rect 169567 112961 169601 112989
rect 169629 112961 173577 112989
rect 173605 112961 173639 112989
rect 173667 112961 173701 112989
rect 173729 112961 173763 112989
rect 173791 112961 184899 112989
rect 184927 112961 184961 112989
rect 184989 112961 188937 112989
rect 188965 112961 188999 112989
rect 189027 112961 189061 112989
rect 189089 112961 189123 112989
rect 189151 112961 200259 112989
rect 200287 112961 200321 112989
rect 200349 112961 204297 112989
rect 204325 112961 204359 112989
rect 204387 112961 204421 112989
rect 204449 112961 204483 112989
rect 204511 112961 215619 112989
rect 215647 112961 215681 112989
rect 215709 112961 219657 112989
rect 219685 112961 219719 112989
rect 219747 112961 219781 112989
rect 219809 112961 219843 112989
rect 219871 112961 230979 112989
rect 231007 112961 231041 112989
rect 231069 112961 235017 112989
rect 235045 112961 235079 112989
rect 235107 112961 235141 112989
rect 235169 112961 235203 112989
rect 235231 112961 246339 112989
rect 246367 112961 246401 112989
rect 246429 112961 250377 112989
rect 250405 112961 250439 112989
rect 250467 112961 250501 112989
rect 250529 112961 250563 112989
rect 250591 112961 261699 112989
rect 261727 112961 261761 112989
rect 261789 112961 265737 112989
rect 265765 112961 265799 112989
rect 265827 112961 265861 112989
rect 265889 112961 265923 112989
rect 265951 112961 277059 112989
rect 277087 112961 277121 112989
rect 277149 112961 281097 112989
rect 281125 112961 281159 112989
rect 281187 112961 281221 112989
rect 281249 112961 281283 112989
rect 281311 112961 296457 112989
rect 296485 112961 296519 112989
rect 296547 112961 296581 112989
rect 296609 112961 296643 112989
rect 296671 112961 298728 112989
rect 298756 112961 298790 112989
rect 298818 112961 298852 112989
rect 298880 112961 298914 112989
rect 298942 112961 298990 112989
rect -958 112913 298990 112961
rect -958 110175 298990 110223
rect -958 110147 -430 110175
rect -402 110147 -368 110175
rect -340 110147 -306 110175
rect -278 110147 -244 110175
rect -216 110147 2757 110175
rect 2785 110147 2819 110175
rect 2847 110147 2881 110175
rect 2909 110147 2943 110175
rect 2971 110147 8259 110175
rect 8287 110147 8321 110175
rect 8349 110147 18117 110175
rect 18145 110147 18179 110175
rect 18207 110147 18241 110175
rect 18269 110147 18303 110175
rect 18331 110147 23619 110175
rect 23647 110147 23681 110175
rect 23709 110147 33477 110175
rect 33505 110147 33539 110175
rect 33567 110147 33601 110175
rect 33629 110147 33663 110175
rect 33691 110147 38979 110175
rect 39007 110147 39041 110175
rect 39069 110147 48837 110175
rect 48865 110147 48899 110175
rect 48927 110147 48961 110175
rect 48989 110147 49023 110175
rect 49051 110147 54339 110175
rect 54367 110147 54401 110175
rect 54429 110147 64197 110175
rect 64225 110147 64259 110175
rect 64287 110147 64321 110175
rect 64349 110147 64383 110175
rect 64411 110147 69699 110175
rect 69727 110147 69761 110175
rect 69789 110147 79557 110175
rect 79585 110147 79619 110175
rect 79647 110147 79681 110175
rect 79709 110147 79743 110175
rect 79771 110147 85059 110175
rect 85087 110147 85121 110175
rect 85149 110147 94917 110175
rect 94945 110147 94979 110175
rect 95007 110147 95041 110175
rect 95069 110147 95103 110175
rect 95131 110147 100419 110175
rect 100447 110147 100481 110175
rect 100509 110147 110277 110175
rect 110305 110147 110339 110175
rect 110367 110147 110401 110175
rect 110429 110147 110463 110175
rect 110491 110147 115779 110175
rect 115807 110147 115841 110175
rect 115869 110147 125637 110175
rect 125665 110147 125699 110175
rect 125727 110147 125761 110175
rect 125789 110147 125823 110175
rect 125851 110147 131139 110175
rect 131167 110147 131201 110175
rect 131229 110147 140997 110175
rect 141025 110147 141059 110175
rect 141087 110147 141121 110175
rect 141149 110147 141183 110175
rect 141211 110147 146499 110175
rect 146527 110147 146561 110175
rect 146589 110147 156357 110175
rect 156385 110147 156419 110175
rect 156447 110147 156481 110175
rect 156509 110147 156543 110175
rect 156571 110147 161859 110175
rect 161887 110147 161921 110175
rect 161949 110147 171717 110175
rect 171745 110147 171779 110175
rect 171807 110147 171841 110175
rect 171869 110147 171903 110175
rect 171931 110147 177219 110175
rect 177247 110147 177281 110175
rect 177309 110147 187077 110175
rect 187105 110147 187139 110175
rect 187167 110147 187201 110175
rect 187229 110147 187263 110175
rect 187291 110147 192579 110175
rect 192607 110147 192641 110175
rect 192669 110147 202437 110175
rect 202465 110147 202499 110175
rect 202527 110147 202561 110175
rect 202589 110147 202623 110175
rect 202651 110147 207939 110175
rect 207967 110147 208001 110175
rect 208029 110147 217797 110175
rect 217825 110147 217859 110175
rect 217887 110147 217921 110175
rect 217949 110147 217983 110175
rect 218011 110147 223299 110175
rect 223327 110147 223361 110175
rect 223389 110147 233157 110175
rect 233185 110147 233219 110175
rect 233247 110147 233281 110175
rect 233309 110147 233343 110175
rect 233371 110147 238659 110175
rect 238687 110147 238721 110175
rect 238749 110147 248517 110175
rect 248545 110147 248579 110175
rect 248607 110147 248641 110175
rect 248669 110147 248703 110175
rect 248731 110147 254019 110175
rect 254047 110147 254081 110175
rect 254109 110147 263877 110175
rect 263905 110147 263939 110175
rect 263967 110147 264001 110175
rect 264029 110147 264063 110175
rect 264091 110147 269379 110175
rect 269407 110147 269441 110175
rect 269469 110147 279237 110175
rect 279265 110147 279299 110175
rect 279327 110147 279361 110175
rect 279389 110147 279423 110175
rect 279451 110147 284739 110175
rect 284767 110147 284801 110175
rect 284829 110147 294597 110175
rect 294625 110147 294659 110175
rect 294687 110147 294721 110175
rect 294749 110147 294783 110175
rect 294811 110147 298248 110175
rect 298276 110147 298310 110175
rect 298338 110147 298372 110175
rect 298400 110147 298434 110175
rect 298462 110147 298990 110175
rect -958 110113 298990 110147
rect -958 110085 -430 110113
rect -402 110085 -368 110113
rect -340 110085 -306 110113
rect -278 110085 -244 110113
rect -216 110085 2757 110113
rect 2785 110085 2819 110113
rect 2847 110085 2881 110113
rect 2909 110085 2943 110113
rect 2971 110085 8259 110113
rect 8287 110085 8321 110113
rect 8349 110085 18117 110113
rect 18145 110085 18179 110113
rect 18207 110085 18241 110113
rect 18269 110085 18303 110113
rect 18331 110085 23619 110113
rect 23647 110085 23681 110113
rect 23709 110085 33477 110113
rect 33505 110085 33539 110113
rect 33567 110085 33601 110113
rect 33629 110085 33663 110113
rect 33691 110085 38979 110113
rect 39007 110085 39041 110113
rect 39069 110085 48837 110113
rect 48865 110085 48899 110113
rect 48927 110085 48961 110113
rect 48989 110085 49023 110113
rect 49051 110085 54339 110113
rect 54367 110085 54401 110113
rect 54429 110085 64197 110113
rect 64225 110085 64259 110113
rect 64287 110085 64321 110113
rect 64349 110085 64383 110113
rect 64411 110085 69699 110113
rect 69727 110085 69761 110113
rect 69789 110085 79557 110113
rect 79585 110085 79619 110113
rect 79647 110085 79681 110113
rect 79709 110085 79743 110113
rect 79771 110085 85059 110113
rect 85087 110085 85121 110113
rect 85149 110085 94917 110113
rect 94945 110085 94979 110113
rect 95007 110085 95041 110113
rect 95069 110085 95103 110113
rect 95131 110085 100419 110113
rect 100447 110085 100481 110113
rect 100509 110085 110277 110113
rect 110305 110085 110339 110113
rect 110367 110085 110401 110113
rect 110429 110085 110463 110113
rect 110491 110085 115779 110113
rect 115807 110085 115841 110113
rect 115869 110085 125637 110113
rect 125665 110085 125699 110113
rect 125727 110085 125761 110113
rect 125789 110085 125823 110113
rect 125851 110085 131139 110113
rect 131167 110085 131201 110113
rect 131229 110085 140997 110113
rect 141025 110085 141059 110113
rect 141087 110085 141121 110113
rect 141149 110085 141183 110113
rect 141211 110085 146499 110113
rect 146527 110085 146561 110113
rect 146589 110085 156357 110113
rect 156385 110085 156419 110113
rect 156447 110085 156481 110113
rect 156509 110085 156543 110113
rect 156571 110085 161859 110113
rect 161887 110085 161921 110113
rect 161949 110085 171717 110113
rect 171745 110085 171779 110113
rect 171807 110085 171841 110113
rect 171869 110085 171903 110113
rect 171931 110085 177219 110113
rect 177247 110085 177281 110113
rect 177309 110085 187077 110113
rect 187105 110085 187139 110113
rect 187167 110085 187201 110113
rect 187229 110085 187263 110113
rect 187291 110085 192579 110113
rect 192607 110085 192641 110113
rect 192669 110085 202437 110113
rect 202465 110085 202499 110113
rect 202527 110085 202561 110113
rect 202589 110085 202623 110113
rect 202651 110085 207939 110113
rect 207967 110085 208001 110113
rect 208029 110085 217797 110113
rect 217825 110085 217859 110113
rect 217887 110085 217921 110113
rect 217949 110085 217983 110113
rect 218011 110085 223299 110113
rect 223327 110085 223361 110113
rect 223389 110085 233157 110113
rect 233185 110085 233219 110113
rect 233247 110085 233281 110113
rect 233309 110085 233343 110113
rect 233371 110085 238659 110113
rect 238687 110085 238721 110113
rect 238749 110085 248517 110113
rect 248545 110085 248579 110113
rect 248607 110085 248641 110113
rect 248669 110085 248703 110113
rect 248731 110085 254019 110113
rect 254047 110085 254081 110113
rect 254109 110085 263877 110113
rect 263905 110085 263939 110113
rect 263967 110085 264001 110113
rect 264029 110085 264063 110113
rect 264091 110085 269379 110113
rect 269407 110085 269441 110113
rect 269469 110085 279237 110113
rect 279265 110085 279299 110113
rect 279327 110085 279361 110113
rect 279389 110085 279423 110113
rect 279451 110085 284739 110113
rect 284767 110085 284801 110113
rect 284829 110085 294597 110113
rect 294625 110085 294659 110113
rect 294687 110085 294721 110113
rect 294749 110085 294783 110113
rect 294811 110085 298248 110113
rect 298276 110085 298310 110113
rect 298338 110085 298372 110113
rect 298400 110085 298434 110113
rect 298462 110085 298990 110113
rect -958 110051 298990 110085
rect -958 110023 -430 110051
rect -402 110023 -368 110051
rect -340 110023 -306 110051
rect -278 110023 -244 110051
rect -216 110023 2757 110051
rect 2785 110023 2819 110051
rect 2847 110023 2881 110051
rect 2909 110023 2943 110051
rect 2971 110023 8259 110051
rect 8287 110023 8321 110051
rect 8349 110023 18117 110051
rect 18145 110023 18179 110051
rect 18207 110023 18241 110051
rect 18269 110023 18303 110051
rect 18331 110023 23619 110051
rect 23647 110023 23681 110051
rect 23709 110023 33477 110051
rect 33505 110023 33539 110051
rect 33567 110023 33601 110051
rect 33629 110023 33663 110051
rect 33691 110023 38979 110051
rect 39007 110023 39041 110051
rect 39069 110023 48837 110051
rect 48865 110023 48899 110051
rect 48927 110023 48961 110051
rect 48989 110023 49023 110051
rect 49051 110023 54339 110051
rect 54367 110023 54401 110051
rect 54429 110023 64197 110051
rect 64225 110023 64259 110051
rect 64287 110023 64321 110051
rect 64349 110023 64383 110051
rect 64411 110023 69699 110051
rect 69727 110023 69761 110051
rect 69789 110023 79557 110051
rect 79585 110023 79619 110051
rect 79647 110023 79681 110051
rect 79709 110023 79743 110051
rect 79771 110023 85059 110051
rect 85087 110023 85121 110051
rect 85149 110023 94917 110051
rect 94945 110023 94979 110051
rect 95007 110023 95041 110051
rect 95069 110023 95103 110051
rect 95131 110023 100419 110051
rect 100447 110023 100481 110051
rect 100509 110023 110277 110051
rect 110305 110023 110339 110051
rect 110367 110023 110401 110051
rect 110429 110023 110463 110051
rect 110491 110023 115779 110051
rect 115807 110023 115841 110051
rect 115869 110023 125637 110051
rect 125665 110023 125699 110051
rect 125727 110023 125761 110051
rect 125789 110023 125823 110051
rect 125851 110023 131139 110051
rect 131167 110023 131201 110051
rect 131229 110023 140997 110051
rect 141025 110023 141059 110051
rect 141087 110023 141121 110051
rect 141149 110023 141183 110051
rect 141211 110023 146499 110051
rect 146527 110023 146561 110051
rect 146589 110023 156357 110051
rect 156385 110023 156419 110051
rect 156447 110023 156481 110051
rect 156509 110023 156543 110051
rect 156571 110023 161859 110051
rect 161887 110023 161921 110051
rect 161949 110023 171717 110051
rect 171745 110023 171779 110051
rect 171807 110023 171841 110051
rect 171869 110023 171903 110051
rect 171931 110023 177219 110051
rect 177247 110023 177281 110051
rect 177309 110023 187077 110051
rect 187105 110023 187139 110051
rect 187167 110023 187201 110051
rect 187229 110023 187263 110051
rect 187291 110023 192579 110051
rect 192607 110023 192641 110051
rect 192669 110023 202437 110051
rect 202465 110023 202499 110051
rect 202527 110023 202561 110051
rect 202589 110023 202623 110051
rect 202651 110023 207939 110051
rect 207967 110023 208001 110051
rect 208029 110023 217797 110051
rect 217825 110023 217859 110051
rect 217887 110023 217921 110051
rect 217949 110023 217983 110051
rect 218011 110023 223299 110051
rect 223327 110023 223361 110051
rect 223389 110023 233157 110051
rect 233185 110023 233219 110051
rect 233247 110023 233281 110051
rect 233309 110023 233343 110051
rect 233371 110023 238659 110051
rect 238687 110023 238721 110051
rect 238749 110023 248517 110051
rect 248545 110023 248579 110051
rect 248607 110023 248641 110051
rect 248669 110023 248703 110051
rect 248731 110023 254019 110051
rect 254047 110023 254081 110051
rect 254109 110023 263877 110051
rect 263905 110023 263939 110051
rect 263967 110023 264001 110051
rect 264029 110023 264063 110051
rect 264091 110023 269379 110051
rect 269407 110023 269441 110051
rect 269469 110023 279237 110051
rect 279265 110023 279299 110051
rect 279327 110023 279361 110051
rect 279389 110023 279423 110051
rect 279451 110023 284739 110051
rect 284767 110023 284801 110051
rect 284829 110023 294597 110051
rect 294625 110023 294659 110051
rect 294687 110023 294721 110051
rect 294749 110023 294783 110051
rect 294811 110023 298248 110051
rect 298276 110023 298310 110051
rect 298338 110023 298372 110051
rect 298400 110023 298434 110051
rect 298462 110023 298990 110051
rect -958 109989 298990 110023
rect -958 109961 -430 109989
rect -402 109961 -368 109989
rect -340 109961 -306 109989
rect -278 109961 -244 109989
rect -216 109961 2757 109989
rect 2785 109961 2819 109989
rect 2847 109961 2881 109989
rect 2909 109961 2943 109989
rect 2971 109961 8259 109989
rect 8287 109961 8321 109989
rect 8349 109961 18117 109989
rect 18145 109961 18179 109989
rect 18207 109961 18241 109989
rect 18269 109961 18303 109989
rect 18331 109961 23619 109989
rect 23647 109961 23681 109989
rect 23709 109961 33477 109989
rect 33505 109961 33539 109989
rect 33567 109961 33601 109989
rect 33629 109961 33663 109989
rect 33691 109961 38979 109989
rect 39007 109961 39041 109989
rect 39069 109961 48837 109989
rect 48865 109961 48899 109989
rect 48927 109961 48961 109989
rect 48989 109961 49023 109989
rect 49051 109961 54339 109989
rect 54367 109961 54401 109989
rect 54429 109961 64197 109989
rect 64225 109961 64259 109989
rect 64287 109961 64321 109989
rect 64349 109961 64383 109989
rect 64411 109961 69699 109989
rect 69727 109961 69761 109989
rect 69789 109961 79557 109989
rect 79585 109961 79619 109989
rect 79647 109961 79681 109989
rect 79709 109961 79743 109989
rect 79771 109961 85059 109989
rect 85087 109961 85121 109989
rect 85149 109961 94917 109989
rect 94945 109961 94979 109989
rect 95007 109961 95041 109989
rect 95069 109961 95103 109989
rect 95131 109961 100419 109989
rect 100447 109961 100481 109989
rect 100509 109961 110277 109989
rect 110305 109961 110339 109989
rect 110367 109961 110401 109989
rect 110429 109961 110463 109989
rect 110491 109961 115779 109989
rect 115807 109961 115841 109989
rect 115869 109961 125637 109989
rect 125665 109961 125699 109989
rect 125727 109961 125761 109989
rect 125789 109961 125823 109989
rect 125851 109961 131139 109989
rect 131167 109961 131201 109989
rect 131229 109961 140997 109989
rect 141025 109961 141059 109989
rect 141087 109961 141121 109989
rect 141149 109961 141183 109989
rect 141211 109961 146499 109989
rect 146527 109961 146561 109989
rect 146589 109961 156357 109989
rect 156385 109961 156419 109989
rect 156447 109961 156481 109989
rect 156509 109961 156543 109989
rect 156571 109961 161859 109989
rect 161887 109961 161921 109989
rect 161949 109961 171717 109989
rect 171745 109961 171779 109989
rect 171807 109961 171841 109989
rect 171869 109961 171903 109989
rect 171931 109961 177219 109989
rect 177247 109961 177281 109989
rect 177309 109961 187077 109989
rect 187105 109961 187139 109989
rect 187167 109961 187201 109989
rect 187229 109961 187263 109989
rect 187291 109961 192579 109989
rect 192607 109961 192641 109989
rect 192669 109961 202437 109989
rect 202465 109961 202499 109989
rect 202527 109961 202561 109989
rect 202589 109961 202623 109989
rect 202651 109961 207939 109989
rect 207967 109961 208001 109989
rect 208029 109961 217797 109989
rect 217825 109961 217859 109989
rect 217887 109961 217921 109989
rect 217949 109961 217983 109989
rect 218011 109961 223299 109989
rect 223327 109961 223361 109989
rect 223389 109961 233157 109989
rect 233185 109961 233219 109989
rect 233247 109961 233281 109989
rect 233309 109961 233343 109989
rect 233371 109961 238659 109989
rect 238687 109961 238721 109989
rect 238749 109961 248517 109989
rect 248545 109961 248579 109989
rect 248607 109961 248641 109989
rect 248669 109961 248703 109989
rect 248731 109961 254019 109989
rect 254047 109961 254081 109989
rect 254109 109961 263877 109989
rect 263905 109961 263939 109989
rect 263967 109961 264001 109989
rect 264029 109961 264063 109989
rect 264091 109961 269379 109989
rect 269407 109961 269441 109989
rect 269469 109961 279237 109989
rect 279265 109961 279299 109989
rect 279327 109961 279361 109989
rect 279389 109961 279423 109989
rect 279451 109961 284739 109989
rect 284767 109961 284801 109989
rect 284829 109961 294597 109989
rect 294625 109961 294659 109989
rect 294687 109961 294721 109989
rect 294749 109961 294783 109989
rect 294811 109961 298248 109989
rect 298276 109961 298310 109989
rect 298338 109961 298372 109989
rect 298400 109961 298434 109989
rect 298462 109961 298990 109989
rect -958 109913 298990 109961
rect -958 104175 298990 104223
rect -958 104147 -910 104175
rect -882 104147 -848 104175
rect -820 104147 -786 104175
rect -758 104147 -724 104175
rect -696 104147 4617 104175
rect 4645 104147 4679 104175
rect 4707 104147 4741 104175
rect 4769 104147 4803 104175
rect 4831 104147 15939 104175
rect 15967 104147 16001 104175
rect 16029 104147 19977 104175
rect 20005 104147 20039 104175
rect 20067 104147 20101 104175
rect 20129 104147 20163 104175
rect 20191 104147 31299 104175
rect 31327 104147 31361 104175
rect 31389 104147 35337 104175
rect 35365 104147 35399 104175
rect 35427 104147 35461 104175
rect 35489 104147 35523 104175
rect 35551 104147 46659 104175
rect 46687 104147 46721 104175
rect 46749 104147 50697 104175
rect 50725 104147 50759 104175
rect 50787 104147 50821 104175
rect 50849 104147 50883 104175
rect 50911 104147 62019 104175
rect 62047 104147 62081 104175
rect 62109 104147 66057 104175
rect 66085 104147 66119 104175
rect 66147 104147 66181 104175
rect 66209 104147 66243 104175
rect 66271 104147 77379 104175
rect 77407 104147 77441 104175
rect 77469 104147 81417 104175
rect 81445 104147 81479 104175
rect 81507 104147 81541 104175
rect 81569 104147 81603 104175
rect 81631 104147 92739 104175
rect 92767 104147 92801 104175
rect 92829 104147 96777 104175
rect 96805 104147 96839 104175
rect 96867 104147 96901 104175
rect 96929 104147 96963 104175
rect 96991 104147 108099 104175
rect 108127 104147 108161 104175
rect 108189 104147 112137 104175
rect 112165 104147 112199 104175
rect 112227 104147 112261 104175
rect 112289 104147 112323 104175
rect 112351 104147 123459 104175
rect 123487 104147 123521 104175
rect 123549 104147 127497 104175
rect 127525 104147 127559 104175
rect 127587 104147 127621 104175
rect 127649 104147 127683 104175
rect 127711 104147 138819 104175
rect 138847 104147 138881 104175
rect 138909 104147 142857 104175
rect 142885 104147 142919 104175
rect 142947 104147 142981 104175
rect 143009 104147 143043 104175
rect 143071 104147 154179 104175
rect 154207 104147 154241 104175
rect 154269 104147 158217 104175
rect 158245 104147 158279 104175
rect 158307 104147 158341 104175
rect 158369 104147 158403 104175
rect 158431 104147 169539 104175
rect 169567 104147 169601 104175
rect 169629 104147 173577 104175
rect 173605 104147 173639 104175
rect 173667 104147 173701 104175
rect 173729 104147 173763 104175
rect 173791 104147 184899 104175
rect 184927 104147 184961 104175
rect 184989 104147 188937 104175
rect 188965 104147 188999 104175
rect 189027 104147 189061 104175
rect 189089 104147 189123 104175
rect 189151 104147 200259 104175
rect 200287 104147 200321 104175
rect 200349 104147 204297 104175
rect 204325 104147 204359 104175
rect 204387 104147 204421 104175
rect 204449 104147 204483 104175
rect 204511 104147 215619 104175
rect 215647 104147 215681 104175
rect 215709 104147 219657 104175
rect 219685 104147 219719 104175
rect 219747 104147 219781 104175
rect 219809 104147 219843 104175
rect 219871 104147 230979 104175
rect 231007 104147 231041 104175
rect 231069 104147 235017 104175
rect 235045 104147 235079 104175
rect 235107 104147 235141 104175
rect 235169 104147 235203 104175
rect 235231 104147 246339 104175
rect 246367 104147 246401 104175
rect 246429 104147 250377 104175
rect 250405 104147 250439 104175
rect 250467 104147 250501 104175
rect 250529 104147 250563 104175
rect 250591 104147 261699 104175
rect 261727 104147 261761 104175
rect 261789 104147 265737 104175
rect 265765 104147 265799 104175
rect 265827 104147 265861 104175
rect 265889 104147 265923 104175
rect 265951 104147 277059 104175
rect 277087 104147 277121 104175
rect 277149 104147 281097 104175
rect 281125 104147 281159 104175
rect 281187 104147 281221 104175
rect 281249 104147 281283 104175
rect 281311 104147 296457 104175
rect 296485 104147 296519 104175
rect 296547 104147 296581 104175
rect 296609 104147 296643 104175
rect 296671 104147 298728 104175
rect 298756 104147 298790 104175
rect 298818 104147 298852 104175
rect 298880 104147 298914 104175
rect 298942 104147 298990 104175
rect -958 104113 298990 104147
rect -958 104085 -910 104113
rect -882 104085 -848 104113
rect -820 104085 -786 104113
rect -758 104085 -724 104113
rect -696 104085 4617 104113
rect 4645 104085 4679 104113
rect 4707 104085 4741 104113
rect 4769 104085 4803 104113
rect 4831 104085 15939 104113
rect 15967 104085 16001 104113
rect 16029 104085 19977 104113
rect 20005 104085 20039 104113
rect 20067 104085 20101 104113
rect 20129 104085 20163 104113
rect 20191 104085 31299 104113
rect 31327 104085 31361 104113
rect 31389 104085 35337 104113
rect 35365 104085 35399 104113
rect 35427 104085 35461 104113
rect 35489 104085 35523 104113
rect 35551 104085 46659 104113
rect 46687 104085 46721 104113
rect 46749 104085 50697 104113
rect 50725 104085 50759 104113
rect 50787 104085 50821 104113
rect 50849 104085 50883 104113
rect 50911 104085 62019 104113
rect 62047 104085 62081 104113
rect 62109 104085 66057 104113
rect 66085 104085 66119 104113
rect 66147 104085 66181 104113
rect 66209 104085 66243 104113
rect 66271 104085 77379 104113
rect 77407 104085 77441 104113
rect 77469 104085 81417 104113
rect 81445 104085 81479 104113
rect 81507 104085 81541 104113
rect 81569 104085 81603 104113
rect 81631 104085 92739 104113
rect 92767 104085 92801 104113
rect 92829 104085 96777 104113
rect 96805 104085 96839 104113
rect 96867 104085 96901 104113
rect 96929 104085 96963 104113
rect 96991 104085 108099 104113
rect 108127 104085 108161 104113
rect 108189 104085 112137 104113
rect 112165 104085 112199 104113
rect 112227 104085 112261 104113
rect 112289 104085 112323 104113
rect 112351 104085 123459 104113
rect 123487 104085 123521 104113
rect 123549 104085 127497 104113
rect 127525 104085 127559 104113
rect 127587 104085 127621 104113
rect 127649 104085 127683 104113
rect 127711 104085 138819 104113
rect 138847 104085 138881 104113
rect 138909 104085 142857 104113
rect 142885 104085 142919 104113
rect 142947 104085 142981 104113
rect 143009 104085 143043 104113
rect 143071 104085 154179 104113
rect 154207 104085 154241 104113
rect 154269 104085 158217 104113
rect 158245 104085 158279 104113
rect 158307 104085 158341 104113
rect 158369 104085 158403 104113
rect 158431 104085 169539 104113
rect 169567 104085 169601 104113
rect 169629 104085 173577 104113
rect 173605 104085 173639 104113
rect 173667 104085 173701 104113
rect 173729 104085 173763 104113
rect 173791 104085 184899 104113
rect 184927 104085 184961 104113
rect 184989 104085 188937 104113
rect 188965 104085 188999 104113
rect 189027 104085 189061 104113
rect 189089 104085 189123 104113
rect 189151 104085 200259 104113
rect 200287 104085 200321 104113
rect 200349 104085 204297 104113
rect 204325 104085 204359 104113
rect 204387 104085 204421 104113
rect 204449 104085 204483 104113
rect 204511 104085 215619 104113
rect 215647 104085 215681 104113
rect 215709 104085 219657 104113
rect 219685 104085 219719 104113
rect 219747 104085 219781 104113
rect 219809 104085 219843 104113
rect 219871 104085 230979 104113
rect 231007 104085 231041 104113
rect 231069 104085 235017 104113
rect 235045 104085 235079 104113
rect 235107 104085 235141 104113
rect 235169 104085 235203 104113
rect 235231 104085 246339 104113
rect 246367 104085 246401 104113
rect 246429 104085 250377 104113
rect 250405 104085 250439 104113
rect 250467 104085 250501 104113
rect 250529 104085 250563 104113
rect 250591 104085 261699 104113
rect 261727 104085 261761 104113
rect 261789 104085 265737 104113
rect 265765 104085 265799 104113
rect 265827 104085 265861 104113
rect 265889 104085 265923 104113
rect 265951 104085 277059 104113
rect 277087 104085 277121 104113
rect 277149 104085 281097 104113
rect 281125 104085 281159 104113
rect 281187 104085 281221 104113
rect 281249 104085 281283 104113
rect 281311 104085 296457 104113
rect 296485 104085 296519 104113
rect 296547 104085 296581 104113
rect 296609 104085 296643 104113
rect 296671 104085 298728 104113
rect 298756 104085 298790 104113
rect 298818 104085 298852 104113
rect 298880 104085 298914 104113
rect 298942 104085 298990 104113
rect -958 104051 298990 104085
rect -958 104023 -910 104051
rect -882 104023 -848 104051
rect -820 104023 -786 104051
rect -758 104023 -724 104051
rect -696 104023 4617 104051
rect 4645 104023 4679 104051
rect 4707 104023 4741 104051
rect 4769 104023 4803 104051
rect 4831 104023 15939 104051
rect 15967 104023 16001 104051
rect 16029 104023 19977 104051
rect 20005 104023 20039 104051
rect 20067 104023 20101 104051
rect 20129 104023 20163 104051
rect 20191 104023 31299 104051
rect 31327 104023 31361 104051
rect 31389 104023 35337 104051
rect 35365 104023 35399 104051
rect 35427 104023 35461 104051
rect 35489 104023 35523 104051
rect 35551 104023 46659 104051
rect 46687 104023 46721 104051
rect 46749 104023 50697 104051
rect 50725 104023 50759 104051
rect 50787 104023 50821 104051
rect 50849 104023 50883 104051
rect 50911 104023 62019 104051
rect 62047 104023 62081 104051
rect 62109 104023 66057 104051
rect 66085 104023 66119 104051
rect 66147 104023 66181 104051
rect 66209 104023 66243 104051
rect 66271 104023 77379 104051
rect 77407 104023 77441 104051
rect 77469 104023 81417 104051
rect 81445 104023 81479 104051
rect 81507 104023 81541 104051
rect 81569 104023 81603 104051
rect 81631 104023 92739 104051
rect 92767 104023 92801 104051
rect 92829 104023 96777 104051
rect 96805 104023 96839 104051
rect 96867 104023 96901 104051
rect 96929 104023 96963 104051
rect 96991 104023 108099 104051
rect 108127 104023 108161 104051
rect 108189 104023 112137 104051
rect 112165 104023 112199 104051
rect 112227 104023 112261 104051
rect 112289 104023 112323 104051
rect 112351 104023 123459 104051
rect 123487 104023 123521 104051
rect 123549 104023 127497 104051
rect 127525 104023 127559 104051
rect 127587 104023 127621 104051
rect 127649 104023 127683 104051
rect 127711 104023 138819 104051
rect 138847 104023 138881 104051
rect 138909 104023 142857 104051
rect 142885 104023 142919 104051
rect 142947 104023 142981 104051
rect 143009 104023 143043 104051
rect 143071 104023 154179 104051
rect 154207 104023 154241 104051
rect 154269 104023 158217 104051
rect 158245 104023 158279 104051
rect 158307 104023 158341 104051
rect 158369 104023 158403 104051
rect 158431 104023 169539 104051
rect 169567 104023 169601 104051
rect 169629 104023 173577 104051
rect 173605 104023 173639 104051
rect 173667 104023 173701 104051
rect 173729 104023 173763 104051
rect 173791 104023 184899 104051
rect 184927 104023 184961 104051
rect 184989 104023 188937 104051
rect 188965 104023 188999 104051
rect 189027 104023 189061 104051
rect 189089 104023 189123 104051
rect 189151 104023 200259 104051
rect 200287 104023 200321 104051
rect 200349 104023 204297 104051
rect 204325 104023 204359 104051
rect 204387 104023 204421 104051
rect 204449 104023 204483 104051
rect 204511 104023 215619 104051
rect 215647 104023 215681 104051
rect 215709 104023 219657 104051
rect 219685 104023 219719 104051
rect 219747 104023 219781 104051
rect 219809 104023 219843 104051
rect 219871 104023 230979 104051
rect 231007 104023 231041 104051
rect 231069 104023 235017 104051
rect 235045 104023 235079 104051
rect 235107 104023 235141 104051
rect 235169 104023 235203 104051
rect 235231 104023 246339 104051
rect 246367 104023 246401 104051
rect 246429 104023 250377 104051
rect 250405 104023 250439 104051
rect 250467 104023 250501 104051
rect 250529 104023 250563 104051
rect 250591 104023 261699 104051
rect 261727 104023 261761 104051
rect 261789 104023 265737 104051
rect 265765 104023 265799 104051
rect 265827 104023 265861 104051
rect 265889 104023 265923 104051
rect 265951 104023 277059 104051
rect 277087 104023 277121 104051
rect 277149 104023 281097 104051
rect 281125 104023 281159 104051
rect 281187 104023 281221 104051
rect 281249 104023 281283 104051
rect 281311 104023 296457 104051
rect 296485 104023 296519 104051
rect 296547 104023 296581 104051
rect 296609 104023 296643 104051
rect 296671 104023 298728 104051
rect 298756 104023 298790 104051
rect 298818 104023 298852 104051
rect 298880 104023 298914 104051
rect 298942 104023 298990 104051
rect -958 103989 298990 104023
rect -958 103961 -910 103989
rect -882 103961 -848 103989
rect -820 103961 -786 103989
rect -758 103961 -724 103989
rect -696 103961 4617 103989
rect 4645 103961 4679 103989
rect 4707 103961 4741 103989
rect 4769 103961 4803 103989
rect 4831 103961 15939 103989
rect 15967 103961 16001 103989
rect 16029 103961 19977 103989
rect 20005 103961 20039 103989
rect 20067 103961 20101 103989
rect 20129 103961 20163 103989
rect 20191 103961 31299 103989
rect 31327 103961 31361 103989
rect 31389 103961 35337 103989
rect 35365 103961 35399 103989
rect 35427 103961 35461 103989
rect 35489 103961 35523 103989
rect 35551 103961 46659 103989
rect 46687 103961 46721 103989
rect 46749 103961 50697 103989
rect 50725 103961 50759 103989
rect 50787 103961 50821 103989
rect 50849 103961 50883 103989
rect 50911 103961 62019 103989
rect 62047 103961 62081 103989
rect 62109 103961 66057 103989
rect 66085 103961 66119 103989
rect 66147 103961 66181 103989
rect 66209 103961 66243 103989
rect 66271 103961 77379 103989
rect 77407 103961 77441 103989
rect 77469 103961 81417 103989
rect 81445 103961 81479 103989
rect 81507 103961 81541 103989
rect 81569 103961 81603 103989
rect 81631 103961 92739 103989
rect 92767 103961 92801 103989
rect 92829 103961 96777 103989
rect 96805 103961 96839 103989
rect 96867 103961 96901 103989
rect 96929 103961 96963 103989
rect 96991 103961 108099 103989
rect 108127 103961 108161 103989
rect 108189 103961 112137 103989
rect 112165 103961 112199 103989
rect 112227 103961 112261 103989
rect 112289 103961 112323 103989
rect 112351 103961 123459 103989
rect 123487 103961 123521 103989
rect 123549 103961 127497 103989
rect 127525 103961 127559 103989
rect 127587 103961 127621 103989
rect 127649 103961 127683 103989
rect 127711 103961 138819 103989
rect 138847 103961 138881 103989
rect 138909 103961 142857 103989
rect 142885 103961 142919 103989
rect 142947 103961 142981 103989
rect 143009 103961 143043 103989
rect 143071 103961 154179 103989
rect 154207 103961 154241 103989
rect 154269 103961 158217 103989
rect 158245 103961 158279 103989
rect 158307 103961 158341 103989
rect 158369 103961 158403 103989
rect 158431 103961 169539 103989
rect 169567 103961 169601 103989
rect 169629 103961 173577 103989
rect 173605 103961 173639 103989
rect 173667 103961 173701 103989
rect 173729 103961 173763 103989
rect 173791 103961 184899 103989
rect 184927 103961 184961 103989
rect 184989 103961 188937 103989
rect 188965 103961 188999 103989
rect 189027 103961 189061 103989
rect 189089 103961 189123 103989
rect 189151 103961 200259 103989
rect 200287 103961 200321 103989
rect 200349 103961 204297 103989
rect 204325 103961 204359 103989
rect 204387 103961 204421 103989
rect 204449 103961 204483 103989
rect 204511 103961 215619 103989
rect 215647 103961 215681 103989
rect 215709 103961 219657 103989
rect 219685 103961 219719 103989
rect 219747 103961 219781 103989
rect 219809 103961 219843 103989
rect 219871 103961 230979 103989
rect 231007 103961 231041 103989
rect 231069 103961 235017 103989
rect 235045 103961 235079 103989
rect 235107 103961 235141 103989
rect 235169 103961 235203 103989
rect 235231 103961 246339 103989
rect 246367 103961 246401 103989
rect 246429 103961 250377 103989
rect 250405 103961 250439 103989
rect 250467 103961 250501 103989
rect 250529 103961 250563 103989
rect 250591 103961 261699 103989
rect 261727 103961 261761 103989
rect 261789 103961 265737 103989
rect 265765 103961 265799 103989
rect 265827 103961 265861 103989
rect 265889 103961 265923 103989
rect 265951 103961 277059 103989
rect 277087 103961 277121 103989
rect 277149 103961 281097 103989
rect 281125 103961 281159 103989
rect 281187 103961 281221 103989
rect 281249 103961 281283 103989
rect 281311 103961 296457 103989
rect 296485 103961 296519 103989
rect 296547 103961 296581 103989
rect 296609 103961 296643 103989
rect 296671 103961 298728 103989
rect 298756 103961 298790 103989
rect 298818 103961 298852 103989
rect 298880 103961 298914 103989
rect 298942 103961 298990 103989
rect -958 103913 298990 103961
rect -958 101175 298990 101223
rect -958 101147 -430 101175
rect -402 101147 -368 101175
rect -340 101147 -306 101175
rect -278 101147 -244 101175
rect -216 101147 2757 101175
rect 2785 101147 2819 101175
rect 2847 101147 2881 101175
rect 2909 101147 2943 101175
rect 2971 101147 8259 101175
rect 8287 101147 8321 101175
rect 8349 101147 18117 101175
rect 18145 101147 18179 101175
rect 18207 101147 18241 101175
rect 18269 101147 18303 101175
rect 18331 101147 23619 101175
rect 23647 101147 23681 101175
rect 23709 101147 33477 101175
rect 33505 101147 33539 101175
rect 33567 101147 33601 101175
rect 33629 101147 33663 101175
rect 33691 101147 38979 101175
rect 39007 101147 39041 101175
rect 39069 101147 48837 101175
rect 48865 101147 48899 101175
rect 48927 101147 48961 101175
rect 48989 101147 49023 101175
rect 49051 101147 54339 101175
rect 54367 101147 54401 101175
rect 54429 101147 64197 101175
rect 64225 101147 64259 101175
rect 64287 101147 64321 101175
rect 64349 101147 64383 101175
rect 64411 101147 69699 101175
rect 69727 101147 69761 101175
rect 69789 101147 79557 101175
rect 79585 101147 79619 101175
rect 79647 101147 79681 101175
rect 79709 101147 79743 101175
rect 79771 101147 85059 101175
rect 85087 101147 85121 101175
rect 85149 101147 94917 101175
rect 94945 101147 94979 101175
rect 95007 101147 95041 101175
rect 95069 101147 95103 101175
rect 95131 101147 100419 101175
rect 100447 101147 100481 101175
rect 100509 101147 110277 101175
rect 110305 101147 110339 101175
rect 110367 101147 110401 101175
rect 110429 101147 110463 101175
rect 110491 101147 115779 101175
rect 115807 101147 115841 101175
rect 115869 101147 125637 101175
rect 125665 101147 125699 101175
rect 125727 101147 125761 101175
rect 125789 101147 125823 101175
rect 125851 101147 131139 101175
rect 131167 101147 131201 101175
rect 131229 101147 140997 101175
rect 141025 101147 141059 101175
rect 141087 101147 141121 101175
rect 141149 101147 141183 101175
rect 141211 101147 146499 101175
rect 146527 101147 146561 101175
rect 146589 101147 156357 101175
rect 156385 101147 156419 101175
rect 156447 101147 156481 101175
rect 156509 101147 156543 101175
rect 156571 101147 161859 101175
rect 161887 101147 161921 101175
rect 161949 101147 171717 101175
rect 171745 101147 171779 101175
rect 171807 101147 171841 101175
rect 171869 101147 171903 101175
rect 171931 101147 177219 101175
rect 177247 101147 177281 101175
rect 177309 101147 187077 101175
rect 187105 101147 187139 101175
rect 187167 101147 187201 101175
rect 187229 101147 187263 101175
rect 187291 101147 192579 101175
rect 192607 101147 192641 101175
rect 192669 101147 202437 101175
rect 202465 101147 202499 101175
rect 202527 101147 202561 101175
rect 202589 101147 202623 101175
rect 202651 101147 207939 101175
rect 207967 101147 208001 101175
rect 208029 101147 217797 101175
rect 217825 101147 217859 101175
rect 217887 101147 217921 101175
rect 217949 101147 217983 101175
rect 218011 101147 223299 101175
rect 223327 101147 223361 101175
rect 223389 101147 233157 101175
rect 233185 101147 233219 101175
rect 233247 101147 233281 101175
rect 233309 101147 233343 101175
rect 233371 101147 238659 101175
rect 238687 101147 238721 101175
rect 238749 101147 248517 101175
rect 248545 101147 248579 101175
rect 248607 101147 248641 101175
rect 248669 101147 248703 101175
rect 248731 101147 254019 101175
rect 254047 101147 254081 101175
rect 254109 101147 263877 101175
rect 263905 101147 263939 101175
rect 263967 101147 264001 101175
rect 264029 101147 264063 101175
rect 264091 101147 269379 101175
rect 269407 101147 269441 101175
rect 269469 101147 279237 101175
rect 279265 101147 279299 101175
rect 279327 101147 279361 101175
rect 279389 101147 279423 101175
rect 279451 101147 284739 101175
rect 284767 101147 284801 101175
rect 284829 101147 294597 101175
rect 294625 101147 294659 101175
rect 294687 101147 294721 101175
rect 294749 101147 294783 101175
rect 294811 101147 298248 101175
rect 298276 101147 298310 101175
rect 298338 101147 298372 101175
rect 298400 101147 298434 101175
rect 298462 101147 298990 101175
rect -958 101113 298990 101147
rect -958 101085 -430 101113
rect -402 101085 -368 101113
rect -340 101085 -306 101113
rect -278 101085 -244 101113
rect -216 101085 2757 101113
rect 2785 101085 2819 101113
rect 2847 101085 2881 101113
rect 2909 101085 2943 101113
rect 2971 101085 8259 101113
rect 8287 101085 8321 101113
rect 8349 101085 18117 101113
rect 18145 101085 18179 101113
rect 18207 101085 18241 101113
rect 18269 101085 18303 101113
rect 18331 101085 23619 101113
rect 23647 101085 23681 101113
rect 23709 101085 33477 101113
rect 33505 101085 33539 101113
rect 33567 101085 33601 101113
rect 33629 101085 33663 101113
rect 33691 101085 38979 101113
rect 39007 101085 39041 101113
rect 39069 101085 48837 101113
rect 48865 101085 48899 101113
rect 48927 101085 48961 101113
rect 48989 101085 49023 101113
rect 49051 101085 54339 101113
rect 54367 101085 54401 101113
rect 54429 101085 64197 101113
rect 64225 101085 64259 101113
rect 64287 101085 64321 101113
rect 64349 101085 64383 101113
rect 64411 101085 69699 101113
rect 69727 101085 69761 101113
rect 69789 101085 79557 101113
rect 79585 101085 79619 101113
rect 79647 101085 79681 101113
rect 79709 101085 79743 101113
rect 79771 101085 85059 101113
rect 85087 101085 85121 101113
rect 85149 101085 94917 101113
rect 94945 101085 94979 101113
rect 95007 101085 95041 101113
rect 95069 101085 95103 101113
rect 95131 101085 100419 101113
rect 100447 101085 100481 101113
rect 100509 101085 110277 101113
rect 110305 101085 110339 101113
rect 110367 101085 110401 101113
rect 110429 101085 110463 101113
rect 110491 101085 115779 101113
rect 115807 101085 115841 101113
rect 115869 101085 125637 101113
rect 125665 101085 125699 101113
rect 125727 101085 125761 101113
rect 125789 101085 125823 101113
rect 125851 101085 131139 101113
rect 131167 101085 131201 101113
rect 131229 101085 140997 101113
rect 141025 101085 141059 101113
rect 141087 101085 141121 101113
rect 141149 101085 141183 101113
rect 141211 101085 146499 101113
rect 146527 101085 146561 101113
rect 146589 101085 156357 101113
rect 156385 101085 156419 101113
rect 156447 101085 156481 101113
rect 156509 101085 156543 101113
rect 156571 101085 161859 101113
rect 161887 101085 161921 101113
rect 161949 101085 171717 101113
rect 171745 101085 171779 101113
rect 171807 101085 171841 101113
rect 171869 101085 171903 101113
rect 171931 101085 177219 101113
rect 177247 101085 177281 101113
rect 177309 101085 187077 101113
rect 187105 101085 187139 101113
rect 187167 101085 187201 101113
rect 187229 101085 187263 101113
rect 187291 101085 192579 101113
rect 192607 101085 192641 101113
rect 192669 101085 202437 101113
rect 202465 101085 202499 101113
rect 202527 101085 202561 101113
rect 202589 101085 202623 101113
rect 202651 101085 207939 101113
rect 207967 101085 208001 101113
rect 208029 101085 217797 101113
rect 217825 101085 217859 101113
rect 217887 101085 217921 101113
rect 217949 101085 217983 101113
rect 218011 101085 223299 101113
rect 223327 101085 223361 101113
rect 223389 101085 233157 101113
rect 233185 101085 233219 101113
rect 233247 101085 233281 101113
rect 233309 101085 233343 101113
rect 233371 101085 238659 101113
rect 238687 101085 238721 101113
rect 238749 101085 248517 101113
rect 248545 101085 248579 101113
rect 248607 101085 248641 101113
rect 248669 101085 248703 101113
rect 248731 101085 254019 101113
rect 254047 101085 254081 101113
rect 254109 101085 263877 101113
rect 263905 101085 263939 101113
rect 263967 101085 264001 101113
rect 264029 101085 264063 101113
rect 264091 101085 269379 101113
rect 269407 101085 269441 101113
rect 269469 101085 279237 101113
rect 279265 101085 279299 101113
rect 279327 101085 279361 101113
rect 279389 101085 279423 101113
rect 279451 101085 284739 101113
rect 284767 101085 284801 101113
rect 284829 101085 294597 101113
rect 294625 101085 294659 101113
rect 294687 101085 294721 101113
rect 294749 101085 294783 101113
rect 294811 101085 298248 101113
rect 298276 101085 298310 101113
rect 298338 101085 298372 101113
rect 298400 101085 298434 101113
rect 298462 101085 298990 101113
rect -958 101051 298990 101085
rect -958 101023 -430 101051
rect -402 101023 -368 101051
rect -340 101023 -306 101051
rect -278 101023 -244 101051
rect -216 101023 2757 101051
rect 2785 101023 2819 101051
rect 2847 101023 2881 101051
rect 2909 101023 2943 101051
rect 2971 101023 8259 101051
rect 8287 101023 8321 101051
rect 8349 101023 18117 101051
rect 18145 101023 18179 101051
rect 18207 101023 18241 101051
rect 18269 101023 18303 101051
rect 18331 101023 23619 101051
rect 23647 101023 23681 101051
rect 23709 101023 33477 101051
rect 33505 101023 33539 101051
rect 33567 101023 33601 101051
rect 33629 101023 33663 101051
rect 33691 101023 38979 101051
rect 39007 101023 39041 101051
rect 39069 101023 48837 101051
rect 48865 101023 48899 101051
rect 48927 101023 48961 101051
rect 48989 101023 49023 101051
rect 49051 101023 54339 101051
rect 54367 101023 54401 101051
rect 54429 101023 64197 101051
rect 64225 101023 64259 101051
rect 64287 101023 64321 101051
rect 64349 101023 64383 101051
rect 64411 101023 69699 101051
rect 69727 101023 69761 101051
rect 69789 101023 79557 101051
rect 79585 101023 79619 101051
rect 79647 101023 79681 101051
rect 79709 101023 79743 101051
rect 79771 101023 85059 101051
rect 85087 101023 85121 101051
rect 85149 101023 94917 101051
rect 94945 101023 94979 101051
rect 95007 101023 95041 101051
rect 95069 101023 95103 101051
rect 95131 101023 100419 101051
rect 100447 101023 100481 101051
rect 100509 101023 110277 101051
rect 110305 101023 110339 101051
rect 110367 101023 110401 101051
rect 110429 101023 110463 101051
rect 110491 101023 115779 101051
rect 115807 101023 115841 101051
rect 115869 101023 125637 101051
rect 125665 101023 125699 101051
rect 125727 101023 125761 101051
rect 125789 101023 125823 101051
rect 125851 101023 131139 101051
rect 131167 101023 131201 101051
rect 131229 101023 140997 101051
rect 141025 101023 141059 101051
rect 141087 101023 141121 101051
rect 141149 101023 141183 101051
rect 141211 101023 146499 101051
rect 146527 101023 146561 101051
rect 146589 101023 156357 101051
rect 156385 101023 156419 101051
rect 156447 101023 156481 101051
rect 156509 101023 156543 101051
rect 156571 101023 161859 101051
rect 161887 101023 161921 101051
rect 161949 101023 171717 101051
rect 171745 101023 171779 101051
rect 171807 101023 171841 101051
rect 171869 101023 171903 101051
rect 171931 101023 177219 101051
rect 177247 101023 177281 101051
rect 177309 101023 187077 101051
rect 187105 101023 187139 101051
rect 187167 101023 187201 101051
rect 187229 101023 187263 101051
rect 187291 101023 192579 101051
rect 192607 101023 192641 101051
rect 192669 101023 202437 101051
rect 202465 101023 202499 101051
rect 202527 101023 202561 101051
rect 202589 101023 202623 101051
rect 202651 101023 207939 101051
rect 207967 101023 208001 101051
rect 208029 101023 217797 101051
rect 217825 101023 217859 101051
rect 217887 101023 217921 101051
rect 217949 101023 217983 101051
rect 218011 101023 223299 101051
rect 223327 101023 223361 101051
rect 223389 101023 233157 101051
rect 233185 101023 233219 101051
rect 233247 101023 233281 101051
rect 233309 101023 233343 101051
rect 233371 101023 238659 101051
rect 238687 101023 238721 101051
rect 238749 101023 248517 101051
rect 248545 101023 248579 101051
rect 248607 101023 248641 101051
rect 248669 101023 248703 101051
rect 248731 101023 254019 101051
rect 254047 101023 254081 101051
rect 254109 101023 263877 101051
rect 263905 101023 263939 101051
rect 263967 101023 264001 101051
rect 264029 101023 264063 101051
rect 264091 101023 269379 101051
rect 269407 101023 269441 101051
rect 269469 101023 279237 101051
rect 279265 101023 279299 101051
rect 279327 101023 279361 101051
rect 279389 101023 279423 101051
rect 279451 101023 284739 101051
rect 284767 101023 284801 101051
rect 284829 101023 294597 101051
rect 294625 101023 294659 101051
rect 294687 101023 294721 101051
rect 294749 101023 294783 101051
rect 294811 101023 298248 101051
rect 298276 101023 298310 101051
rect 298338 101023 298372 101051
rect 298400 101023 298434 101051
rect 298462 101023 298990 101051
rect -958 100989 298990 101023
rect -958 100961 -430 100989
rect -402 100961 -368 100989
rect -340 100961 -306 100989
rect -278 100961 -244 100989
rect -216 100961 2757 100989
rect 2785 100961 2819 100989
rect 2847 100961 2881 100989
rect 2909 100961 2943 100989
rect 2971 100961 8259 100989
rect 8287 100961 8321 100989
rect 8349 100961 18117 100989
rect 18145 100961 18179 100989
rect 18207 100961 18241 100989
rect 18269 100961 18303 100989
rect 18331 100961 23619 100989
rect 23647 100961 23681 100989
rect 23709 100961 33477 100989
rect 33505 100961 33539 100989
rect 33567 100961 33601 100989
rect 33629 100961 33663 100989
rect 33691 100961 38979 100989
rect 39007 100961 39041 100989
rect 39069 100961 48837 100989
rect 48865 100961 48899 100989
rect 48927 100961 48961 100989
rect 48989 100961 49023 100989
rect 49051 100961 54339 100989
rect 54367 100961 54401 100989
rect 54429 100961 64197 100989
rect 64225 100961 64259 100989
rect 64287 100961 64321 100989
rect 64349 100961 64383 100989
rect 64411 100961 69699 100989
rect 69727 100961 69761 100989
rect 69789 100961 79557 100989
rect 79585 100961 79619 100989
rect 79647 100961 79681 100989
rect 79709 100961 79743 100989
rect 79771 100961 85059 100989
rect 85087 100961 85121 100989
rect 85149 100961 94917 100989
rect 94945 100961 94979 100989
rect 95007 100961 95041 100989
rect 95069 100961 95103 100989
rect 95131 100961 100419 100989
rect 100447 100961 100481 100989
rect 100509 100961 110277 100989
rect 110305 100961 110339 100989
rect 110367 100961 110401 100989
rect 110429 100961 110463 100989
rect 110491 100961 115779 100989
rect 115807 100961 115841 100989
rect 115869 100961 125637 100989
rect 125665 100961 125699 100989
rect 125727 100961 125761 100989
rect 125789 100961 125823 100989
rect 125851 100961 131139 100989
rect 131167 100961 131201 100989
rect 131229 100961 140997 100989
rect 141025 100961 141059 100989
rect 141087 100961 141121 100989
rect 141149 100961 141183 100989
rect 141211 100961 146499 100989
rect 146527 100961 146561 100989
rect 146589 100961 156357 100989
rect 156385 100961 156419 100989
rect 156447 100961 156481 100989
rect 156509 100961 156543 100989
rect 156571 100961 161859 100989
rect 161887 100961 161921 100989
rect 161949 100961 171717 100989
rect 171745 100961 171779 100989
rect 171807 100961 171841 100989
rect 171869 100961 171903 100989
rect 171931 100961 177219 100989
rect 177247 100961 177281 100989
rect 177309 100961 187077 100989
rect 187105 100961 187139 100989
rect 187167 100961 187201 100989
rect 187229 100961 187263 100989
rect 187291 100961 192579 100989
rect 192607 100961 192641 100989
rect 192669 100961 202437 100989
rect 202465 100961 202499 100989
rect 202527 100961 202561 100989
rect 202589 100961 202623 100989
rect 202651 100961 207939 100989
rect 207967 100961 208001 100989
rect 208029 100961 217797 100989
rect 217825 100961 217859 100989
rect 217887 100961 217921 100989
rect 217949 100961 217983 100989
rect 218011 100961 223299 100989
rect 223327 100961 223361 100989
rect 223389 100961 233157 100989
rect 233185 100961 233219 100989
rect 233247 100961 233281 100989
rect 233309 100961 233343 100989
rect 233371 100961 238659 100989
rect 238687 100961 238721 100989
rect 238749 100961 248517 100989
rect 248545 100961 248579 100989
rect 248607 100961 248641 100989
rect 248669 100961 248703 100989
rect 248731 100961 254019 100989
rect 254047 100961 254081 100989
rect 254109 100961 263877 100989
rect 263905 100961 263939 100989
rect 263967 100961 264001 100989
rect 264029 100961 264063 100989
rect 264091 100961 269379 100989
rect 269407 100961 269441 100989
rect 269469 100961 279237 100989
rect 279265 100961 279299 100989
rect 279327 100961 279361 100989
rect 279389 100961 279423 100989
rect 279451 100961 284739 100989
rect 284767 100961 284801 100989
rect 284829 100961 294597 100989
rect 294625 100961 294659 100989
rect 294687 100961 294721 100989
rect 294749 100961 294783 100989
rect 294811 100961 298248 100989
rect 298276 100961 298310 100989
rect 298338 100961 298372 100989
rect 298400 100961 298434 100989
rect 298462 100961 298990 100989
rect -958 100913 298990 100961
rect -958 95175 298990 95223
rect -958 95147 -910 95175
rect -882 95147 -848 95175
rect -820 95147 -786 95175
rect -758 95147 -724 95175
rect -696 95147 4617 95175
rect 4645 95147 4679 95175
rect 4707 95147 4741 95175
rect 4769 95147 4803 95175
rect 4831 95147 15939 95175
rect 15967 95147 16001 95175
rect 16029 95147 19977 95175
rect 20005 95147 20039 95175
rect 20067 95147 20101 95175
rect 20129 95147 20163 95175
rect 20191 95147 31299 95175
rect 31327 95147 31361 95175
rect 31389 95147 35337 95175
rect 35365 95147 35399 95175
rect 35427 95147 35461 95175
rect 35489 95147 35523 95175
rect 35551 95147 46659 95175
rect 46687 95147 46721 95175
rect 46749 95147 50697 95175
rect 50725 95147 50759 95175
rect 50787 95147 50821 95175
rect 50849 95147 50883 95175
rect 50911 95147 62019 95175
rect 62047 95147 62081 95175
rect 62109 95147 66057 95175
rect 66085 95147 66119 95175
rect 66147 95147 66181 95175
rect 66209 95147 66243 95175
rect 66271 95147 77379 95175
rect 77407 95147 77441 95175
rect 77469 95147 81417 95175
rect 81445 95147 81479 95175
rect 81507 95147 81541 95175
rect 81569 95147 81603 95175
rect 81631 95147 92739 95175
rect 92767 95147 92801 95175
rect 92829 95147 96777 95175
rect 96805 95147 96839 95175
rect 96867 95147 96901 95175
rect 96929 95147 96963 95175
rect 96991 95147 108099 95175
rect 108127 95147 108161 95175
rect 108189 95147 112137 95175
rect 112165 95147 112199 95175
rect 112227 95147 112261 95175
rect 112289 95147 112323 95175
rect 112351 95147 123459 95175
rect 123487 95147 123521 95175
rect 123549 95147 127497 95175
rect 127525 95147 127559 95175
rect 127587 95147 127621 95175
rect 127649 95147 127683 95175
rect 127711 95147 138819 95175
rect 138847 95147 138881 95175
rect 138909 95147 142857 95175
rect 142885 95147 142919 95175
rect 142947 95147 142981 95175
rect 143009 95147 143043 95175
rect 143071 95147 154179 95175
rect 154207 95147 154241 95175
rect 154269 95147 158217 95175
rect 158245 95147 158279 95175
rect 158307 95147 158341 95175
rect 158369 95147 158403 95175
rect 158431 95147 169539 95175
rect 169567 95147 169601 95175
rect 169629 95147 173577 95175
rect 173605 95147 173639 95175
rect 173667 95147 173701 95175
rect 173729 95147 173763 95175
rect 173791 95147 184899 95175
rect 184927 95147 184961 95175
rect 184989 95147 188937 95175
rect 188965 95147 188999 95175
rect 189027 95147 189061 95175
rect 189089 95147 189123 95175
rect 189151 95147 200259 95175
rect 200287 95147 200321 95175
rect 200349 95147 204297 95175
rect 204325 95147 204359 95175
rect 204387 95147 204421 95175
rect 204449 95147 204483 95175
rect 204511 95147 215619 95175
rect 215647 95147 215681 95175
rect 215709 95147 219657 95175
rect 219685 95147 219719 95175
rect 219747 95147 219781 95175
rect 219809 95147 219843 95175
rect 219871 95147 230979 95175
rect 231007 95147 231041 95175
rect 231069 95147 235017 95175
rect 235045 95147 235079 95175
rect 235107 95147 235141 95175
rect 235169 95147 235203 95175
rect 235231 95147 246339 95175
rect 246367 95147 246401 95175
rect 246429 95147 250377 95175
rect 250405 95147 250439 95175
rect 250467 95147 250501 95175
rect 250529 95147 250563 95175
rect 250591 95147 261699 95175
rect 261727 95147 261761 95175
rect 261789 95147 265737 95175
rect 265765 95147 265799 95175
rect 265827 95147 265861 95175
rect 265889 95147 265923 95175
rect 265951 95147 277059 95175
rect 277087 95147 277121 95175
rect 277149 95147 281097 95175
rect 281125 95147 281159 95175
rect 281187 95147 281221 95175
rect 281249 95147 281283 95175
rect 281311 95147 296457 95175
rect 296485 95147 296519 95175
rect 296547 95147 296581 95175
rect 296609 95147 296643 95175
rect 296671 95147 298728 95175
rect 298756 95147 298790 95175
rect 298818 95147 298852 95175
rect 298880 95147 298914 95175
rect 298942 95147 298990 95175
rect -958 95113 298990 95147
rect -958 95085 -910 95113
rect -882 95085 -848 95113
rect -820 95085 -786 95113
rect -758 95085 -724 95113
rect -696 95085 4617 95113
rect 4645 95085 4679 95113
rect 4707 95085 4741 95113
rect 4769 95085 4803 95113
rect 4831 95085 15939 95113
rect 15967 95085 16001 95113
rect 16029 95085 19977 95113
rect 20005 95085 20039 95113
rect 20067 95085 20101 95113
rect 20129 95085 20163 95113
rect 20191 95085 31299 95113
rect 31327 95085 31361 95113
rect 31389 95085 35337 95113
rect 35365 95085 35399 95113
rect 35427 95085 35461 95113
rect 35489 95085 35523 95113
rect 35551 95085 46659 95113
rect 46687 95085 46721 95113
rect 46749 95085 50697 95113
rect 50725 95085 50759 95113
rect 50787 95085 50821 95113
rect 50849 95085 50883 95113
rect 50911 95085 62019 95113
rect 62047 95085 62081 95113
rect 62109 95085 66057 95113
rect 66085 95085 66119 95113
rect 66147 95085 66181 95113
rect 66209 95085 66243 95113
rect 66271 95085 77379 95113
rect 77407 95085 77441 95113
rect 77469 95085 81417 95113
rect 81445 95085 81479 95113
rect 81507 95085 81541 95113
rect 81569 95085 81603 95113
rect 81631 95085 92739 95113
rect 92767 95085 92801 95113
rect 92829 95085 96777 95113
rect 96805 95085 96839 95113
rect 96867 95085 96901 95113
rect 96929 95085 96963 95113
rect 96991 95085 108099 95113
rect 108127 95085 108161 95113
rect 108189 95085 112137 95113
rect 112165 95085 112199 95113
rect 112227 95085 112261 95113
rect 112289 95085 112323 95113
rect 112351 95085 123459 95113
rect 123487 95085 123521 95113
rect 123549 95085 127497 95113
rect 127525 95085 127559 95113
rect 127587 95085 127621 95113
rect 127649 95085 127683 95113
rect 127711 95085 138819 95113
rect 138847 95085 138881 95113
rect 138909 95085 142857 95113
rect 142885 95085 142919 95113
rect 142947 95085 142981 95113
rect 143009 95085 143043 95113
rect 143071 95085 154179 95113
rect 154207 95085 154241 95113
rect 154269 95085 158217 95113
rect 158245 95085 158279 95113
rect 158307 95085 158341 95113
rect 158369 95085 158403 95113
rect 158431 95085 169539 95113
rect 169567 95085 169601 95113
rect 169629 95085 173577 95113
rect 173605 95085 173639 95113
rect 173667 95085 173701 95113
rect 173729 95085 173763 95113
rect 173791 95085 184899 95113
rect 184927 95085 184961 95113
rect 184989 95085 188937 95113
rect 188965 95085 188999 95113
rect 189027 95085 189061 95113
rect 189089 95085 189123 95113
rect 189151 95085 200259 95113
rect 200287 95085 200321 95113
rect 200349 95085 204297 95113
rect 204325 95085 204359 95113
rect 204387 95085 204421 95113
rect 204449 95085 204483 95113
rect 204511 95085 215619 95113
rect 215647 95085 215681 95113
rect 215709 95085 219657 95113
rect 219685 95085 219719 95113
rect 219747 95085 219781 95113
rect 219809 95085 219843 95113
rect 219871 95085 230979 95113
rect 231007 95085 231041 95113
rect 231069 95085 235017 95113
rect 235045 95085 235079 95113
rect 235107 95085 235141 95113
rect 235169 95085 235203 95113
rect 235231 95085 246339 95113
rect 246367 95085 246401 95113
rect 246429 95085 250377 95113
rect 250405 95085 250439 95113
rect 250467 95085 250501 95113
rect 250529 95085 250563 95113
rect 250591 95085 261699 95113
rect 261727 95085 261761 95113
rect 261789 95085 265737 95113
rect 265765 95085 265799 95113
rect 265827 95085 265861 95113
rect 265889 95085 265923 95113
rect 265951 95085 277059 95113
rect 277087 95085 277121 95113
rect 277149 95085 281097 95113
rect 281125 95085 281159 95113
rect 281187 95085 281221 95113
rect 281249 95085 281283 95113
rect 281311 95085 296457 95113
rect 296485 95085 296519 95113
rect 296547 95085 296581 95113
rect 296609 95085 296643 95113
rect 296671 95085 298728 95113
rect 298756 95085 298790 95113
rect 298818 95085 298852 95113
rect 298880 95085 298914 95113
rect 298942 95085 298990 95113
rect -958 95051 298990 95085
rect -958 95023 -910 95051
rect -882 95023 -848 95051
rect -820 95023 -786 95051
rect -758 95023 -724 95051
rect -696 95023 4617 95051
rect 4645 95023 4679 95051
rect 4707 95023 4741 95051
rect 4769 95023 4803 95051
rect 4831 95023 15939 95051
rect 15967 95023 16001 95051
rect 16029 95023 19977 95051
rect 20005 95023 20039 95051
rect 20067 95023 20101 95051
rect 20129 95023 20163 95051
rect 20191 95023 31299 95051
rect 31327 95023 31361 95051
rect 31389 95023 35337 95051
rect 35365 95023 35399 95051
rect 35427 95023 35461 95051
rect 35489 95023 35523 95051
rect 35551 95023 46659 95051
rect 46687 95023 46721 95051
rect 46749 95023 50697 95051
rect 50725 95023 50759 95051
rect 50787 95023 50821 95051
rect 50849 95023 50883 95051
rect 50911 95023 62019 95051
rect 62047 95023 62081 95051
rect 62109 95023 66057 95051
rect 66085 95023 66119 95051
rect 66147 95023 66181 95051
rect 66209 95023 66243 95051
rect 66271 95023 77379 95051
rect 77407 95023 77441 95051
rect 77469 95023 81417 95051
rect 81445 95023 81479 95051
rect 81507 95023 81541 95051
rect 81569 95023 81603 95051
rect 81631 95023 92739 95051
rect 92767 95023 92801 95051
rect 92829 95023 96777 95051
rect 96805 95023 96839 95051
rect 96867 95023 96901 95051
rect 96929 95023 96963 95051
rect 96991 95023 108099 95051
rect 108127 95023 108161 95051
rect 108189 95023 112137 95051
rect 112165 95023 112199 95051
rect 112227 95023 112261 95051
rect 112289 95023 112323 95051
rect 112351 95023 123459 95051
rect 123487 95023 123521 95051
rect 123549 95023 127497 95051
rect 127525 95023 127559 95051
rect 127587 95023 127621 95051
rect 127649 95023 127683 95051
rect 127711 95023 138819 95051
rect 138847 95023 138881 95051
rect 138909 95023 142857 95051
rect 142885 95023 142919 95051
rect 142947 95023 142981 95051
rect 143009 95023 143043 95051
rect 143071 95023 154179 95051
rect 154207 95023 154241 95051
rect 154269 95023 158217 95051
rect 158245 95023 158279 95051
rect 158307 95023 158341 95051
rect 158369 95023 158403 95051
rect 158431 95023 169539 95051
rect 169567 95023 169601 95051
rect 169629 95023 173577 95051
rect 173605 95023 173639 95051
rect 173667 95023 173701 95051
rect 173729 95023 173763 95051
rect 173791 95023 184899 95051
rect 184927 95023 184961 95051
rect 184989 95023 188937 95051
rect 188965 95023 188999 95051
rect 189027 95023 189061 95051
rect 189089 95023 189123 95051
rect 189151 95023 200259 95051
rect 200287 95023 200321 95051
rect 200349 95023 204297 95051
rect 204325 95023 204359 95051
rect 204387 95023 204421 95051
rect 204449 95023 204483 95051
rect 204511 95023 215619 95051
rect 215647 95023 215681 95051
rect 215709 95023 219657 95051
rect 219685 95023 219719 95051
rect 219747 95023 219781 95051
rect 219809 95023 219843 95051
rect 219871 95023 230979 95051
rect 231007 95023 231041 95051
rect 231069 95023 235017 95051
rect 235045 95023 235079 95051
rect 235107 95023 235141 95051
rect 235169 95023 235203 95051
rect 235231 95023 246339 95051
rect 246367 95023 246401 95051
rect 246429 95023 250377 95051
rect 250405 95023 250439 95051
rect 250467 95023 250501 95051
rect 250529 95023 250563 95051
rect 250591 95023 261699 95051
rect 261727 95023 261761 95051
rect 261789 95023 265737 95051
rect 265765 95023 265799 95051
rect 265827 95023 265861 95051
rect 265889 95023 265923 95051
rect 265951 95023 277059 95051
rect 277087 95023 277121 95051
rect 277149 95023 281097 95051
rect 281125 95023 281159 95051
rect 281187 95023 281221 95051
rect 281249 95023 281283 95051
rect 281311 95023 296457 95051
rect 296485 95023 296519 95051
rect 296547 95023 296581 95051
rect 296609 95023 296643 95051
rect 296671 95023 298728 95051
rect 298756 95023 298790 95051
rect 298818 95023 298852 95051
rect 298880 95023 298914 95051
rect 298942 95023 298990 95051
rect -958 94989 298990 95023
rect -958 94961 -910 94989
rect -882 94961 -848 94989
rect -820 94961 -786 94989
rect -758 94961 -724 94989
rect -696 94961 4617 94989
rect 4645 94961 4679 94989
rect 4707 94961 4741 94989
rect 4769 94961 4803 94989
rect 4831 94961 15939 94989
rect 15967 94961 16001 94989
rect 16029 94961 19977 94989
rect 20005 94961 20039 94989
rect 20067 94961 20101 94989
rect 20129 94961 20163 94989
rect 20191 94961 31299 94989
rect 31327 94961 31361 94989
rect 31389 94961 35337 94989
rect 35365 94961 35399 94989
rect 35427 94961 35461 94989
rect 35489 94961 35523 94989
rect 35551 94961 46659 94989
rect 46687 94961 46721 94989
rect 46749 94961 50697 94989
rect 50725 94961 50759 94989
rect 50787 94961 50821 94989
rect 50849 94961 50883 94989
rect 50911 94961 62019 94989
rect 62047 94961 62081 94989
rect 62109 94961 66057 94989
rect 66085 94961 66119 94989
rect 66147 94961 66181 94989
rect 66209 94961 66243 94989
rect 66271 94961 77379 94989
rect 77407 94961 77441 94989
rect 77469 94961 81417 94989
rect 81445 94961 81479 94989
rect 81507 94961 81541 94989
rect 81569 94961 81603 94989
rect 81631 94961 92739 94989
rect 92767 94961 92801 94989
rect 92829 94961 96777 94989
rect 96805 94961 96839 94989
rect 96867 94961 96901 94989
rect 96929 94961 96963 94989
rect 96991 94961 108099 94989
rect 108127 94961 108161 94989
rect 108189 94961 112137 94989
rect 112165 94961 112199 94989
rect 112227 94961 112261 94989
rect 112289 94961 112323 94989
rect 112351 94961 123459 94989
rect 123487 94961 123521 94989
rect 123549 94961 127497 94989
rect 127525 94961 127559 94989
rect 127587 94961 127621 94989
rect 127649 94961 127683 94989
rect 127711 94961 138819 94989
rect 138847 94961 138881 94989
rect 138909 94961 142857 94989
rect 142885 94961 142919 94989
rect 142947 94961 142981 94989
rect 143009 94961 143043 94989
rect 143071 94961 154179 94989
rect 154207 94961 154241 94989
rect 154269 94961 158217 94989
rect 158245 94961 158279 94989
rect 158307 94961 158341 94989
rect 158369 94961 158403 94989
rect 158431 94961 169539 94989
rect 169567 94961 169601 94989
rect 169629 94961 173577 94989
rect 173605 94961 173639 94989
rect 173667 94961 173701 94989
rect 173729 94961 173763 94989
rect 173791 94961 184899 94989
rect 184927 94961 184961 94989
rect 184989 94961 188937 94989
rect 188965 94961 188999 94989
rect 189027 94961 189061 94989
rect 189089 94961 189123 94989
rect 189151 94961 200259 94989
rect 200287 94961 200321 94989
rect 200349 94961 204297 94989
rect 204325 94961 204359 94989
rect 204387 94961 204421 94989
rect 204449 94961 204483 94989
rect 204511 94961 215619 94989
rect 215647 94961 215681 94989
rect 215709 94961 219657 94989
rect 219685 94961 219719 94989
rect 219747 94961 219781 94989
rect 219809 94961 219843 94989
rect 219871 94961 230979 94989
rect 231007 94961 231041 94989
rect 231069 94961 235017 94989
rect 235045 94961 235079 94989
rect 235107 94961 235141 94989
rect 235169 94961 235203 94989
rect 235231 94961 246339 94989
rect 246367 94961 246401 94989
rect 246429 94961 250377 94989
rect 250405 94961 250439 94989
rect 250467 94961 250501 94989
rect 250529 94961 250563 94989
rect 250591 94961 261699 94989
rect 261727 94961 261761 94989
rect 261789 94961 265737 94989
rect 265765 94961 265799 94989
rect 265827 94961 265861 94989
rect 265889 94961 265923 94989
rect 265951 94961 277059 94989
rect 277087 94961 277121 94989
rect 277149 94961 281097 94989
rect 281125 94961 281159 94989
rect 281187 94961 281221 94989
rect 281249 94961 281283 94989
rect 281311 94961 296457 94989
rect 296485 94961 296519 94989
rect 296547 94961 296581 94989
rect 296609 94961 296643 94989
rect 296671 94961 298728 94989
rect 298756 94961 298790 94989
rect 298818 94961 298852 94989
rect 298880 94961 298914 94989
rect 298942 94961 298990 94989
rect -958 94913 298990 94961
rect -958 92175 298990 92223
rect -958 92147 -430 92175
rect -402 92147 -368 92175
rect -340 92147 -306 92175
rect -278 92147 -244 92175
rect -216 92147 2757 92175
rect 2785 92147 2819 92175
rect 2847 92147 2881 92175
rect 2909 92147 2943 92175
rect 2971 92147 8259 92175
rect 8287 92147 8321 92175
rect 8349 92147 18117 92175
rect 18145 92147 18179 92175
rect 18207 92147 18241 92175
rect 18269 92147 18303 92175
rect 18331 92147 23619 92175
rect 23647 92147 23681 92175
rect 23709 92147 33477 92175
rect 33505 92147 33539 92175
rect 33567 92147 33601 92175
rect 33629 92147 33663 92175
rect 33691 92147 38979 92175
rect 39007 92147 39041 92175
rect 39069 92147 48837 92175
rect 48865 92147 48899 92175
rect 48927 92147 48961 92175
rect 48989 92147 49023 92175
rect 49051 92147 54339 92175
rect 54367 92147 54401 92175
rect 54429 92147 64197 92175
rect 64225 92147 64259 92175
rect 64287 92147 64321 92175
rect 64349 92147 64383 92175
rect 64411 92147 69699 92175
rect 69727 92147 69761 92175
rect 69789 92147 79557 92175
rect 79585 92147 79619 92175
rect 79647 92147 79681 92175
rect 79709 92147 79743 92175
rect 79771 92147 85059 92175
rect 85087 92147 85121 92175
rect 85149 92147 94917 92175
rect 94945 92147 94979 92175
rect 95007 92147 95041 92175
rect 95069 92147 95103 92175
rect 95131 92147 100419 92175
rect 100447 92147 100481 92175
rect 100509 92147 110277 92175
rect 110305 92147 110339 92175
rect 110367 92147 110401 92175
rect 110429 92147 110463 92175
rect 110491 92147 115779 92175
rect 115807 92147 115841 92175
rect 115869 92147 125637 92175
rect 125665 92147 125699 92175
rect 125727 92147 125761 92175
rect 125789 92147 125823 92175
rect 125851 92147 131139 92175
rect 131167 92147 131201 92175
rect 131229 92147 140997 92175
rect 141025 92147 141059 92175
rect 141087 92147 141121 92175
rect 141149 92147 141183 92175
rect 141211 92147 146499 92175
rect 146527 92147 146561 92175
rect 146589 92147 156357 92175
rect 156385 92147 156419 92175
rect 156447 92147 156481 92175
rect 156509 92147 156543 92175
rect 156571 92147 161859 92175
rect 161887 92147 161921 92175
rect 161949 92147 171717 92175
rect 171745 92147 171779 92175
rect 171807 92147 171841 92175
rect 171869 92147 171903 92175
rect 171931 92147 177219 92175
rect 177247 92147 177281 92175
rect 177309 92147 187077 92175
rect 187105 92147 187139 92175
rect 187167 92147 187201 92175
rect 187229 92147 187263 92175
rect 187291 92147 192579 92175
rect 192607 92147 192641 92175
rect 192669 92147 202437 92175
rect 202465 92147 202499 92175
rect 202527 92147 202561 92175
rect 202589 92147 202623 92175
rect 202651 92147 207939 92175
rect 207967 92147 208001 92175
rect 208029 92147 217797 92175
rect 217825 92147 217859 92175
rect 217887 92147 217921 92175
rect 217949 92147 217983 92175
rect 218011 92147 223299 92175
rect 223327 92147 223361 92175
rect 223389 92147 233157 92175
rect 233185 92147 233219 92175
rect 233247 92147 233281 92175
rect 233309 92147 233343 92175
rect 233371 92147 238659 92175
rect 238687 92147 238721 92175
rect 238749 92147 248517 92175
rect 248545 92147 248579 92175
rect 248607 92147 248641 92175
rect 248669 92147 248703 92175
rect 248731 92147 254019 92175
rect 254047 92147 254081 92175
rect 254109 92147 263877 92175
rect 263905 92147 263939 92175
rect 263967 92147 264001 92175
rect 264029 92147 264063 92175
rect 264091 92147 269379 92175
rect 269407 92147 269441 92175
rect 269469 92147 279237 92175
rect 279265 92147 279299 92175
rect 279327 92147 279361 92175
rect 279389 92147 279423 92175
rect 279451 92147 284739 92175
rect 284767 92147 284801 92175
rect 284829 92147 294597 92175
rect 294625 92147 294659 92175
rect 294687 92147 294721 92175
rect 294749 92147 294783 92175
rect 294811 92147 298248 92175
rect 298276 92147 298310 92175
rect 298338 92147 298372 92175
rect 298400 92147 298434 92175
rect 298462 92147 298990 92175
rect -958 92113 298990 92147
rect -958 92085 -430 92113
rect -402 92085 -368 92113
rect -340 92085 -306 92113
rect -278 92085 -244 92113
rect -216 92085 2757 92113
rect 2785 92085 2819 92113
rect 2847 92085 2881 92113
rect 2909 92085 2943 92113
rect 2971 92085 8259 92113
rect 8287 92085 8321 92113
rect 8349 92085 18117 92113
rect 18145 92085 18179 92113
rect 18207 92085 18241 92113
rect 18269 92085 18303 92113
rect 18331 92085 23619 92113
rect 23647 92085 23681 92113
rect 23709 92085 33477 92113
rect 33505 92085 33539 92113
rect 33567 92085 33601 92113
rect 33629 92085 33663 92113
rect 33691 92085 38979 92113
rect 39007 92085 39041 92113
rect 39069 92085 48837 92113
rect 48865 92085 48899 92113
rect 48927 92085 48961 92113
rect 48989 92085 49023 92113
rect 49051 92085 54339 92113
rect 54367 92085 54401 92113
rect 54429 92085 64197 92113
rect 64225 92085 64259 92113
rect 64287 92085 64321 92113
rect 64349 92085 64383 92113
rect 64411 92085 69699 92113
rect 69727 92085 69761 92113
rect 69789 92085 79557 92113
rect 79585 92085 79619 92113
rect 79647 92085 79681 92113
rect 79709 92085 79743 92113
rect 79771 92085 85059 92113
rect 85087 92085 85121 92113
rect 85149 92085 94917 92113
rect 94945 92085 94979 92113
rect 95007 92085 95041 92113
rect 95069 92085 95103 92113
rect 95131 92085 100419 92113
rect 100447 92085 100481 92113
rect 100509 92085 110277 92113
rect 110305 92085 110339 92113
rect 110367 92085 110401 92113
rect 110429 92085 110463 92113
rect 110491 92085 115779 92113
rect 115807 92085 115841 92113
rect 115869 92085 125637 92113
rect 125665 92085 125699 92113
rect 125727 92085 125761 92113
rect 125789 92085 125823 92113
rect 125851 92085 131139 92113
rect 131167 92085 131201 92113
rect 131229 92085 140997 92113
rect 141025 92085 141059 92113
rect 141087 92085 141121 92113
rect 141149 92085 141183 92113
rect 141211 92085 146499 92113
rect 146527 92085 146561 92113
rect 146589 92085 156357 92113
rect 156385 92085 156419 92113
rect 156447 92085 156481 92113
rect 156509 92085 156543 92113
rect 156571 92085 161859 92113
rect 161887 92085 161921 92113
rect 161949 92085 171717 92113
rect 171745 92085 171779 92113
rect 171807 92085 171841 92113
rect 171869 92085 171903 92113
rect 171931 92085 177219 92113
rect 177247 92085 177281 92113
rect 177309 92085 187077 92113
rect 187105 92085 187139 92113
rect 187167 92085 187201 92113
rect 187229 92085 187263 92113
rect 187291 92085 192579 92113
rect 192607 92085 192641 92113
rect 192669 92085 202437 92113
rect 202465 92085 202499 92113
rect 202527 92085 202561 92113
rect 202589 92085 202623 92113
rect 202651 92085 207939 92113
rect 207967 92085 208001 92113
rect 208029 92085 217797 92113
rect 217825 92085 217859 92113
rect 217887 92085 217921 92113
rect 217949 92085 217983 92113
rect 218011 92085 223299 92113
rect 223327 92085 223361 92113
rect 223389 92085 233157 92113
rect 233185 92085 233219 92113
rect 233247 92085 233281 92113
rect 233309 92085 233343 92113
rect 233371 92085 238659 92113
rect 238687 92085 238721 92113
rect 238749 92085 248517 92113
rect 248545 92085 248579 92113
rect 248607 92085 248641 92113
rect 248669 92085 248703 92113
rect 248731 92085 254019 92113
rect 254047 92085 254081 92113
rect 254109 92085 263877 92113
rect 263905 92085 263939 92113
rect 263967 92085 264001 92113
rect 264029 92085 264063 92113
rect 264091 92085 269379 92113
rect 269407 92085 269441 92113
rect 269469 92085 279237 92113
rect 279265 92085 279299 92113
rect 279327 92085 279361 92113
rect 279389 92085 279423 92113
rect 279451 92085 284739 92113
rect 284767 92085 284801 92113
rect 284829 92085 294597 92113
rect 294625 92085 294659 92113
rect 294687 92085 294721 92113
rect 294749 92085 294783 92113
rect 294811 92085 298248 92113
rect 298276 92085 298310 92113
rect 298338 92085 298372 92113
rect 298400 92085 298434 92113
rect 298462 92085 298990 92113
rect -958 92051 298990 92085
rect -958 92023 -430 92051
rect -402 92023 -368 92051
rect -340 92023 -306 92051
rect -278 92023 -244 92051
rect -216 92023 2757 92051
rect 2785 92023 2819 92051
rect 2847 92023 2881 92051
rect 2909 92023 2943 92051
rect 2971 92023 8259 92051
rect 8287 92023 8321 92051
rect 8349 92023 18117 92051
rect 18145 92023 18179 92051
rect 18207 92023 18241 92051
rect 18269 92023 18303 92051
rect 18331 92023 23619 92051
rect 23647 92023 23681 92051
rect 23709 92023 33477 92051
rect 33505 92023 33539 92051
rect 33567 92023 33601 92051
rect 33629 92023 33663 92051
rect 33691 92023 38979 92051
rect 39007 92023 39041 92051
rect 39069 92023 48837 92051
rect 48865 92023 48899 92051
rect 48927 92023 48961 92051
rect 48989 92023 49023 92051
rect 49051 92023 54339 92051
rect 54367 92023 54401 92051
rect 54429 92023 64197 92051
rect 64225 92023 64259 92051
rect 64287 92023 64321 92051
rect 64349 92023 64383 92051
rect 64411 92023 69699 92051
rect 69727 92023 69761 92051
rect 69789 92023 79557 92051
rect 79585 92023 79619 92051
rect 79647 92023 79681 92051
rect 79709 92023 79743 92051
rect 79771 92023 85059 92051
rect 85087 92023 85121 92051
rect 85149 92023 94917 92051
rect 94945 92023 94979 92051
rect 95007 92023 95041 92051
rect 95069 92023 95103 92051
rect 95131 92023 100419 92051
rect 100447 92023 100481 92051
rect 100509 92023 110277 92051
rect 110305 92023 110339 92051
rect 110367 92023 110401 92051
rect 110429 92023 110463 92051
rect 110491 92023 115779 92051
rect 115807 92023 115841 92051
rect 115869 92023 125637 92051
rect 125665 92023 125699 92051
rect 125727 92023 125761 92051
rect 125789 92023 125823 92051
rect 125851 92023 131139 92051
rect 131167 92023 131201 92051
rect 131229 92023 140997 92051
rect 141025 92023 141059 92051
rect 141087 92023 141121 92051
rect 141149 92023 141183 92051
rect 141211 92023 146499 92051
rect 146527 92023 146561 92051
rect 146589 92023 156357 92051
rect 156385 92023 156419 92051
rect 156447 92023 156481 92051
rect 156509 92023 156543 92051
rect 156571 92023 161859 92051
rect 161887 92023 161921 92051
rect 161949 92023 171717 92051
rect 171745 92023 171779 92051
rect 171807 92023 171841 92051
rect 171869 92023 171903 92051
rect 171931 92023 177219 92051
rect 177247 92023 177281 92051
rect 177309 92023 187077 92051
rect 187105 92023 187139 92051
rect 187167 92023 187201 92051
rect 187229 92023 187263 92051
rect 187291 92023 192579 92051
rect 192607 92023 192641 92051
rect 192669 92023 202437 92051
rect 202465 92023 202499 92051
rect 202527 92023 202561 92051
rect 202589 92023 202623 92051
rect 202651 92023 207939 92051
rect 207967 92023 208001 92051
rect 208029 92023 217797 92051
rect 217825 92023 217859 92051
rect 217887 92023 217921 92051
rect 217949 92023 217983 92051
rect 218011 92023 223299 92051
rect 223327 92023 223361 92051
rect 223389 92023 233157 92051
rect 233185 92023 233219 92051
rect 233247 92023 233281 92051
rect 233309 92023 233343 92051
rect 233371 92023 238659 92051
rect 238687 92023 238721 92051
rect 238749 92023 248517 92051
rect 248545 92023 248579 92051
rect 248607 92023 248641 92051
rect 248669 92023 248703 92051
rect 248731 92023 254019 92051
rect 254047 92023 254081 92051
rect 254109 92023 263877 92051
rect 263905 92023 263939 92051
rect 263967 92023 264001 92051
rect 264029 92023 264063 92051
rect 264091 92023 269379 92051
rect 269407 92023 269441 92051
rect 269469 92023 279237 92051
rect 279265 92023 279299 92051
rect 279327 92023 279361 92051
rect 279389 92023 279423 92051
rect 279451 92023 284739 92051
rect 284767 92023 284801 92051
rect 284829 92023 294597 92051
rect 294625 92023 294659 92051
rect 294687 92023 294721 92051
rect 294749 92023 294783 92051
rect 294811 92023 298248 92051
rect 298276 92023 298310 92051
rect 298338 92023 298372 92051
rect 298400 92023 298434 92051
rect 298462 92023 298990 92051
rect -958 91989 298990 92023
rect -958 91961 -430 91989
rect -402 91961 -368 91989
rect -340 91961 -306 91989
rect -278 91961 -244 91989
rect -216 91961 2757 91989
rect 2785 91961 2819 91989
rect 2847 91961 2881 91989
rect 2909 91961 2943 91989
rect 2971 91961 8259 91989
rect 8287 91961 8321 91989
rect 8349 91961 18117 91989
rect 18145 91961 18179 91989
rect 18207 91961 18241 91989
rect 18269 91961 18303 91989
rect 18331 91961 23619 91989
rect 23647 91961 23681 91989
rect 23709 91961 33477 91989
rect 33505 91961 33539 91989
rect 33567 91961 33601 91989
rect 33629 91961 33663 91989
rect 33691 91961 38979 91989
rect 39007 91961 39041 91989
rect 39069 91961 48837 91989
rect 48865 91961 48899 91989
rect 48927 91961 48961 91989
rect 48989 91961 49023 91989
rect 49051 91961 54339 91989
rect 54367 91961 54401 91989
rect 54429 91961 64197 91989
rect 64225 91961 64259 91989
rect 64287 91961 64321 91989
rect 64349 91961 64383 91989
rect 64411 91961 69699 91989
rect 69727 91961 69761 91989
rect 69789 91961 79557 91989
rect 79585 91961 79619 91989
rect 79647 91961 79681 91989
rect 79709 91961 79743 91989
rect 79771 91961 85059 91989
rect 85087 91961 85121 91989
rect 85149 91961 94917 91989
rect 94945 91961 94979 91989
rect 95007 91961 95041 91989
rect 95069 91961 95103 91989
rect 95131 91961 100419 91989
rect 100447 91961 100481 91989
rect 100509 91961 110277 91989
rect 110305 91961 110339 91989
rect 110367 91961 110401 91989
rect 110429 91961 110463 91989
rect 110491 91961 115779 91989
rect 115807 91961 115841 91989
rect 115869 91961 125637 91989
rect 125665 91961 125699 91989
rect 125727 91961 125761 91989
rect 125789 91961 125823 91989
rect 125851 91961 131139 91989
rect 131167 91961 131201 91989
rect 131229 91961 140997 91989
rect 141025 91961 141059 91989
rect 141087 91961 141121 91989
rect 141149 91961 141183 91989
rect 141211 91961 146499 91989
rect 146527 91961 146561 91989
rect 146589 91961 156357 91989
rect 156385 91961 156419 91989
rect 156447 91961 156481 91989
rect 156509 91961 156543 91989
rect 156571 91961 161859 91989
rect 161887 91961 161921 91989
rect 161949 91961 171717 91989
rect 171745 91961 171779 91989
rect 171807 91961 171841 91989
rect 171869 91961 171903 91989
rect 171931 91961 177219 91989
rect 177247 91961 177281 91989
rect 177309 91961 187077 91989
rect 187105 91961 187139 91989
rect 187167 91961 187201 91989
rect 187229 91961 187263 91989
rect 187291 91961 192579 91989
rect 192607 91961 192641 91989
rect 192669 91961 202437 91989
rect 202465 91961 202499 91989
rect 202527 91961 202561 91989
rect 202589 91961 202623 91989
rect 202651 91961 207939 91989
rect 207967 91961 208001 91989
rect 208029 91961 217797 91989
rect 217825 91961 217859 91989
rect 217887 91961 217921 91989
rect 217949 91961 217983 91989
rect 218011 91961 223299 91989
rect 223327 91961 223361 91989
rect 223389 91961 233157 91989
rect 233185 91961 233219 91989
rect 233247 91961 233281 91989
rect 233309 91961 233343 91989
rect 233371 91961 238659 91989
rect 238687 91961 238721 91989
rect 238749 91961 248517 91989
rect 248545 91961 248579 91989
rect 248607 91961 248641 91989
rect 248669 91961 248703 91989
rect 248731 91961 254019 91989
rect 254047 91961 254081 91989
rect 254109 91961 263877 91989
rect 263905 91961 263939 91989
rect 263967 91961 264001 91989
rect 264029 91961 264063 91989
rect 264091 91961 269379 91989
rect 269407 91961 269441 91989
rect 269469 91961 279237 91989
rect 279265 91961 279299 91989
rect 279327 91961 279361 91989
rect 279389 91961 279423 91989
rect 279451 91961 284739 91989
rect 284767 91961 284801 91989
rect 284829 91961 294597 91989
rect 294625 91961 294659 91989
rect 294687 91961 294721 91989
rect 294749 91961 294783 91989
rect 294811 91961 298248 91989
rect 298276 91961 298310 91989
rect 298338 91961 298372 91989
rect 298400 91961 298434 91989
rect 298462 91961 298990 91989
rect -958 91913 298990 91961
rect -958 86175 298990 86223
rect -958 86147 -910 86175
rect -882 86147 -848 86175
rect -820 86147 -786 86175
rect -758 86147 -724 86175
rect -696 86147 4617 86175
rect 4645 86147 4679 86175
rect 4707 86147 4741 86175
rect 4769 86147 4803 86175
rect 4831 86147 15939 86175
rect 15967 86147 16001 86175
rect 16029 86147 19977 86175
rect 20005 86147 20039 86175
rect 20067 86147 20101 86175
rect 20129 86147 20163 86175
rect 20191 86147 31299 86175
rect 31327 86147 31361 86175
rect 31389 86147 35337 86175
rect 35365 86147 35399 86175
rect 35427 86147 35461 86175
rect 35489 86147 35523 86175
rect 35551 86147 46659 86175
rect 46687 86147 46721 86175
rect 46749 86147 50697 86175
rect 50725 86147 50759 86175
rect 50787 86147 50821 86175
rect 50849 86147 50883 86175
rect 50911 86147 62019 86175
rect 62047 86147 62081 86175
rect 62109 86147 66057 86175
rect 66085 86147 66119 86175
rect 66147 86147 66181 86175
rect 66209 86147 66243 86175
rect 66271 86147 77379 86175
rect 77407 86147 77441 86175
rect 77469 86147 81417 86175
rect 81445 86147 81479 86175
rect 81507 86147 81541 86175
rect 81569 86147 81603 86175
rect 81631 86147 92739 86175
rect 92767 86147 92801 86175
rect 92829 86147 96777 86175
rect 96805 86147 96839 86175
rect 96867 86147 96901 86175
rect 96929 86147 96963 86175
rect 96991 86147 108099 86175
rect 108127 86147 108161 86175
rect 108189 86147 112137 86175
rect 112165 86147 112199 86175
rect 112227 86147 112261 86175
rect 112289 86147 112323 86175
rect 112351 86147 123459 86175
rect 123487 86147 123521 86175
rect 123549 86147 127497 86175
rect 127525 86147 127559 86175
rect 127587 86147 127621 86175
rect 127649 86147 127683 86175
rect 127711 86147 138819 86175
rect 138847 86147 138881 86175
rect 138909 86147 142857 86175
rect 142885 86147 142919 86175
rect 142947 86147 142981 86175
rect 143009 86147 143043 86175
rect 143071 86147 154179 86175
rect 154207 86147 154241 86175
rect 154269 86147 158217 86175
rect 158245 86147 158279 86175
rect 158307 86147 158341 86175
rect 158369 86147 158403 86175
rect 158431 86147 169539 86175
rect 169567 86147 169601 86175
rect 169629 86147 173577 86175
rect 173605 86147 173639 86175
rect 173667 86147 173701 86175
rect 173729 86147 173763 86175
rect 173791 86147 184899 86175
rect 184927 86147 184961 86175
rect 184989 86147 188937 86175
rect 188965 86147 188999 86175
rect 189027 86147 189061 86175
rect 189089 86147 189123 86175
rect 189151 86147 200259 86175
rect 200287 86147 200321 86175
rect 200349 86147 204297 86175
rect 204325 86147 204359 86175
rect 204387 86147 204421 86175
rect 204449 86147 204483 86175
rect 204511 86147 215619 86175
rect 215647 86147 215681 86175
rect 215709 86147 219657 86175
rect 219685 86147 219719 86175
rect 219747 86147 219781 86175
rect 219809 86147 219843 86175
rect 219871 86147 230979 86175
rect 231007 86147 231041 86175
rect 231069 86147 235017 86175
rect 235045 86147 235079 86175
rect 235107 86147 235141 86175
rect 235169 86147 235203 86175
rect 235231 86147 246339 86175
rect 246367 86147 246401 86175
rect 246429 86147 250377 86175
rect 250405 86147 250439 86175
rect 250467 86147 250501 86175
rect 250529 86147 250563 86175
rect 250591 86147 261699 86175
rect 261727 86147 261761 86175
rect 261789 86147 265737 86175
rect 265765 86147 265799 86175
rect 265827 86147 265861 86175
rect 265889 86147 265923 86175
rect 265951 86147 277059 86175
rect 277087 86147 277121 86175
rect 277149 86147 281097 86175
rect 281125 86147 281159 86175
rect 281187 86147 281221 86175
rect 281249 86147 281283 86175
rect 281311 86147 296457 86175
rect 296485 86147 296519 86175
rect 296547 86147 296581 86175
rect 296609 86147 296643 86175
rect 296671 86147 298728 86175
rect 298756 86147 298790 86175
rect 298818 86147 298852 86175
rect 298880 86147 298914 86175
rect 298942 86147 298990 86175
rect -958 86113 298990 86147
rect -958 86085 -910 86113
rect -882 86085 -848 86113
rect -820 86085 -786 86113
rect -758 86085 -724 86113
rect -696 86085 4617 86113
rect 4645 86085 4679 86113
rect 4707 86085 4741 86113
rect 4769 86085 4803 86113
rect 4831 86085 15939 86113
rect 15967 86085 16001 86113
rect 16029 86085 19977 86113
rect 20005 86085 20039 86113
rect 20067 86085 20101 86113
rect 20129 86085 20163 86113
rect 20191 86085 31299 86113
rect 31327 86085 31361 86113
rect 31389 86085 35337 86113
rect 35365 86085 35399 86113
rect 35427 86085 35461 86113
rect 35489 86085 35523 86113
rect 35551 86085 46659 86113
rect 46687 86085 46721 86113
rect 46749 86085 50697 86113
rect 50725 86085 50759 86113
rect 50787 86085 50821 86113
rect 50849 86085 50883 86113
rect 50911 86085 62019 86113
rect 62047 86085 62081 86113
rect 62109 86085 66057 86113
rect 66085 86085 66119 86113
rect 66147 86085 66181 86113
rect 66209 86085 66243 86113
rect 66271 86085 77379 86113
rect 77407 86085 77441 86113
rect 77469 86085 81417 86113
rect 81445 86085 81479 86113
rect 81507 86085 81541 86113
rect 81569 86085 81603 86113
rect 81631 86085 92739 86113
rect 92767 86085 92801 86113
rect 92829 86085 96777 86113
rect 96805 86085 96839 86113
rect 96867 86085 96901 86113
rect 96929 86085 96963 86113
rect 96991 86085 108099 86113
rect 108127 86085 108161 86113
rect 108189 86085 112137 86113
rect 112165 86085 112199 86113
rect 112227 86085 112261 86113
rect 112289 86085 112323 86113
rect 112351 86085 123459 86113
rect 123487 86085 123521 86113
rect 123549 86085 127497 86113
rect 127525 86085 127559 86113
rect 127587 86085 127621 86113
rect 127649 86085 127683 86113
rect 127711 86085 138819 86113
rect 138847 86085 138881 86113
rect 138909 86085 142857 86113
rect 142885 86085 142919 86113
rect 142947 86085 142981 86113
rect 143009 86085 143043 86113
rect 143071 86085 154179 86113
rect 154207 86085 154241 86113
rect 154269 86085 158217 86113
rect 158245 86085 158279 86113
rect 158307 86085 158341 86113
rect 158369 86085 158403 86113
rect 158431 86085 169539 86113
rect 169567 86085 169601 86113
rect 169629 86085 173577 86113
rect 173605 86085 173639 86113
rect 173667 86085 173701 86113
rect 173729 86085 173763 86113
rect 173791 86085 184899 86113
rect 184927 86085 184961 86113
rect 184989 86085 188937 86113
rect 188965 86085 188999 86113
rect 189027 86085 189061 86113
rect 189089 86085 189123 86113
rect 189151 86085 200259 86113
rect 200287 86085 200321 86113
rect 200349 86085 204297 86113
rect 204325 86085 204359 86113
rect 204387 86085 204421 86113
rect 204449 86085 204483 86113
rect 204511 86085 215619 86113
rect 215647 86085 215681 86113
rect 215709 86085 219657 86113
rect 219685 86085 219719 86113
rect 219747 86085 219781 86113
rect 219809 86085 219843 86113
rect 219871 86085 230979 86113
rect 231007 86085 231041 86113
rect 231069 86085 235017 86113
rect 235045 86085 235079 86113
rect 235107 86085 235141 86113
rect 235169 86085 235203 86113
rect 235231 86085 246339 86113
rect 246367 86085 246401 86113
rect 246429 86085 250377 86113
rect 250405 86085 250439 86113
rect 250467 86085 250501 86113
rect 250529 86085 250563 86113
rect 250591 86085 261699 86113
rect 261727 86085 261761 86113
rect 261789 86085 265737 86113
rect 265765 86085 265799 86113
rect 265827 86085 265861 86113
rect 265889 86085 265923 86113
rect 265951 86085 277059 86113
rect 277087 86085 277121 86113
rect 277149 86085 281097 86113
rect 281125 86085 281159 86113
rect 281187 86085 281221 86113
rect 281249 86085 281283 86113
rect 281311 86085 296457 86113
rect 296485 86085 296519 86113
rect 296547 86085 296581 86113
rect 296609 86085 296643 86113
rect 296671 86085 298728 86113
rect 298756 86085 298790 86113
rect 298818 86085 298852 86113
rect 298880 86085 298914 86113
rect 298942 86085 298990 86113
rect -958 86051 298990 86085
rect -958 86023 -910 86051
rect -882 86023 -848 86051
rect -820 86023 -786 86051
rect -758 86023 -724 86051
rect -696 86023 4617 86051
rect 4645 86023 4679 86051
rect 4707 86023 4741 86051
rect 4769 86023 4803 86051
rect 4831 86023 15939 86051
rect 15967 86023 16001 86051
rect 16029 86023 19977 86051
rect 20005 86023 20039 86051
rect 20067 86023 20101 86051
rect 20129 86023 20163 86051
rect 20191 86023 31299 86051
rect 31327 86023 31361 86051
rect 31389 86023 35337 86051
rect 35365 86023 35399 86051
rect 35427 86023 35461 86051
rect 35489 86023 35523 86051
rect 35551 86023 46659 86051
rect 46687 86023 46721 86051
rect 46749 86023 50697 86051
rect 50725 86023 50759 86051
rect 50787 86023 50821 86051
rect 50849 86023 50883 86051
rect 50911 86023 62019 86051
rect 62047 86023 62081 86051
rect 62109 86023 66057 86051
rect 66085 86023 66119 86051
rect 66147 86023 66181 86051
rect 66209 86023 66243 86051
rect 66271 86023 77379 86051
rect 77407 86023 77441 86051
rect 77469 86023 81417 86051
rect 81445 86023 81479 86051
rect 81507 86023 81541 86051
rect 81569 86023 81603 86051
rect 81631 86023 92739 86051
rect 92767 86023 92801 86051
rect 92829 86023 96777 86051
rect 96805 86023 96839 86051
rect 96867 86023 96901 86051
rect 96929 86023 96963 86051
rect 96991 86023 108099 86051
rect 108127 86023 108161 86051
rect 108189 86023 112137 86051
rect 112165 86023 112199 86051
rect 112227 86023 112261 86051
rect 112289 86023 112323 86051
rect 112351 86023 123459 86051
rect 123487 86023 123521 86051
rect 123549 86023 127497 86051
rect 127525 86023 127559 86051
rect 127587 86023 127621 86051
rect 127649 86023 127683 86051
rect 127711 86023 138819 86051
rect 138847 86023 138881 86051
rect 138909 86023 142857 86051
rect 142885 86023 142919 86051
rect 142947 86023 142981 86051
rect 143009 86023 143043 86051
rect 143071 86023 154179 86051
rect 154207 86023 154241 86051
rect 154269 86023 158217 86051
rect 158245 86023 158279 86051
rect 158307 86023 158341 86051
rect 158369 86023 158403 86051
rect 158431 86023 169539 86051
rect 169567 86023 169601 86051
rect 169629 86023 173577 86051
rect 173605 86023 173639 86051
rect 173667 86023 173701 86051
rect 173729 86023 173763 86051
rect 173791 86023 184899 86051
rect 184927 86023 184961 86051
rect 184989 86023 188937 86051
rect 188965 86023 188999 86051
rect 189027 86023 189061 86051
rect 189089 86023 189123 86051
rect 189151 86023 200259 86051
rect 200287 86023 200321 86051
rect 200349 86023 204297 86051
rect 204325 86023 204359 86051
rect 204387 86023 204421 86051
rect 204449 86023 204483 86051
rect 204511 86023 215619 86051
rect 215647 86023 215681 86051
rect 215709 86023 219657 86051
rect 219685 86023 219719 86051
rect 219747 86023 219781 86051
rect 219809 86023 219843 86051
rect 219871 86023 230979 86051
rect 231007 86023 231041 86051
rect 231069 86023 235017 86051
rect 235045 86023 235079 86051
rect 235107 86023 235141 86051
rect 235169 86023 235203 86051
rect 235231 86023 246339 86051
rect 246367 86023 246401 86051
rect 246429 86023 250377 86051
rect 250405 86023 250439 86051
rect 250467 86023 250501 86051
rect 250529 86023 250563 86051
rect 250591 86023 261699 86051
rect 261727 86023 261761 86051
rect 261789 86023 265737 86051
rect 265765 86023 265799 86051
rect 265827 86023 265861 86051
rect 265889 86023 265923 86051
rect 265951 86023 277059 86051
rect 277087 86023 277121 86051
rect 277149 86023 281097 86051
rect 281125 86023 281159 86051
rect 281187 86023 281221 86051
rect 281249 86023 281283 86051
rect 281311 86023 296457 86051
rect 296485 86023 296519 86051
rect 296547 86023 296581 86051
rect 296609 86023 296643 86051
rect 296671 86023 298728 86051
rect 298756 86023 298790 86051
rect 298818 86023 298852 86051
rect 298880 86023 298914 86051
rect 298942 86023 298990 86051
rect -958 85989 298990 86023
rect -958 85961 -910 85989
rect -882 85961 -848 85989
rect -820 85961 -786 85989
rect -758 85961 -724 85989
rect -696 85961 4617 85989
rect 4645 85961 4679 85989
rect 4707 85961 4741 85989
rect 4769 85961 4803 85989
rect 4831 85961 15939 85989
rect 15967 85961 16001 85989
rect 16029 85961 19977 85989
rect 20005 85961 20039 85989
rect 20067 85961 20101 85989
rect 20129 85961 20163 85989
rect 20191 85961 31299 85989
rect 31327 85961 31361 85989
rect 31389 85961 35337 85989
rect 35365 85961 35399 85989
rect 35427 85961 35461 85989
rect 35489 85961 35523 85989
rect 35551 85961 46659 85989
rect 46687 85961 46721 85989
rect 46749 85961 50697 85989
rect 50725 85961 50759 85989
rect 50787 85961 50821 85989
rect 50849 85961 50883 85989
rect 50911 85961 62019 85989
rect 62047 85961 62081 85989
rect 62109 85961 66057 85989
rect 66085 85961 66119 85989
rect 66147 85961 66181 85989
rect 66209 85961 66243 85989
rect 66271 85961 77379 85989
rect 77407 85961 77441 85989
rect 77469 85961 81417 85989
rect 81445 85961 81479 85989
rect 81507 85961 81541 85989
rect 81569 85961 81603 85989
rect 81631 85961 92739 85989
rect 92767 85961 92801 85989
rect 92829 85961 96777 85989
rect 96805 85961 96839 85989
rect 96867 85961 96901 85989
rect 96929 85961 96963 85989
rect 96991 85961 108099 85989
rect 108127 85961 108161 85989
rect 108189 85961 112137 85989
rect 112165 85961 112199 85989
rect 112227 85961 112261 85989
rect 112289 85961 112323 85989
rect 112351 85961 123459 85989
rect 123487 85961 123521 85989
rect 123549 85961 127497 85989
rect 127525 85961 127559 85989
rect 127587 85961 127621 85989
rect 127649 85961 127683 85989
rect 127711 85961 138819 85989
rect 138847 85961 138881 85989
rect 138909 85961 142857 85989
rect 142885 85961 142919 85989
rect 142947 85961 142981 85989
rect 143009 85961 143043 85989
rect 143071 85961 154179 85989
rect 154207 85961 154241 85989
rect 154269 85961 158217 85989
rect 158245 85961 158279 85989
rect 158307 85961 158341 85989
rect 158369 85961 158403 85989
rect 158431 85961 169539 85989
rect 169567 85961 169601 85989
rect 169629 85961 173577 85989
rect 173605 85961 173639 85989
rect 173667 85961 173701 85989
rect 173729 85961 173763 85989
rect 173791 85961 184899 85989
rect 184927 85961 184961 85989
rect 184989 85961 188937 85989
rect 188965 85961 188999 85989
rect 189027 85961 189061 85989
rect 189089 85961 189123 85989
rect 189151 85961 200259 85989
rect 200287 85961 200321 85989
rect 200349 85961 204297 85989
rect 204325 85961 204359 85989
rect 204387 85961 204421 85989
rect 204449 85961 204483 85989
rect 204511 85961 215619 85989
rect 215647 85961 215681 85989
rect 215709 85961 219657 85989
rect 219685 85961 219719 85989
rect 219747 85961 219781 85989
rect 219809 85961 219843 85989
rect 219871 85961 230979 85989
rect 231007 85961 231041 85989
rect 231069 85961 235017 85989
rect 235045 85961 235079 85989
rect 235107 85961 235141 85989
rect 235169 85961 235203 85989
rect 235231 85961 246339 85989
rect 246367 85961 246401 85989
rect 246429 85961 250377 85989
rect 250405 85961 250439 85989
rect 250467 85961 250501 85989
rect 250529 85961 250563 85989
rect 250591 85961 261699 85989
rect 261727 85961 261761 85989
rect 261789 85961 265737 85989
rect 265765 85961 265799 85989
rect 265827 85961 265861 85989
rect 265889 85961 265923 85989
rect 265951 85961 277059 85989
rect 277087 85961 277121 85989
rect 277149 85961 281097 85989
rect 281125 85961 281159 85989
rect 281187 85961 281221 85989
rect 281249 85961 281283 85989
rect 281311 85961 296457 85989
rect 296485 85961 296519 85989
rect 296547 85961 296581 85989
rect 296609 85961 296643 85989
rect 296671 85961 298728 85989
rect 298756 85961 298790 85989
rect 298818 85961 298852 85989
rect 298880 85961 298914 85989
rect 298942 85961 298990 85989
rect -958 85913 298990 85961
rect -958 83175 298990 83223
rect -958 83147 -430 83175
rect -402 83147 -368 83175
rect -340 83147 -306 83175
rect -278 83147 -244 83175
rect -216 83147 2757 83175
rect 2785 83147 2819 83175
rect 2847 83147 2881 83175
rect 2909 83147 2943 83175
rect 2971 83147 8259 83175
rect 8287 83147 8321 83175
rect 8349 83147 18117 83175
rect 18145 83147 18179 83175
rect 18207 83147 18241 83175
rect 18269 83147 18303 83175
rect 18331 83147 23619 83175
rect 23647 83147 23681 83175
rect 23709 83147 33477 83175
rect 33505 83147 33539 83175
rect 33567 83147 33601 83175
rect 33629 83147 33663 83175
rect 33691 83147 38979 83175
rect 39007 83147 39041 83175
rect 39069 83147 48837 83175
rect 48865 83147 48899 83175
rect 48927 83147 48961 83175
rect 48989 83147 49023 83175
rect 49051 83147 54339 83175
rect 54367 83147 54401 83175
rect 54429 83147 64197 83175
rect 64225 83147 64259 83175
rect 64287 83147 64321 83175
rect 64349 83147 64383 83175
rect 64411 83147 69699 83175
rect 69727 83147 69761 83175
rect 69789 83147 79557 83175
rect 79585 83147 79619 83175
rect 79647 83147 79681 83175
rect 79709 83147 79743 83175
rect 79771 83147 85059 83175
rect 85087 83147 85121 83175
rect 85149 83147 94917 83175
rect 94945 83147 94979 83175
rect 95007 83147 95041 83175
rect 95069 83147 95103 83175
rect 95131 83147 100419 83175
rect 100447 83147 100481 83175
rect 100509 83147 110277 83175
rect 110305 83147 110339 83175
rect 110367 83147 110401 83175
rect 110429 83147 110463 83175
rect 110491 83147 115779 83175
rect 115807 83147 115841 83175
rect 115869 83147 125637 83175
rect 125665 83147 125699 83175
rect 125727 83147 125761 83175
rect 125789 83147 125823 83175
rect 125851 83147 131139 83175
rect 131167 83147 131201 83175
rect 131229 83147 140997 83175
rect 141025 83147 141059 83175
rect 141087 83147 141121 83175
rect 141149 83147 141183 83175
rect 141211 83147 146499 83175
rect 146527 83147 146561 83175
rect 146589 83147 156357 83175
rect 156385 83147 156419 83175
rect 156447 83147 156481 83175
rect 156509 83147 156543 83175
rect 156571 83147 161859 83175
rect 161887 83147 161921 83175
rect 161949 83147 171717 83175
rect 171745 83147 171779 83175
rect 171807 83147 171841 83175
rect 171869 83147 171903 83175
rect 171931 83147 177219 83175
rect 177247 83147 177281 83175
rect 177309 83147 187077 83175
rect 187105 83147 187139 83175
rect 187167 83147 187201 83175
rect 187229 83147 187263 83175
rect 187291 83147 192579 83175
rect 192607 83147 192641 83175
rect 192669 83147 202437 83175
rect 202465 83147 202499 83175
rect 202527 83147 202561 83175
rect 202589 83147 202623 83175
rect 202651 83147 207939 83175
rect 207967 83147 208001 83175
rect 208029 83147 217797 83175
rect 217825 83147 217859 83175
rect 217887 83147 217921 83175
rect 217949 83147 217983 83175
rect 218011 83147 223299 83175
rect 223327 83147 223361 83175
rect 223389 83147 233157 83175
rect 233185 83147 233219 83175
rect 233247 83147 233281 83175
rect 233309 83147 233343 83175
rect 233371 83147 238659 83175
rect 238687 83147 238721 83175
rect 238749 83147 248517 83175
rect 248545 83147 248579 83175
rect 248607 83147 248641 83175
rect 248669 83147 248703 83175
rect 248731 83147 254019 83175
rect 254047 83147 254081 83175
rect 254109 83147 263877 83175
rect 263905 83147 263939 83175
rect 263967 83147 264001 83175
rect 264029 83147 264063 83175
rect 264091 83147 269379 83175
rect 269407 83147 269441 83175
rect 269469 83147 279237 83175
rect 279265 83147 279299 83175
rect 279327 83147 279361 83175
rect 279389 83147 279423 83175
rect 279451 83147 284739 83175
rect 284767 83147 284801 83175
rect 284829 83147 294597 83175
rect 294625 83147 294659 83175
rect 294687 83147 294721 83175
rect 294749 83147 294783 83175
rect 294811 83147 298248 83175
rect 298276 83147 298310 83175
rect 298338 83147 298372 83175
rect 298400 83147 298434 83175
rect 298462 83147 298990 83175
rect -958 83113 298990 83147
rect -958 83085 -430 83113
rect -402 83085 -368 83113
rect -340 83085 -306 83113
rect -278 83085 -244 83113
rect -216 83085 2757 83113
rect 2785 83085 2819 83113
rect 2847 83085 2881 83113
rect 2909 83085 2943 83113
rect 2971 83085 8259 83113
rect 8287 83085 8321 83113
rect 8349 83085 18117 83113
rect 18145 83085 18179 83113
rect 18207 83085 18241 83113
rect 18269 83085 18303 83113
rect 18331 83085 23619 83113
rect 23647 83085 23681 83113
rect 23709 83085 33477 83113
rect 33505 83085 33539 83113
rect 33567 83085 33601 83113
rect 33629 83085 33663 83113
rect 33691 83085 38979 83113
rect 39007 83085 39041 83113
rect 39069 83085 48837 83113
rect 48865 83085 48899 83113
rect 48927 83085 48961 83113
rect 48989 83085 49023 83113
rect 49051 83085 54339 83113
rect 54367 83085 54401 83113
rect 54429 83085 64197 83113
rect 64225 83085 64259 83113
rect 64287 83085 64321 83113
rect 64349 83085 64383 83113
rect 64411 83085 69699 83113
rect 69727 83085 69761 83113
rect 69789 83085 79557 83113
rect 79585 83085 79619 83113
rect 79647 83085 79681 83113
rect 79709 83085 79743 83113
rect 79771 83085 85059 83113
rect 85087 83085 85121 83113
rect 85149 83085 94917 83113
rect 94945 83085 94979 83113
rect 95007 83085 95041 83113
rect 95069 83085 95103 83113
rect 95131 83085 100419 83113
rect 100447 83085 100481 83113
rect 100509 83085 110277 83113
rect 110305 83085 110339 83113
rect 110367 83085 110401 83113
rect 110429 83085 110463 83113
rect 110491 83085 115779 83113
rect 115807 83085 115841 83113
rect 115869 83085 125637 83113
rect 125665 83085 125699 83113
rect 125727 83085 125761 83113
rect 125789 83085 125823 83113
rect 125851 83085 131139 83113
rect 131167 83085 131201 83113
rect 131229 83085 140997 83113
rect 141025 83085 141059 83113
rect 141087 83085 141121 83113
rect 141149 83085 141183 83113
rect 141211 83085 146499 83113
rect 146527 83085 146561 83113
rect 146589 83085 156357 83113
rect 156385 83085 156419 83113
rect 156447 83085 156481 83113
rect 156509 83085 156543 83113
rect 156571 83085 161859 83113
rect 161887 83085 161921 83113
rect 161949 83085 171717 83113
rect 171745 83085 171779 83113
rect 171807 83085 171841 83113
rect 171869 83085 171903 83113
rect 171931 83085 177219 83113
rect 177247 83085 177281 83113
rect 177309 83085 187077 83113
rect 187105 83085 187139 83113
rect 187167 83085 187201 83113
rect 187229 83085 187263 83113
rect 187291 83085 192579 83113
rect 192607 83085 192641 83113
rect 192669 83085 202437 83113
rect 202465 83085 202499 83113
rect 202527 83085 202561 83113
rect 202589 83085 202623 83113
rect 202651 83085 207939 83113
rect 207967 83085 208001 83113
rect 208029 83085 217797 83113
rect 217825 83085 217859 83113
rect 217887 83085 217921 83113
rect 217949 83085 217983 83113
rect 218011 83085 223299 83113
rect 223327 83085 223361 83113
rect 223389 83085 233157 83113
rect 233185 83085 233219 83113
rect 233247 83085 233281 83113
rect 233309 83085 233343 83113
rect 233371 83085 238659 83113
rect 238687 83085 238721 83113
rect 238749 83085 248517 83113
rect 248545 83085 248579 83113
rect 248607 83085 248641 83113
rect 248669 83085 248703 83113
rect 248731 83085 254019 83113
rect 254047 83085 254081 83113
rect 254109 83085 263877 83113
rect 263905 83085 263939 83113
rect 263967 83085 264001 83113
rect 264029 83085 264063 83113
rect 264091 83085 269379 83113
rect 269407 83085 269441 83113
rect 269469 83085 279237 83113
rect 279265 83085 279299 83113
rect 279327 83085 279361 83113
rect 279389 83085 279423 83113
rect 279451 83085 284739 83113
rect 284767 83085 284801 83113
rect 284829 83085 294597 83113
rect 294625 83085 294659 83113
rect 294687 83085 294721 83113
rect 294749 83085 294783 83113
rect 294811 83085 298248 83113
rect 298276 83085 298310 83113
rect 298338 83085 298372 83113
rect 298400 83085 298434 83113
rect 298462 83085 298990 83113
rect -958 83051 298990 83085
rect -958 83023 -430 83051
rect -402 83023 -368 83051
rect -340 83023 -306 83051
rect -278 83023 -244 83051
rect -216 83023 2757 83051
rect 2785 83023 2819 83051
rect 2847 83023 2881 83051
rect 2909 83023 2943 83051
rect 2971 83023 8259 83051
rect 8287 83023 8321 83051
rect 8349 83023 18117 83051
rect 18145 83023 18179 83051
rect 18207 83023 18241 83051
rect 18269 83023 18303 83051
rect 18331 83023 23619 83051
rect 23647 83023 23681 83051
rect 23709 83023 33477 83051
rect 33505 83023 33539 83051
rect 33567 83023 33601 83051
rect 33629 83023 33663 83051
rect 33691 83023 38979 83051
rect 39007 83023 39041 83051
rect 39069 83023 48837 83051
rect 48865 83023 48899 83051
rect 48927 83023 48961 83051
rect 48989 83023 49023 83051
rect 49051 83023 54339 83051
rect 54367 83023 54401 83051
rect 54429 83023 64197 83051
rect 64225 83023 64259 83051
rect 64287 83023 64321 83051
rect 64349 83023 64383 83051
rect 64411 83023 69699 83051
rect 69727 83023 69761 83051
rect 69789 83023 79557 83051
rect 79585 83023 79619 83051
rect 79647 83023 79681 83051
rect 79709 83023 79743 83051
rect 79771 83023 85059 83051
rect 85087 83023 85121 83051
rect 85149 83023 94917 83051
rect 94945 83023 94979 83051
rect 95007 83023 95041 83051
rect 95069 83023 95103 83051
rect 95131 83023 100419 83051
rect 100447 83023 100481 83051
rect 100509 83023 110277 83051
rect 110305 83023 110339 83051
rect 110367 83023 110401 83051
rect 110429 83023 110463 83051
rect 110491 83023 115779 83051
rect 115807 83023 115841 83051
rect 115869 83023 125637 83051
rect 125665 83023 125699 83051
rect 125727 83023 125761 83051
rect 125789 83023 125823 83051
rect 125851 83023 131139 83051
rect 131167 83023 131201 83051
rect 131229 83023 140997 83051
rect 141025 83023 141059 83051
rect 141087 83023 141121 83051
rect 141149 83023 141183 83051
rect 141211 83023 146499 83051
rect 146527 83023 146561 83051
rect 146589 83023 156357 83051
rect 156385 83023 156419 83051
rect 156447 83023 156481 83051
rect 156509 83023 156543 83051
rect 156571 83023 161859 83051
rect 161887 83023 161921 83051
rect 161949 83023 171717 83051
rect 171745 83023 171779 83051
rect 171807 83023 171841 83051
rect 171869 83023 171903 83051
rect 171931 83023 177219 83051
rect 177247 83023 177281 83051
rect 177309 83023 187077 83051
rect 187105 83023 187139 83051
rect 187167 83023 187201 83051
rect 187229 83023 187263 83051
rect 187291 83023 192579 83051
rect 192607 83023 192641 83051
rect 192669 83023 202437 83051
rect 202465 83023 202499 83051
rect 202527 83023 202561 83051
rect 202589 83023 202623 83051
rect 202651 83023 207939 83051
rect 207967 83023 208001 83051
rect 208029 83023 217797 83051
rect 217825 83023 217859 83051
rect 217887 83023 217921 83051
rect 217949 83023 217983 83051
rect 218011 83023 223299 83051
rect 223327 83023 223361 83051
rect 223389 83023 233157 83051
rect 233185 83023 233219 83051
rect 233247 83023 233281 83051
rect 233309 83023 233343 83051
rect 233371 83023 238659 83051
rect 238687 83023 238721 83051
rect 238749 83023 248517 83051
rect 248545 83023 248579 83051
rect 248607 83023 248641 83051
rect 248669 83023 248703 83051
rect 248731 83023 254019 83051
rect 254047 83023 254081 83051
rect 254109 83023 263877 83051
rect 263905 83023 263939 83051
rect 263967 83023 264001 83051
rect 264029 83023 264063 83051
rect 264091 83023 269379 83051
rect 269407 83023 269441 83051
rect 269469 83023 279237 83051
rect 279265 83023 279299 83051
rect 279327 83023 279361 83051
rect 279389 83023 279423 83051
rect 279451 83023 284739 83051
rect 284767 83023 284801 83051
rect 284829 83023 294597 83051
rect 294625 83023 294659 83051
rect 294687 83023 294721 83051
rect 294749 83023 294783 83051
rect 294811 83023 298248 83051
rect 298276 83023 298310 83051
rect 298338 83023 298372 83051
rect 298400 83023 298434 83051
rect 298462 83023 298990 83051
rect -958 82989 298990 83023
rect -958 82961 -430 82989
rect -402 82961 -368 82989
rect -340 82961 -306 82989
rect -278 82961 -244 82989
rect -216 82961 2757 82989
rect 2785 82961 2819 82989
rect 2847 82961 2881 82989
rect 2909 82961 2943 82989
rect 2971 82961 8259 82989
rect 8287 82961 8321 82989
rect 8349 82961 18117 82989
rect 18145 82961 18179 82989
rect 18207 82961 18241 82989
rect 18269 82961 18303 82989
rect 18331 82961 23619 82989
rect 23647 82961 23681 82989
rect 23709 82961 33477 82989
rect 33505 82961 33539 82989
rect 33567 82961 33601 82989
rect 33629 82961 33663 82989
rect 33691 82961 38979 82989
rect 39007 82961 39041 82989
rect 39069 82961 48837 82989
rect 48865 82961 48899 82989
rect 48927 82961 48961 82989
rect 48989 82961 49023 82989
rect 49051 82961 54339 82989
rect 54367 82961 54401 82989
rect 54429 82961 64197 82989
rect 64225 82961 64259 82989
rect 64287 82961 64321 82989
rect 64349 82961 64383 82989
rect 64411 82961 69699 82989
rect 69727 82961 69761 82989
rect 69789 82961 79557 82989
rect 79585 82961 79619 82989
rect 79647 82961 79681 82989
rect 79709 82961 79743 82989
rect 79771 82961 85059 82989
rect 85087 82961 85121 82989
rect 85149 82961 94917 82989
rect 94945 82961 94979 82989
rect 95007 82961 95041 82989
rect 95069 82961 95103 82989
rect 95131 82961 100419 82989
rect 100447 82961 100481 82989
rect 100509 82961 110277 82989
rect 110305 82961 110339 82989
rect 110367 82961 110401 82989
rect 110429 82961 110463 82989
rect 110491 82961 115779 82989
rect 115807 82961 115841 82989
rect 115869 82961 125637 82989
rect 125665 82961 125699 82989
rect 125727 82961 125761 82989
rect 125789 82961 125823 82989
rect 125851 82961 131139 82989
rect 131167 82961 131201 82989
rect 131229 82961 140997 82989
rect 141025 82961 141059 82989
rect 141087 82961 141121 82989
rect 141149 82961 141183 82989
rect 141211 82961 146499 82989
rect 146527 82961 146561 82989
rect 146589 82961 156357 82989
rect 156385 82961 156419 82989
rect 156447 82961 156481 82989
rect 156509 82961 156543 82989
rect 156571 82961 161859 82989
rect 161887 82961 161921 82989
rect 161949 82961 171717 82989
rect 171745 82961 171779 82989
rect 171807 82961 171841 82989
rect 171869 82961 171903 82989
rect 171931 82961 177219 82989
rect 177247 82961 177281 82989
rect 177309 82961 187077 82989
rect 187105 82961 187139 82989
rect 187167 82961 187201 82989
rect 187229 82961 187263 82989
rect 187291 82961 192579 82989
rect 192607 82961 192641 82989
rect 192669 82961 202437 82989
rect 202465 82961 202499 82989
rect 202527 82961 202561 82989
rect 202589 82961 202623 82989
rect 202651 82961 207939 82989
rect 207967 82961 208001 82989
rect 208029 82961 217797 82989
rect 217825 82961 217859 82989
rect 217887 82961 217921 82989
rect 217949 82961 217983 82989
rect 218011 82961 223299 82989
rect 223327 82961 223361 82989
rect 223389 82961 233157 82989
rect 233185 82961 233219 82989
rect 233247 82961 233281 82989
rect 233309 82961 233343 82989
rect 233371 82961 238659 82989
rect 238687 82961 238721 82989
rect 238749 82961 248517 82989
rect 248545 82961 248579 82989
rect 248607 82961 248641 82989
rect 248669 82961 248703 82989
rect 248731 82961 254019 82989
rect 254047 82961 254081 82989
rect 254109 82961 263877 82989
rect 263905 82961 263939 82989
rect 263967 82961 264001 82989
rect 264029 82961 264063 82989
rect 264091 82961 269379 82989
rect 269407 82961 269441 82989
rect 269469 82961 279237 82989
rect 279265 82961 279299 82989
rect 279327 82961 279361 82989
rect 279389 82961 279423 82989
rect 279451 82961 284739 82989
rect 284767 82961 284801 82989
rect 284829 82961 294597 82989
rect 294625 82961 294659 82989
rect 294687 82961 294721 82989
rect 294749 82961 294783 82989
rect 294811 82961 298248 82989
rect 298276 82961 298310 82989
rect 298338 82961 298372 82989
rect 298400 82961 298434 82989
rect 298462 82961 298990 82989
rect -958 82913 298990 82961
rect -958 77175 298990 77223
rect -958 77147 -910 77175
rect -882 77147 -848 77175
rect -820 77147 -786 77175
rect -758 77147 -724 77175
rect -696 77147 4617 77175
rect 4645 77147 4679 77175
rect 4707 77147 4741 77175
rect 4769 77147 4803 77175
rect 4831 77147 15939 77175
rect 15967 77147 16001 77175
rect 16029 77147 19977 77175
rect 20005 77147 20039 77175
rect 20067 77147 20101 77175
rect 20129 77147 20163 77175
rect 20191 77147 31299 77175
rect 31327 77147 31361 77175
rect 31389 77147 35337 77175
rect 35365 77147 35399 77175
rect 35427 77147 35461 77175
rect 35489 77147 35523 77175
rect 35551 77147 46659 77175
rect 46687 77147 46721 77175
rect 46749 77147 50697 77175
rect 50725 77147 50759 77175
rect 50787 77147 50821 77175
rect 50849 77147 50883 77175
rect 50911 77147 62019 77175
rect 62047 77147 62081 77175
rect 62109 77147 66057 77175
rect 66085 77147 66119 77175
rect 66147 77147 66181 77175
rect 66209 77147 66243 77175
rect 66271 77147 77379 77175
rect 77407 77147 77441 77175
rect 77469 77147 81417 77175
rect 81445 77147 81479 77175
rect 81507 77147 81541 77175
rect 81569 77147 81603 77175
rect 81631 77147 92739 77175
rect 92767 77147 92801 77175
rect 92829 77147 96777 77175
rect 96805 77147 96839 77175
rect 96867 77147 96901 77175
rect 96929 77147 96963 77175
rect 96991 77147 108099 77175
rect 108127 77147 108161 77175
rect 108189 77147 112137 77175
rect 112165 77147 112199 77175
rect 112227 77147 112261 77175
rect 112289 77147 112323 77175
rect 112351 77147 123459 77175
rect 123487 77147 123521 77175
rect 123549 77147 127497 77175
rect 127525 77147 127559 77175
rect 127587 77147 127621 77175
rect 127649 77147 127683 77175
rect 127711 77147 138819 77175
rect 138847 77147 138881 77175
rect 138909 77147 142857 77175
rect 142885 77147 142919 77175
rect 142947 77147 142981 77175
rect 143009 77147 143043 77175
rect 143071 77147 154179 77175
rect 154207 77147 154241 77175
rect 154269 77147 158217 77175
rect 158245 77147 158279 77175
rect 158307 77147 158341 77175
rect 158369 77147 158403 77175
rect 158431 77147 169539 77175
rect 169567 77147 169601 77175
rect 169629 77147 173577 77175
rect 173605 77147 173639 77175
rect 173667 77147 173701 77175
rect 173729 77147 173763 77175
rect 173791 77147 184899 77175
rect 184927 77147 184961 77175
rect 184989 77147 188937 77175
rect 188965 77147 188999 77175
rect 189027 77147 189061 77175
rect 189089 77147 189123 77175
rect 189151 77147 200259 77175
rect 200287 77147 200321 77175
rect 200349 77147 204297 77175
rect 204325 77147 204359 77175
rect 204387 77147 204421 77175
rect 204449 77147 204483 77175
rect 204511 77147 215619 77175
rect 215647 77147 215681 77175
rect 215709 77147 219657 77175
rect 219685 77147 219719 77175
rect 219747 77147 219781 77175
rect 219809 77147 219843 77175
rect 219871 77147 230979 77175
rect 231007 77147 231041 77175
rect 231069 77147 235017 77175
rect 235045 77147 235079 77175
rect 235107 77147 235141 77175
rect 235169 77147 235203 77175
rect 235231 77147 246339 77175
rect 246367 77147 246401 77175
rect 246429 77147 250377 77175
rect 250405 77147 250439 77175
rect 250467 77147 250501 77175
rect 250529 77147 250563 77175
rect 250591 77147 261699 77175
rect 261727 77147 261761 77175
rect 261789 77147 265737 77175
rect 265765 77147 265799 77175
rect 265827 77147 265861 77175
rect 265889 77147 265923 77175
rect 265951 77147 277059 77175
rect 277087 77147 277121 77175
rect 277149 77147 281097 77175
rect 281125 77147 281159 77175
rect 281187 77147 281221 77175
rect 281249 77147 281283 77175
rect 281311 77147 296457 77175
rect 296485 77147 296519 77175
rect 296547 77147 296581 77175
rect 296609 77147 296643 77175
rect 296671 77147 298728 77175
rect 298756 77147 298790 77175
rect 298818 77147 298852 77175
rect 298880 77147 298914 77175
rect 298942 77147 298990 77175
rect -958 77113 298990 77147
rect -958 77085 -910 77113
rect -882 77085 -848 77113
rect -820 77085 -786 77113
rect -758 77085 -724 77113
rect -696 77085 4617 77113
rect 4645 77085 4679 77113
rect 4707 77085 4741 77113
rect 4769 77085 4803 77113
rect 4831 77085 15939 77113
rect 15967 77085 16001 77113
rect 16029 77085 19977 77113
rect 20005 77085 20039 77113
rect 20067 77085 20101 77113
rect 20129 77085 20163 77113
rect 20191 77085 31299 77113
rect 31327 77085 31361 77113
rect 31389 77085 35337 77113
rect 35365 77085 35399 77113
rect 35427 77085 35461 77113
rect 35489 77085 35523 77113
rect 35551 77085 46659 77113
rect 46687 77085 46721 77113
rect 46749 77085 50697 77113
rect 50725 77085 50759 77113
rect 50787 77085 50821 77113
rect 50849 77085 50883 77113
rect 50911 77085 62019 77113
rect 62047 77085 62081 77113
rect 62109 77085 66057 77113
rect 66085 77085 66119 77113
rect 66147 77085 66181 77113
rect 66209 77085 66243 77113
rect 66271 77085 77379 77113
rect 77407 77085 77441 77113
rect 77469 77085 81417 77113
rect 81445 77085 81479 77113
rect 81507 77085 81541 77113
rect 81569 77085 81603 77113
rect 81631 77085 92739 77113
rect 92767 77085 92801 77113
rect 92829 77085 96777 77113
rect 96805 77085 96839 77113
rect 96867 77085 96901 77113
rect 96929 77085 96963 77113
rect 96991 77085 108099 77113
rect 108127 77085 108161 77113
rect 108189 77085 112137 77113
rect 112165 77085 112199 77113
rect 112227 77085 112261 77113
rect 112289 77085 112323 77113
rect 112351 77085 123459 77113
rect 123487 77085 123521 77113
rect 123549 77085 127497 77113
rect 127525 77085 127559 77113
rect 127587 77085 127621 77113
rect 127649 77085 127683 77113
rect 127711 77085 138819 77113
rect 138847 77085 138881 77113
rect 138909 77085 142857 77113
rect 142885 77085 142919 77113
rect 142947 77085 142981 77113
rect 143009 77085 143043 77113
rect 143071 77085 154179 77113
rect 154207 77085 154241 77113
rect 154269 77085 158217 77113
rect 158245 77085 158279 77113
rect 158307 77085 158341 77113
rect 158369 77085 158403 77113
rect 158431 77085 169539 77113
rect 169567 77085 169601 77113
rect 169629 77085 173577 77113
rect 173605 77085 173639 77113
rect 173667 77085 173701 77113
rect 173729 77085 173763 77113
rect 173791 77085 184899 77113
rect 184927 77085 184961 77113
rect 184989 77085 188937 77113
rect 188965 77085 188999 77113
rect 189027 77085 189061 77113
rect 189089 77085 189123 77113
rect 189151 77085 200259 77113
rect 200287 77085 200321 77113
rect 200349 77085 204297 77113
rect 204325 77085 204359 77113
rect 204387 77085 204421 77113
rect 204449 77085 204483 77113
rect 204511 77085 215619 77113
rect 215647 77085 215681 77113
rect 215709 77085 219657 77113
rect 219685 77085 219719 77113
rect 219747 77085 219781 77113
rect 219809 77085 219843 77113
rect 219871 77085 230979 77113
rect 231007 77085 231041 77113
rect 231069 77085 235017 77113
rect 235045 77085 235079 77113
rect 235107 77085 235141 77113
rect 235169 77085 235203 77113
rect 235231 77085 246339 77113
rect 246367 77085 246401 77113
rect 246429 77085 250377 77113
rect 250405 77085 250439 77113
rect 250467 77085 250501 77113
rect 250529 77085 250563 77113
rect 250591 77085 261699 77113
rect 261727 77085 261761 77113
rect 261789 77085 265737 77113
rect 265765 77085 265799 77113
rect 265827 77085 265861 77113
rect 265889 77085 265923 77113
rect 265951 77085 277059 77113
rect 277087 77085 277121 77113
rect 277149 77085 281097 77113
rect 281125 77085 281159 77113
rect 281187 77085 281221 77113
rect 281249 77085 281283 77113
rect 281311 77085 296457 77113
rect 296485 77085 296519 77113
rect 296547 77085 296581 77113
rect 296609 77085 296643 77113
rect 296671 77085 298728 77113
rect 298756 77085 298790 77113
rect 298818 77085 298852 77113
rect 298880 77085 298914 77113
rect 298942 77085 298990 77113
rect -958 77051 298990 77085
rect -958 77023 -910 77051
rect -882 77023 -848 77051
rect -820 77023 -786 77051
rect -758 77023 -724 77051
rect -696 77023 4617 77051
rect 4645 77023 4679 77051
rect 4707 77023 4741 77051
rect 4769 77023 4803 77051
rect 4831 77023 15939 77051
rect 15967 77023 16001 77051
rect 16029 77023 19977 77051
rect 20005 77023 20039 77051
rect 20067 77023 20101 77051
rect 20129 77023 20163 77051
rect 20191 77023 31299 77051
rect 31327 77023 31361 77051
rect 31389 77023 35337 77051
rect 35365 77023 35399 77051
rect 35427 77023 35461 77051
rect 35489 77023 35523 77051
rect 35551 77023 46659 77051
rect 46687 77023 46721 77051
rect 46749 77023 50697 77051
rect 50725 77023 50759 77051
rect 50787 77023 50821 77051
rect 50849 77023 50883 77051
rect 50911 77023 62019 77051
rect 62047 77023 62081 77051
rect 62109 77023 66057 77051
rect 66085 77023 66119 77051
rect 66147 77023 66181 77051
rect 66209 77023 66243 77051
rect 66271 77023 77379 77051
rect 77407 77023 77441 77051
rect 77469 77023 81417 77051
rect 81445 77023 81479 77051
rect 81507 77023 81541 77051
rect 81569 77023 81603 77051
rect 81631 77023 92739 77051
rect 92767 77023 92801 77051
rect 92829 77023 96777 77051
rect 96805 77023 96839 77051
rect 96867 77023 96901 77051
rect 96929 77023 96963 77051
rect 96991 77023 108099 77051
rect 108127 77023 108161 77051
rect 108189 77023 112137 77051
rect 112165 77023 112199 77051
rect 112227 77023 112261 77051
rect 112289 77023 112323 77051
rect 112351 77023 123459 77051
rect 123487 77023 123521 77051
rect 123549 77023 127497 77051
rect 127525 77023 127559 77051
rect 127587 77023 127621 77051
rect 127649 77023 127683 77051
rect 127711 77023 138819 77051
rect 138847 77023 138881 77051
rect 138909 77023 142857 77051
rect 142885 77023 142919 77051
rect 142947 77023 142981 77051
rect 143009 77023 143043 77051
rect 143071 77023 154179 77051
rect 154207 77023 154241 77051
rect 154269 77023 158217 77051
rect 158245 77023 158279 77051
rect 158307 77023 158341 77051
rect 158369 77023 158403 77051
rect 158431 77023 169539 77051
rect 169567 77023 169601 77051
rect 169629 77023 173577 77051
rect 173605 77023 173639 77051
rect 173667 77023 173701 77051
rect 173729 77023 173763 77051
rect 173791 77023 184899 77051
rect 184927 77023 184961 77051
rect 184989 77023 188937 77051
rect 188965 77023 188999 77051
rect 189027 77023 189061 77051
rect 189089 77023 189123 77051
rect 189151 77023 200259 77051
rect 200287 77023 200321 77051
rect 200349 77023 204297 77051
rect 204325 77023 204359 77051
rect 204387 77023 204421 77051
rect 204449 77023 204483 77051
rect 204511 77023 215619 77051
rect 215647 77023 215681 77051
rect 215709 77023 219657 77051
rect 219685 77023 219719 77051
rect 219747 77023 219781 77051
rect 219809 77023 219843 77051
rect 219871 77023 230979 77051
rect 231007 77023 231041 77051
rect 231069 77023 235017 77051
rect 235045 77023 235079 77051
rect 235107 77023 235141 77051
rect 235169 77023 235203 77051
rect 235231 77023 246339 77051
rect 246367 77023 246401 77051
rect 246429 77023 250377 77051
rect 250405 77023 250439 77051
rect 250467 77023 250501 77051
rect 250529 77023 250563 77051
rect 250591 77023 261699 77051
rect 261727 77023 261761 77051
rect 261789 77023 265737 77051
rect 265765 77023 265799 77051
rect 265827 77023 265861 77051
rect 265889 77023 265923 77051
rect 265951 77023 277059 77051
rect 277087 77023 277121 77051
rect 277149 77023 281097 77051
rect 281125 77023 281159 77051
rect 281187 77023 281221 77051
rect 281249 77023 281283 77051
rect 281311 77023 296457 77051
rect 296485 77023 296519 77051
rect 296547 77023 296581 77051
rect 296609 77023 296643 77051
rect 296671 77023 298728 77051
rect 298756 77023 298790 77051
rect 298818 77023 298852 77051
rect 298880 77023 298914 77051
rect 298942 77023 298990 77051
rect -958 76989 298990 77023
rect -958 76961 -910 76989
rect -882 76961 -848 76989
rect -820 76961 -786 76989
rect -758 76961 -724 76989
rect -696 76961 4617 76989
rect 4645 76961 4679 76989
rect 4707 76961 4741 76989
rect 4769 76961 4803 76989
rect 4831 76961 15939 76989
rect 15967 76961 16001 76989
rect 16029 76961 19977 76989
rect 20005 76961 20039 76989
rect 20067 76961 20101 76989
rect 20129 76961 20163 76989
rect 20191 76961 31299 76989
rect 31327 76961 31361 76989
rect 31389 76961 35337 76989
rect 35365 76961 35399 76989
rect 35427 76961 35461 76989
rect 35489 76961 35523 76989
rect 35551 76961 46659 76989
rect 46687 76961 46721 76989
rect 46749 76961 50697 76989
rect 50725 76961 50759 76989
rect 50787 76961 50821 76989
rect 50849 76961 50883 76989
rect 50911 76961 62019 76989
rect 62047 76961 62081 76989
rect 62109 76961 66057 76989
rect 66085 76961 66119 76989
rect 66147 76961 66181 76989
rect 66209 76961 66243 76989
rect 66271 76961 77379 76989
rect 77407 76961 77441 76989
rect 77469 76961 81417 76989
rect 81445 76961 81479 76989
rect 81507 76961 81541 76989
rect 81569 76961 81603 76989
rect 81631 76961 92739 76989
rect 92767 76961 92801 76989
rect 92829 76961 96777 76989
rect 96805 76961 96839 76989
rect 96867 76961 96901 76989
rect 96929 76961 96963 76989
rect 96991 76961 108099 76989
rect 108127 76961 108161 76989
rect 108189 76961 112137 76989
rect 112165 76961 112199 76989
rect 112227 76961 112261 76989
rect 112289 76961 112323 76989
rect 112351 76961 123459 76989
rect 123487 76961 123521 76989
rect 123549 76961 127497 76989
rect 127525 76961 127559 76989
rect 127587 76961 127621 76989
rect 127649 76961 127683 76989
rect 127711 76961 138819 76989
rect 138847 76961 138881 76989
rect 138909 76961 142857 76989
rect 142885 76961 142919 76989
rect 142947 76961 142981 76989
rect 143009 76961 143043 76989
rect 143071 76961 154179 76989
rect 154207 76961 154241 76989
rect 154269 76961 158217 76989
rect 158245 76961 158279 76989
rect 158307 76961 158341 76989
rect 158369 76961 158403 76989
rect 158431 76961 169539 76989
rect 169567 76961 169601 76989
rect 169629 76961 173577 76989
rect 173605 76961 173639 76989
rect 173667 76961 173701 76989
rect 173729 76961 173763 76989
rect 173791 76961 184899 76989
rect 184927 76961 184961 76989
rect 184989 76961 188937 76989
rect 188965 76961 188999 76989
rect 189027 76961 189061 76989
rect 189089 76961 189123 76989
rect 189151 76961 200259 76989
rect 200287 76961 200321 76989
rect 200349 76961 204297 76989
rect 204325 76961 204359 76989
rect 204387 76961 204421 76989
rect 204449 76961 204483 76989
rect 204511 76961 215619 76989
rect 215647 76961 215681 76989
rect 215709 76961 219657 76989
rect 219685 76961 219719 76989
rect 219747 76961 219781 76989
rect 219809 76961 219843 76989
rect 219871 76961 230979 76989
rect 231007 76961 231041 76989
rect 231069 76961 235017 76989
rect 235045 76961 235079 76989
rect 235107 76961 235141 76989
rect 235169 76961 235203 76989
rect 235231 76961 246339 76989
rect 246367 76961 246401 76989
rect 246429 76961 250377 76989
rect 250405 76961 250439 76989
rect 250467 76961 250501 76989
rect 250529 76961 250563 76989
rect 250591 76961 261699 76989
rect 261727 76961 261761 76989
rect 261789 76961 265737 76989
rect 265765 76961 265799 76989
rect 265827 76961 265861 76989
rect 265889 76961 265923 76989
rect 265951 76961 277059 76989
rect 277087 76961 277121 76989
rect 277149 76961 281097 76989
rect 281125 76961 281159 76989
rect 281187 76961 281221 76989
rect 281249 76961 281283 76989
rect 281311 76961 296457 76989
rect 296485 76961 296519 76989
rect 296547 76961 296581 76989
rect 296609 76961 296643 76989
rect 296671 76961 298728 76989
rect 298756 76961 298790 76989
rect 298818 76961 298852 76989
rect 298880 76961 298914 76989
rect 298942 76961 298990 76989
rect -958 76913 298990 76961
rect -958 74175 298990 74223
rect -958 74147 -430 74175
rect -402 74147 -368 74175
rect -340 74147 -306 74175
rect -278 74147 -244 74175
rect -216 74147 2757 74175
rect 2785 74147 2819 74175
rect 2847 74147 2881 74175
rect 2909 74147 2943 74175
rect 2971 74147 8259 74175
rect 8287 74147 8321 74175
rect 8349 74147 18117 74175
rect 18145 74147 18179 74175
rect 18207 74147 18241 74175
rect 18269 74147 18303 74175
rect 18331 74147 23619 74175
rect 23647 74147 23681 74175
rect 23709 74147 33477 74175
rect 33505 74147 33539 74175
rect 33567 74147 33601 74175
rect 33629 74147 33663 74175
rect 33691 74147 38979 74175
rect 39007 74147 39041 74175
rect 39069 74147 48837 74175
rect 48865 74147 48899 74175
rect 48927 74147 48961 74175
rect 48989 74147 49023 74175
rect 49051 74147 54339 74175
rect 54367 74147 54401 74175
rect 54429 74147 64197 74175
rect 64225 74147 64259 74175
rect 64287 74147 64321 74175
rect 64349 74147 64383 74175
rect 64411 74147 69699 74175
rect 69727 74147 69761 74175
rect 69789 74147 79557 74175
rect 79585 74147 79619 74175
rect 79647 74147 79681 74175
rect 79709 74147 79743 74175
rect 79771 74147 85059 74175
rect 85087 74147 85121 74175
rect 85149 74147 94917 74175
rect 94945 74147 94979 74175
rect 95007 74147 95041 74175
rect 95069 74147 95103 74175
rect 95131 74147 100419 74175
rect 100447 74147 100481 74175
rect 100509 74147 110277 74175
rect 110305 74147 110339 74175
rect 110367 74147 110401 74175
rect 110429 74147 110463 74175
rect 110491 74147 115779 74175
rect 115807 74147 115841 74175
rect 115869 74147 125637 74175
rect 125665 74147 125699 74175
rect 125727 74147 125761 74175
rect 125789 74147 125823 74175
rect 125851 74147 131139 74175
rect 131167 74147 131201 74175
rect 131229 74147 140997 74175
rect 141025 74147 141059 74175
rect 141087 74147 141121 74175
rect 141149 74147 141183 74175
rect 141211 74147 146499 74175
rect 146527 74147 146561 74175
rect 146589 74147 156357 74175
rect 156385 74147 156419 74175
rect 156447 74147 156481 74175
rect 156509 74147 156543 74175
rect 156571 74147 161859 74175
rect 161887 74147 161921 74175
rect 161949 74147 171717 74175
rect 171745 74147 171779 74175
rect 171807 74147 171841 74175
rect 171869 74147 171903 74175
rect 171931 74147 177219 74175
rect 177247 74147 177281 74175
rect 177309 74147 187077 74175
rect 187105 74147 187139 74175
rect 187167 74147 187201 74175
rect 187229 74147 187263 74175
rect 187291 74147 192579 74175
rect 192607 74147 192641 74175
rect 192669 74147 202437 74175
rect 202465 74147 202499 74175
rect 202527 74147 202561 74175
rect 202589 74147 202623 74175
rect 202651 74147 207939 74175
rect 207967 74147 208001 74175
rect 208029 74147 217797 74175
rect 217825 74147 217859 74175
rect 217887 74147 217921 74175
rect 217949 74147 217983 74175
rect 218011 74147 223299 74175
rect 223327 74147 223361 74175
rect 223389 74147 233157 74175
rect 233185 74147 233219 74175
rect 233247 74147 233281 74175
rect 233309 74147 233343 74175
rect 233371 74147 238659 74175
rect 238687 74147 238721 74175
rect 238749 74147 248517 74175
rect 248545 74147 248579 74175
rect 248607 74147 248641 74175
rect 248669 74147 248703 74175
rect 248731 74147 254019 74175
rect 254047 74147 254081 74175
rect 254109 74147 263877 74175
rect 263905 74147 263939 74175
rect 263967 74147 264001 74175
rect 264029 74147 264063 74175
rect 264091 74147 269379 74175
rect 269407 74147 269441 74175
rect 269469 74147 279237 74175
rect 279265 74147 279299 74175
rect 279327 74147 279361 74175
rect 279389 74147 279423 74175
rect 279451 74147 284739 74175
rect 284767 74147 284801 74175
rect 284829 74147 294597 74175
rect 294625 74147 294659 74175
rect 294687 74147 294721 74175
rect 294749 74147 294783 74175
rect 294811 74147 298248 74175
rect 298276 74147 298310 74175
rect 298338 74147 298372 74175
rect 298400 74147 298434 74175
rect 298462 74147 298990 74175
rect -958 74113 298990 74147
rect -958 74085 -430 74113
rect -402 74085 -368 74113
rect -340 74085 -306 74113
rect -278 74085 -244 74113
rect -216 74085 2757 74113
rect 2785 74085 2819 74113
rect 2847 74085 2881 74113
rect 2909 74085 2943 74113
rect 2971 74085 8259 74113
rect 8287 74085 8321 74113
rect 8349 74085 18117 74113
rect 18145 74085 18179 74113
rect 18207 74085 18241 74113
rect 18269 74085 18303 74113
rect 18331 74085 23619 74113
rect 23647 74085 23681 74113
rect 23709 74085 33477 74113
rect 33505 74085 33539 74113
rect 33567 74085 33601 74113
rect 33629 74085 33663 74113
rect 33691 74085 38979 74113
rect 39007 74085 39041 74113
rect 39069 74085 48837 74113
rect 48865 74085 48899 74113
rect 48927 74085 48961 74113
rect 48989 74085 49023 74113
rect 49051 74085 54339 74113
rect 54367 74085 54401 74113
rect 54429 74085 64197 74113
rect 64225 74085 64259 74113
rect 64287 74085 64321 74113
rect 64349 74085 64383 74113
rect 64411 74085 69699 74113
rect 69727 74085 69761 74113
rect 69789 74085 79557 74113
rect 79585 74085 79619 74113
rect 79647 74085 79681 74113
rect 79709 74085 79743 74113
rect 79771 74085 85059 74113
rect 85087 74085 85121 74113
rect 85149 74085 94917 74113
rect 94945 74085 94979 74113
rect 95007 74085 95041 74113
rect 95069 74085 95103 74113
rect 95131 74085 100419 74113
rect 100447 74085 100481 74113
rect 100509 74085 110277 74113
rect 110305 74085 110339 74113
rect 110367 74085 110401 74113
rect 110429 74085 110463 74113
rect 110491 74085 115779 74113
rect 115807 74085 115841 74113
rect 115869 74085 125637 74113
rect 125665 74085 125699 74113
rect 125727 74085 125761 74113
rect 125789 74085 125823 74113
rect 125851 74085 131139 74113
rect 131167 74085 131201 74113
rect 131229 74085 140997 74113
rect 141025 74085 141059 74113
rect 141087 74085 141121 74113
rect 141149 74085 141183 74113
rect 141211 74085 146499 74113
rect 146527 74085 146561 74113
rect 146589 74085 156357 74113
rect 156385 74085 156419 74113
rect 156447 74085 156481 74113
rect 156509 74085 156543 74113
rect 156571 74085 161859 74113
rect 161887 74085 161921 74113
rect 161949 74085 171717 74113
rect 171745 74085 171779 74113
rect 171807 74085 171841 74113
rect 171869 74085 171903 74113
rect 171931 74085 177219 74113
rect 177247 74085 177281 74113
rect 177309 74085 187077 74113
rect 187105 74085 187139 74113
rect 187167 74085 187201 74113
rect 187229 74085 187263 74113
rect 187291 74085 192579 74113
rect 192607 74085 192641 74113
rect 192669 74085 202437 74113
rect 202465 74085 202499 74113
rect 202527 74085 202561 74113
rect 202589 74085 202623 74113
rect 202651 74085 207939 74113
rect 207967 74085 208001 74113
rect 208029 74085 217797 74113
rect 217825 74085 217859 74113
rect 217887 74085 217921 74113
rect 217949 74085 217983 74113
rect 218011 74085 223299 74113
rect 223327 74085 223361 74113
rect 223389 74085 233157 74113
rect 233185 74085 233219 74113
rect 233247 74085 233281 74113
rect 233309 74085 233343 74113
rect 233371 74085 238659 74113
rect 238687 74085 238721 74113
rect 238749 74085 248517 74113
rect 248545 74085 248579 74113
rect 248607 74085 248641 74113
rect 248669 74085 248703 74113
rect 248731 74085 254019 74113
rect 254047 74085 254081 74113
rect 254109 74085 263877 74113
rect 263905 74085 263939 74113
rect 263967 74085 264001 74113
rect 264029 74085 264063 74113
rect 264091 74085 269379 74113
rect 269407 74085 269441 74113
rect 269469 74085 279237 74113
rect 279265 74085 279299 74113
rect 279327 74085 279361 74113
rect 279389 74085 279423 74113
rect 279451 74085 284739 74113
rect 284767 74085 284801 74113
rect 284829 74085 294597 74113
rect 294625 74085 294659 74113
rect 294687 74085 294721 74113
rect 294749 74085 294783 74113
rect 294811 74085 298248 74113
rect 298276 74085 298310 74113
rect 298338 74085 298372 74113
rect 298400 74085 298434 74113
rect 298462 74085 298990 74113
rect -958 74051 298990 74085
rect -958 74023 -430 74051
rect -402 74023 -368 74051
rect -340 74023 -306 74051
rect -278 74023 -244 74051
rect -216 74023 2757 74051
rect 2785 74023 2819 74051
rect 2847 74023 2881 74051
rect 2909 74023 2943 74051
rect 2971 74023 8259 74051
rect 8287 74023 8321 74051
rect 8349 74023 18117 74051
rect 18145 74023 18179 74051
rect 18207 74023 18241 74051
rect 18269 74023 18303 74051
rect 18331 74023 23619 74051
rect 23647 74023 23681 74051
rect 23709 74023 33477 74051
rect 33505 74023 33539 74051
rect 33567 74023 33601 74051
rect 33629 74023 33663 74051
rect 33691 74023 38979 74051
rect 39007 74023 39041 74051
rect 39069 74023 48837 74051
rect 48865 74023 48899 74051
rect 48927 74023 48961 74051
rect 48989 74023 49023 74051
rect 49051 74023 54339 74051
rect 54367 74023 54401 74051
rect 54429 74023 64197 74051
rect 64225 74023 64259 74051
rect 64287 74023 64321 74051
rect 64349 74023 64383 74051
rect 64411 74023 69699 74051
rect 69727 74023 69761 74051
rect 69789 74023 79557 74051
rect 79585 74023 79619 74051
rect 79647 74023 79681 74051
rect 79709 74023 79743 74051
rect 79771 74023 85059 74051
rect 85087 74023 85121 74051
rect 85149 74023 94917 74051
rect 94945 74023 94979 74051
rect 95007 74023 95041 74051
rect 95069 74023 95103 74051
rect 95131 74023 100419 74051
rect 100447 74023 100481 74051
rect 100509 74023 110277 74051
rect 110305 74023 110339 74051
rect 110367 74023 110401 74051
rect 110429 74023 110463 74051
rect 110491 74023 115779 74051
rect 115807 74023 115841 74051
rect 115869 74023 125637 74051
rect 125665 74023 125699 74051
rect 125727 74023 125761 74051
rect 125789 74023 125823 74051
rect 125851 74023 131139 74051
rect 131167 74023 131201 74051
rect 131229 74023 140997 74051
rect 141025 74023 141059 74051
rect 141087 74023 141121 74051
rect 141149 74023 141183 74051
rect 141211 74023 146499 74051
rect 146527 74023 146561 74051
rect 146589 74023 156357 74051
rect 156385 74023 156419 74051
rect 156447 74023 156481 74051
rect 156509 74023 156543 74051
rect 156571 74023 161859 74051
rect 161887 74023 161921 74051
rect 161949 74023 171717 74051
rect 171745 74023 171779 74051
rect 171807 74023 171841 74051
rect 171869 74023 171903 74051
rect 171931 74023 177219 74051
rect 177247 74023 177281 74051
rect 177309 74023 187077 74051
rect 187105 74023 187139 74051
rect 187167 74023 187201 74051
rect 187229 74023 187263 74051
rect 187291 74023 192579 74051
rect 192607 74023 192641 74051
rect 192669 74023 202437 74051
rect 202465 74023 202499 74051
rect 202527 74023 202561 74051
rect 202589 74023 202623 74051
rect 202651 74023 207939 74051
rect 207967 74023 208001 74051
rect 208029 74023 217797 74051
rect 217825 74023 217859 74051
rect 217887 74023 217921 74051
rect 217949 74023 217983 74051
rect 218011 74023 223299 74051
rect 223327 74023 223361 74051
rect 223389 74023 233157 74051
rect 233185 74023 233219 74051
rect 233247 74023 233281 74051
rect 233309 74023 233343 74051
rect 233371 74023 238659 74051
rect 238687 74023 238721 74051
rect 238749 74023 248517 74051
rect 248545 74023 248579 74051
rect 248607 74023 248641 74051
rect 248669 74023 248703 74051
rect 248731 74023 254019 74051
rect 254047 74023 254081 74051
rect 254109 74023 263877 74051
rect 263905 74023 263939 74051
rect 263967 74023 264001 74051
rect 264029 74023 264063 74051
rect 264091 74023 269379 74051
rect 269407 74023 269441 74051
rect 269469 74023 279237 74051
rect 279265 74023 279299 74051
rect 279327 74023 279361 74051
rect 279389 74023 279423 74051
rect 279451 74023 284739 74051
rect 284767 74023 284801 74051
rect 284829 74023 294597 74051
rect 294625 74023 294659 74051
rect 294687 74023 294721 74051
rect 294749 74023 294783 74051
rect 294811 74023 298248 74051
rect 298276 74023 298310 74051
rect 298338 74023 298372 74051
rect 298400 74023 298434 74051
rect 298462 74023 298990 74051
rect -958 73989 298990 74023
rect -958 73961 -430 73989
rect -402 73961 -368 73989
rect -340 73961 -306 73989
rect -278 73961 -244 73989
rect -216 73961 2757 73989
rect 2785 73961 2819 73989
rect 2847 73961 2881 73989
rect 2909 73961 2943 73989
rect 2971 73961 8259 73989
rect 8287 73961 8321 73989
rect 8349 73961 18117 73989
rect 18145 73961 18179 73989
rect 18207 73961 18241 73989
rect 18269 73961 18303 73989
rect 18331 73961 23619 73989
rect 23647 73961 23681 73989
rect 23709 73961 33477 73989
rect 33505 73961 33539 73989
rect 33567 73961 33601 73989
rect 33629 73961 33663 73989
rect 33691 73961 38979 73989
rect 39007 73961 39041 73989
rect 39069 73961 48837 73989
rect 48865 73961 48899 73989
rect 48927 73961 48961 73989
rect 48989 73961 49023 73989
rect 49051 73961 54339 73989
rect 54367 73961 54401 73989
rect 54429 73961 64197 73989
rect 64225 73961 64259 73989
rect 64287 73961 64321 73989
rect 64349 73961 64383 73989
rect 64411 73961 69699 73989
rect 69727 73961 69761 73989
rect 69789 73961 79557 73989
rect 79585 73961 79619 73989
rect 79647 73961 79681 73989
rect 79709 73961 79743 73989
rect 79771 73961 85059 73989
rect 85087 73961 85121 73989
rect 85149 73961 94917 73989
rect 94945 73961 94979 73989
rect 95007 73961 95041 73989
rect 95069 73961 95103 73989
rect 95131 73961 100419 73989
rect 100447 73961 100481 73989
rect 100509 73961 110277 73989
rect 110305 73961 110339 73989
rect 110367 73961 110401 73989
rect 110429 73961 110463 73989
rect 110491 73961 115779 73989
rect 115807 73961 115841 73989
rect 115869 73961 125637 73989
rect 125665 73961 125699 73989
rect 125727 73961 125761 73989
rect 125789 73961 125823 73989
rect 125851 73961 131139 73989
rect 131167 73961 131201 73989
rect 131229 73961 140997 73989
rect 141025 73961 141059 73989
rect 141087 73961 141121 73989
rect 141149 73961 141183 73989
rect 141211 73961 146499 73989
rect 146527 73961 146561 73989
rect 146589 73961 156357 73989
rect 156385 73961 156419 73989
rect 156447 73961 156481 73989
rect 156509 73961 156543 73989
rect 156571 73961 161859 73989
rect 161887 73961 161921 73989
rect 161949 73961 171717 73989
rect 171745 73961 171779 73989
rect 171807 73961 171841 73989
rect 171869 73961 171903 73989
rect 171931 73961 177219 73989
rect 177247 73961 177281 73989
rect 177309 73961 187077 73989
rect 187105 73961 187139 73989
rect 187167 73961 187201 73989
rect 187229 73961 187263 73989
rect 187291 73961 192579 73989
rect 192607 73961 192641 73989
rect 192669 73961 202437 73989
rect 202465 73961 202499 73989
rect 202527 73961 202561 73989
rect 202589 73961 202623 73989
rect 202651 73961 207939 73989
rect 207967 73961 208001 73989
rect 208029 73961 217797 73989
rect 217825 73961 217859 73989
rect 217887 73961 217921 73989
rect 217949 73961 217983 73989
rect 218011 73961 223299 73989
rect 223327 73961 223361 73989
rect 223389 73961 233157 73989
rect 233185 73961 233219 73989
rect 233247 73961 233281 73989
rect 233309 73961 233343 73989
rect 233371 73961 238659 73989
rect 238687 73961 238721 73989
rect 238749 73961 248517 73989
rect 248545 73961 248579 73989
rect 248607 73961 248641 73989
rect 248669 73961 248703 73989
rect 248731 73961 254019 73989
rect 254047 73961 254081 73989
rect 254109 73961 263877 73989
rect 263905 73961 263939 73989
rect 263967 73961 264001 73989
rect 264029 73961 264063 73989
rect 264091 73961 269379 73989
rect 269407 73961 269441 73989
rect 269469 73961 279237 73989
rect 279265 73961 279299 73989
rect 279327 73961 279361 73989
rect 279389 73961 279423 73989
rect 279451 73961 284739 73989
rect 284767 73961 284801 73989
rect 284829 73961 294597 73989
rect 294625 73961 294659 73989
rect 294687 73961 294721 73989
rect 294749 73961 294783 73989
rect 294811 73961 298248 73989
rect 298276 73961 298310 73989
rect 298338 73961 298372 73989
rect 298400 73961 298434 73989
rect 298462 73961 298990 73989
rect -958 73913 298990 73961
rect -958 68175 298990 68223
rect -958 68147 -910 68175
rect -882 68147 -848 68175
rect -820 68147 -786 68175
rect -758 68147 -724 68175
rect -696 68147 4617 68175
rect 4645 68147 4679 68175
rect 4707 68147 4741 68175
rect 4769 68147 4803 68175
rect 4831 68147 15939 68175
rect 15967 68147 16001 68175
rect 16029 68147 19977 68175
rect 20005 68147 20039 68175
rect 20067 68147 20101 68175
rect 20129 68147 20163 68175
rect 20191 68147 31299 68175
rect 31327 68147 31361 68175
rect 31389 68147 35337 68175
rect 35365 68147 35399 68175
rect 35427 68147 35461 68175
rect 35489 68147 35523 68175
rect 35551 68147 46659 68175
rect 46687 68147 46721 68175
rect 46749 68147 50697 68175
rect 50725 68147 50759 68175
rect 50787 68147 50821 68175
rect 50849 68147 50883 68175
rect 50911 68147 62019 68175
rect 62047 68147 62081 68175
rect 62109 68147 66057 68175
rect 66085 68147 66119 68175
rect 66147 68147 66181 68175
rect 66209 68147 66243 68175
rect 66271 68147 77379 68175
rect 77407 68147 77441 68175
rect 77469 68147 81417 68175
rect 81445 68147 81479 68175
rect 81507 68147 81541 68175
rect 81569 68147 81603 68175
rect 81631 68147 92739 68175
rect 92767 68147 92801 68175
rect 92829 68147 96777 68175
rect 96805 68147 96839 68175
rect 96867 68147 96901 68175
rect 96929 68147 96963 68175
rect 96991 68147 108099 68175
rect 108127 68147 108161 68175
rect 108189 68147 112137 68175
rect 112165 68147 112199 68175
rect 112227 68147 112261 68175
rect 112289 68147 112323 68175
rect 112351 68147 123459 68175
rect 123487 68147 123521 68175
rect 123549 68147 127497 68175
rect 127525 68147 127559 68175
rect 127587 68147 127621 68175
rect 127649 68147 127683 68175
rect 127711 68147 138819 68175
rect 138847 68147 138881 68175
rect 138909 68147 142857 68175
rect 142885 68147 142919 68175
rect 142947 68147 142981 68175
rect 143009 68147 143043 68175
rect 143071 68147 154179 68175
rect 154207 68147 154241 68175
rect 154269 68147 158217 68175
rect 158245 68147 158279 68175
rect 158307 68147 158341 68175
rect 158369 68147 158403 68175
rect 158431 68147 169539 68175
rect 169567 68147 169601 68175
rect 169629 68147 173577 68175
rect 173605 68147 173639 68175
rect 173667 68147 173701 68175
rect 173729 68147 173763 68175
rect 173791 68147 184899 68175
rect 184927 68147 184961 68175
rect 184989 68147 188937 68175
rect 188965 68147 188999 68175
rect 189027 68147 189061 68175
rect 189089 68147 189123 68175
rect 189151 68147 200259 68175
rect 200287 68147 200321 68175
rect 200349 68147 204297 68175
rect 204325 68147 204359 68175
rect 204387 68147 204421 68175
rect 204449 68147 204483 68175
rect 204511 68147 215619 68175
rect 215647 68147 215681 68175
rect 215709 68147 219657 68175
rect 219685 68147 219719 68175
rect 219747 68147 219781 68175
rect 219809 68147 219843 68175
rect 219871 68147 230979 68175
rect 231007 68147 231041 68175
rect 231069 68147 235017 68175
rect 235045 68147 235079 68175
rect 235107 68147 235141 68175
rect 235169 68147 235203 68175
rect 235231 68147 246339 68175
rect 246367 68147 246401 68175
rect 246429 68147 250377 68175
rect 250405 68147 250439 68175
rect 250467 68147 250501 68175
rect 250529 68147 250563 68175
rect 250591 68147 261699 68175
rect 261727 68147 261761 68175
rect 261789 68147 265737 68175
rect 265765 68147 265799 68175
rect 265827 68147 265861 68175
rect 265889 68147 265923 68175
rect 265951 68147 277059 68175
rect 277087 68147 277121 68175
rect 277149 68147 281097 68175
rect 281125 68147 281159 68175
rect 281187 68147 281221 68175
rect 281249 68147 281283 68175
rect 281311 68147 296457 68175
rect 296485 68147 296519 68175
rect 296547 68147 296581 68175
rect 296609 68147 296643 68175
rect 296671 68147 298728 68175
rect 298756 68147 298790 68175
rect 298818 68147 298852 68175
rect 298880 68147 298914 68175
rect 298942 68147 298990 68175
rect -958 68113 298990 68147
rect -958 68085 -910 68113
rect -882 68085 -848 68113
rect -820 68085 -786 68113
rect -758 68085 -724 68113
rect -696 68085 4617 68113
rect 4645 68085 4679 68113
rect 4707 68085 4741 68113
rect 4769 68085 4803 68113
rect 4831 68085 15939 68113
rect 15967 68085 16001 68113
rect 16029 68085 19977 68113
rect 20005 68085 20039 68113
rect 20067 68085 20101 68113
rect 20129 68085 20163 68113
rect 20191 68085 31299 68113
rect 31327 68085 31361 68113
rect 31389 68085 35337 68113
rect 35365 68085 35399 68113
rect 35427 68085 35461 68113
rect 35489 68085 35523 68113
rect 35551 68085 46659 68113
rect 46687 68085 46721 68113
rect 46749 68085 50697 68113
rect 50725 68085 50759 68113
rect 50787 68085 50821 68113
rect 50849 68085 50883 68113
rect 50911 68085 62019 68113
rect 62047 68085 62081 68113
rect 62109 68085 66057 68113
rect 66085 68085 66119 68113
rect 66147 68085 66181 68113
rect 66209 68085 66243 68113
rect 66271 68085 77379 68113
rect 77407 68085 77441 68113
rect 77469 68085 81417 68113
rect 81445 68085 81479 68113
rect 81507 68085 81541 68113
rect 81569 68085 81603 68113
rect 81631 68085 92739 68113
rect 92767 68085 92801 68113
rect 92829 68085 96777 68113
rect 96805 68085 96839 68113
rect 96867 68085 96901 68113
rect 96929 68085 96963 68113
rect 96991 68085 108099 68113
rect 108127 68085 108161 68113
rect 108189 68085 112137 68113
rect 112165 68085 112199 68113
rect 112227 68085 112261 68113
rect 112289 68085 112323 68113
rect 112351 68085 123459 68113
rect 123487 68085 123521 68113
rect 123549 68085 127497 68113
rect 127525 68085 127559 68113
rect 127587 68085 127621 68113
rect 127649 68085 127683 68113
rect 127711 68085 138819 68113
rect 138847 68085 138881 68113
rect 138909 68085 142857 68113
rect 142885 68085 142919 68113
rect 142947 68085 142981 68113
rect 143009 68085 143043 68113
rect 143071 68085 154179 68113
rect 154207 68085 154241 68113
rect 154269 68085 158217 68113
rect 158245 68085 158279 68113
rect 158307 68085 158341 68113
rect 158369 68085 158403 68113
rect 158431 68085 169539 68113
rect 169567 68085 169601 68113
rect 169629 68085 173577 68113
rect 173605 68085 173639 68113
rect 173667 68085 173701 68113
rect 173729 68085 173763 68113
rect 173791 68085 184899 68113
rect 184927 68085 184961 68113
rect 184989 68085 188937 68113
rect 188965 68085 188999 68113
rect 189027 68085 189061 68113
rect 189089 68085 189123 68113
rect 189151 68085 200259 68113
rect 200287 68085 200321 68113
rect 200349 68085 204297 68113
rect 204325 68085 204359 68113
rect 204387 68085 204421 68113
rect 204449 68085 204483 68113
rect 204511 68085 215619 68113
rect 215647 68085 215681 68113
rect 215709 68085 219657 68113
rect 219685 68085 219719 68113
rect 219747 68085 219781 68113
rect 219809 68085 219843 68113
rect 219871 68085 230979 68113
rect 231007 68085 231041 68113
rect 231069 68085 235017 68113
rect 235045 68085 235079 68113
rect 235107 68085 235141 68113
rect 235169 68085 235203 68113
rect 235231 68085 246339 68113
rect 246367 68085 246401 68113
rect 246429 68085 250377 68113
rect 250405 68085 250439 68113
rect 250467 68085 250501 68113
rect 250529 68085 250563 68113
rect 250591 68085 261699 68113
rect 261727 68085 261761 68113
rect 261789 68085 265737 68113
rect 265765 68085 265799 68113
rect 265827 68085 265861 68113
rect 265889 68085 265923 68113
rect 265951 68085 277059 68113
rect 277087 68085 277121 68113
rect 277149 68085 281097 68113
rect 281125 68085 281159 68113
rect 281187 68085 281221 68113
rect 281249 68085 281283 68113
rect 281311 68085 296457 68113
rect 296485 68085 296519 68113
rect 296547 68085 296581 68113
rect 296609 68085 296643 68113
rect 296671 68085 298728 68113
rect 298756 68085 298790 68113
rect 298818 68085 298852 68113
rect 298880 68085 298914 68113
rect 298942 68085 298990 68113
rect -958 68051 298990 68085
rect -958 68023 -910 68051
rect -882 68023 -848 68051
rect -820 68023 -786 68051
rect -758 68023 -724 68051
rect -696 68023 4617 68051
rect 4645 68023 4679 68051
rect 4707 68023 4741 68051
rect 4769 68023 4803 68051
rect 4831 68023 15939 68051
rect 15967 68023 16001 68051
rect 16029 68023 19977 68051
rect 20005 68023 20039 68051
rect 20067 68023 20101 68051
rect 20129 68023 20163 68051
rect 20191 68023 31299 68051
rect 31327 68023 31361 68051
rect 31389 68023 35337 68051
rect 35365 68023 35399 68051
rect 35427 68023 35461 68051
rect 35489 68023 35523 68051
rect 35551 68023 46659 68051
rect 46687 68023 46721 68051
rect 46749 68023 50697 68051
rect 50725 68023 50759 68051
rect 50787 68023 50821 68051
rect 50849 68023 50883 68051
rect 50911 68023 62019 68051
rect 62047 68023 62081 68051
rect 62109 68023 66057 68051
rect 66085 68023 66119 68051
rect 66147 68023 66181 68051
rect 66209 68023 66243 68051
rect 66271 68023 77379 68051
rect 77407 68023 77441 68051
rect 77469 68023 81417 68051
rect 81445 68023 81479 68051
rect 81507 68023 81541 68051
rect 81569 68023 81603 68051
rect 81631 68023 92739 68051
rect 92767 68023 92801 68051
rect 92829 68023 96777 68051
rect 96805 68023 96839 68051
rect 96867 68023 96901 68051
rect 96929 68023 96963 68051
rect 96991 68023 108099 68051
rect 108127 68023 108161 68051
rect 108189 68023 112137 68051
rect 112165 68023 112199 68051
rect 112227 68023 112261 68051
rect 112289 68023 112323 68051
rect 112351 68023 123459 68051
rect 123487 68023 123521 68051
rect 123549 68023 127497 68051
rect 127525 68023 127559 68051
rect 127587 68023 127621 68051
rect 127649 68023 127683 68051
rect 127711 68023 138819 68051
rect 138847 68023 138881 68051
rect 138909 68023 142857 68051
rect 142885 68023 142919 68051
rect 142947 68023 142981 68051
rect 143009 68023 143043 68051
rect 143071 68023 154179 68051
rect 154207 68023 154241 68051
rect 154269 68023 158217 68051
rect 158245 68023 158279 68051
rect 158307 68023 158341 68051
rect 158369 68023 158403 68051
rect 158431 68023 169539 68051
rect 169567 68023 169601 68051
rect 169629 68023 173577 68051
rect 173605 68023 173639 68051
rect 173667 68023 173701 68051
rect 173729 68023 173763 68051
rect 173791 68023 184899 68051
rect 184927 68023 184961 68051
rect 184989 68023 188937 68051
rect 188965 68023 188999 68051
rect 189027 68023 189061 68051
rect 189089 68023 189123 68051
rect 189151 68023 200259 68051
rect 200287 68023 200321 68051
rect 200349 68023 204297 68051
rect 204325 68023 204359 68051
rect 204387 68023 204421 68051
rect 204449 68023 204483 68051
rect 204511 68023 215619 68051
rect 215647 68023 215681 68051
rect 215709 68023 219657 68051
rect 219685 68023 219719 68051
rect 219747 68023 219781 68051
rect 219809 68023 219843 68051
rect 219871 68023 230979 68051
rect 231007 68023 231041 68051
rect 231069 68023 235017 68051
rect 235045 68023 235079 68051
rect 235107 68023 235141 68051
rect 235169 68023 235203 68051
rect 235231 68023 246339 68051
rect 246367 68023 246401 68051
rect 246429 68023 250377 68051
rect 250405 68023 250439 68051
rect 250467 68023 250501 68051
rect 250529 68023 250563 68051
rect 250591 68023 261699 68051
rect 261727 68023 261761 68051
rect 261789 68023 265737 68051
rect 265765 68023 265799 68051
rect 265827 68023 265861 68051
rect 265889 68023 265923 68051
rect 265951 68023 277059 68051
rect 277087 68023 277121 68051
rect 277149 68023 281097 68051
rect 281125 68023 281159 68051
rect 281187 68023 281221 68051
rect 281249 68023 281283 68051
rect 281311 68023 296457 68051
rect 296485 68023 296519 68051
rect 296547 68023 296581 68051
rect 296609 68023 296643 68051
rect 296671 68023 298728 68051
rect 298756 68023 298790 68051
rect 298818 68023 298852 68051
rect 298880 68023 298914 68051
rect 298942 68023 298990 68051
rect -958 67989 298990 68023
rect -958 67961 -910 67989
rect -882 67961 -848 67989
rect -820 67961 -786 67989
rect -758 67961 -724 67989
rect -696 67961 4617 67989
rect 4645 67961 4679 67989
rect 4707 67961 4741 67989
rect 4769 67961 4803 67989
rect 4831 67961 15939 67989
rect 15967 67961 16001 67989
rect 16029 67961 19977 67989
rect 20005 67961 20039 67989
rect 20067 67961 20101 67989
rect 20129 67961 20163 67989
rect 20191 67961 31299 67989
rect 31327 67961 31361 67989
rect 31389 67961 35337 67989
rect 35365 67961 35399 67989
rect 35427 67961 35461 67989
rect 35489 67961 35523 67989
rect 35551 67961 46659 67989
rect 46687 67961 46721 67989
rect 46749 67961 50697 67989
rect 50725 67961 50759 67989
rect 50787 67961 50821 67989
rect 50849 67961 50883 67989
rect 50911 67961 62019 67989
rect 62047 67961 62081 67989
rect 62109 67961 66057 67989
rect 66085 67961 66119 67989
rect 66147 67961 66181 67989
rect 66209 67961 66243 67989
rect 66271 67961 77379 67989
rect 77407 67961 77441 67989
rect 77469 67961 81417 67989
rect 81445 67961 81479 67989
rect 81507 67961 81541 67989
rect 81569 67961 81603 67989
rect 81631 67961 92739 67989
rect 92767 67961 92801 67989
rect 92829 67961 96777 67989
rect 96805 67961 96839 67989
rect 96867 67961 96901 67989
rect 96929 67961 96963 67989
rect 96991 67961 108099 67989
rect 108127 67961 108161 67989
rect 108189 67961 112137 67989
rect 112165 67961 112199 67989
rect 112227 67961 112261 67989
rect 112289 67961 112323 67989
rect 112351 67961 123459 67989
rect 123487 67961 123521 67989
rect 123549 67961 127497 67989
rect 127525 67961 127559 67989
rect 127587 67961 127621 67989
rect 127649 67961 127683 67989
rect 127711 67961 138819 67989
rect 138847 67961 138881 67989
rect 138909 67961 142857 67989
rect 142885 67961 142919 67989
rect 142947 67961 142981 67989
rect 143009 67961 143043 67989
rect 143071 67961 154179 67989
rect 154207 67961 154241 67989
rect 154269 67961 158217 67989
rect 158245 67961 158279 67989
rect 158307 67961 158341 67989
rect 158369 67961 158403 67989
rect 158431 67961 169539 67989
rect 169567 67961 169601 67989
rect 169629 67961 173577 67989
rect 173605 67961 173639 67989
rect 173667 67961 173701 67989
rect 173729 67961 173763 67989
rect 173791 67961 184899 67989
rect 184927 67961 184961 67989
rect 184989 67961 188937 67989
rect 188965 67961 188999 67989
rect 189027 67961 189061 67989
rect 189089 67961 189123 67989
rect 189151 67961 200259 67989
rect 200287 67961 200321 67989
rect 200349 67961 204297 67989
rect 204325 67961 204359 67989
rect 204387 67961 204421 67989
rect 204449 67961 204483 67989
rect 204511 67961 215619 67989
rect 215647 67961 215681 67989
rect 215709 67961 219657 67989
rect 219685 67961 219719 67989
rect 219747 67961 219781 67989
rect 219809 67961 219843 67989
rect 219871 67961 230979 67989
rect 231007 67961 231041 67989
rect 231069 67961 235017 67989
rect 235045 67961 235079 67989
rect 235107 67961 235141 67989
rect 235169 67961 235203 67989
rect 235231 67961 246339 67989
rect 246367 67961 246401 67989
rect 246429 67961 250377 67989
rect 250405 67961 250439 67989
rect 250467 67961 250501 67989
rect 250529 67961 250563 67989
rect 250591 67961 261699 67989
rect 261727 67961 261761 67989
rect 261789 67961 265737 67989
rect 265765 67961 265799 67989
rect 265827 67961 265861 67989
rect 265889 67961 265923 67989
rect 265951 67961 277059 67989
rect 277087 67961 277121 67989
rect 277149 67961 281097 67989
rect 281125 67961 281159 67989
rect 281187 67961 281221 67989
rect 281249 67961 281283 67989
rect 281311 67961 296457 67989
rect 296485 67961 296519 67989
rect 296547 67961 296581 67989
rect 296609 67961 296643 67989
rect 296671 67961 298728 67989
rect 298756 67961 298790 67989
rect 298818 67961 298852 67989
rect 298880 67961 298914 67989
rect 298942 67961 298990 67989
rect -958 67913 298990 67961
rect -958 65175 298990 65223
rect -958 65147 -430 65175
rect -402 65147 -368 65175
rect -340 65147 -306 65175
rect -278 65147 -244 65175
rect -216 65147 2757 65175
rect 2785 65147 2819 65175
rect 2847 65147 2881 65175
rect 2909 65147 2943 65175
rect 2971 65147 8259 65175
rect 8287 65147 8321 65175
rect 8349 65147 18117 65175
rect 18145 65147 18179 65175
rect 18207 65147 18241 65175
rect 18269 65147 18303 65175
rect 18331 65147 23619 65175
rect 23647 65147 23681 65175
rect 23709 65147 33477 65175
rect 33505 65147 33539 65175
rect 33567 65147 33601 65175
rect 33629 65147 33663 65175
rect 33691 65147 38979 65175
rect 39007 65147 39041 65175
rect 39069 65147 48837 65175
rect 48865 65147 48899 65175
rect 48927 65147 48961 65175
rect 48989 65147 49023 65175
rect 49051 65147 54339 65175
rect 54367 65147 54401 65175
rect 54429 65147 64197 65175
rect 64225 65147 64259 65175
rect 64287 65147 64321 65175
rect 64349 65147 64383 65175
rect 64411 65147 69699 65175
rect 69727 65147 69761 65175
rect 69789 65147 79557 65175
rect 79585 65147 79619 65175
rect 79647 65147 79681 65175
rect 79709 65147 79743 65175
rect 79771 65147 85059 65175
rect 85087 65147 85121 65175
rect 85149 65147 94917 65175
rect 94945 65147 94979 65175
rect 95007 65147 95041 65175
rect 95069 65147 95103 65175
rect 95131 65147 100419 65175
rect 100447 65147 100481 65175
rect 100509 65147 110277 65175
rect 110305 65147 110339 65175
rect 110367 65147 110401 65175
rect 110429 65147 110463 65175
rect 110491 65147 115779 65175
rect 115807 65147 115841 65175
rect 115869 65147 125637 65175
rect 125665 65147 125699 65175
rect 125727 65147 125761 65175
rect 125789 65147 125823 65175
rect 125851 65147 131139 65175
rect 131167 65147 131201 65175
rect 131229 65147 140997 65175
rect 141025 65147 141059 65175
rect 141087 65147 141121 65175
rect 141149 65147 141183 65175
rect 141211 65147 146499 65175
rect 146527 65147 146561 65175
rect 146589 65147 156357 65175
rect 156385 65147 156419 65175
rect 156447 65147 156481 65175
rect 156509 65147 156543 65175
rect 156571 65147 161859 65175
rect 161887 65147 161921 65175
rect 161949 65147 171717 65175
rect 171745 65147 171779 65175
rect 171807 65147 171841 65175
rect 171869 65147 171903 65175
rect 171931 65147 177219 65175
rect 177247 65147 177281 65175
rect 177309 65147 187077 65175
rect 187105 65147 187139 65175
rect 187167 65147 187201 65175
rect 187229 65147 187263 65175
rect 187291 65147 192579 65175
rect 192607 65147 192641 65175
rect 192669 65147 202437 65175
rect 202465 65147 202499 65175
rect 202527 65147 202561 65175
rect 202589 65147 202623 65175
rect 202651 65147 207939 65175
rect 207967 65147 208001 65175
rect 208029 65147 217797 65175
rect 217825 65147 217859 65175
rect 217887 65147 217921 65175
rect 217949 65147 217983 65175
rect 218011 65147 223299 65175
rect 223327 65147 223361 65175
rect 223389 65147 233157 65175
rect 233185 65147 233219 65175
rect 233247 65147 233281 65175
rect 233309 65147 233343 65175
rect 233371 65147 238659 65175
rect 238687 65147 238721 65175
rect 238749 65147 248517 65175
rect 248545 65147 248579 65175
rect 248607 65147 248641 65175
rect 248669 65147 248703 65175
rect 248731 65147 254019 65175
rect 254047 65147 254081 65175
rect 254109 65147 263877 65175
rect 263905 65147 263939 65175
rect 263967 65147 264001 65175
rect 264029 65147 264063 65175
rect 264091 65147 269379 65175
rect 269407 65147 269441 65175
rect 269469 65147 279237 65175
rect 279265 65147 279299 65175
rect 279327 65147 279361 65175
rect 279389 65147 279423 65175
rect 279451 65147 284739 65175
rect 284767 65147 284801 65175
rect 284829 65147 294597 65175
rect 294625 65147 294659 65175
rect 294687 65147 294721 65175
rect 294749 65147 294783 65175
rect 294811 65147 298248 65175
rect 298276 65147 298310 65175
rect 298338 65147 298372 65175
rect 298400 65147 298434 65175
rect 298462 65147 298990 65175
rect -958 65113 298990 65147
rect -958 65085 -430 65113
rect -402 65085 -368 65113
rect -340 65085 -306 65113
rect -278 65085 -244 65113
rect -216 65085 2757 65113
rect 2785 65085 2819 65113
rect 2847 65085 2881 65113
rect 2909 65085 2943 65113
rect 2971 65085 8259 65113
rect 8287 65085 8321 65113
rect 8349 65085 18117 65113
rect 18145 65085 18179 65113
rect 18207 65085 18241 65113
rect 18269 65085 18303 65113
rect 18331 65085 23619 65113
rect 23647 65085 23681 65113
rect 23709 65085 33477 65113
rect 33505 65085 33539 65113
rect 33567 65085 33601 65113
rect 33629 65085 33663 65113
rect 33691 65085 38979 65113
rect 39007 65085 39041 65113
rect 39069 65085 48837 65113
rect 48865 65085 48899 65113
rect 48927 65085 48961 65113
rect 48989 65085 49023 65113
rect 49051 65085 54339 65113
rect 54367 65085 54401 65113
rect 54429 65085 64197 65113
rect 64225 65085 64259 65113
rect 64287 65085 64321 65113
rect 64349 65085 64383 65113
rect 64411 65085 69699 65113
rect 69727 65085 69761 65113
rect 69789 65085 79557 65113
rect 79585 65085 79619 65113
rect 79647 65085 79681 65113
rect 79709 65085 79743 65113
rect 79771 65085 85059 65113
rect 85087 65085 85121 65113
rect 85149 65085 94917 65113
rect 94945 65085 94979 65113
rect 95007 65085 95041 65113
rect 95069 65085 95103 65113
rect 95131 65085 100419 65113
rect 100447 65085 100481 65113
rect 100509 65085 110277 65113
rect 110305 65085 110339 65113
rect 110367 65085 110401 65113
rect 110429 65085 110463 65113
rect 110491 65085 115779 65113
rect 115807 65085 115841 65113
rect 115869 65085 125637 65113
rect 125665 65085 125699 65113
rect 125727 65085 125761 65113
rect 125789 65085 125823 65113
rect 125851 65085 131139 65113
rect 131167 65085 131201 65113
rect 131229 65085 140997 65113
rect 141025 65085 141059 65113
rect 141087 65085 141121 65113
rect 141149 65085 141183 65113
rect 141211 65085 146499 65113
rect 146527 65085 146561 65113
rect 146589 65085 156357 65113
rect 156385 65085 156419 65113
rect 156447 65085 156481 65113
rect 156509 65085 156543 65113
rect 156571 65085 161859 65113
rect 161887 65085 161921 65113
rect 161949 65085 171717 65113
rect 171745 65085 171779 65113
rect 171807 65085 171841 65113
rect 171869 65085 171903 65113
rect 171931 65085 177219 65113
rect 177247 65085 177281 65113
rect 177309 65085 187077 65113
rect 187105 65085 187139 65113
rect 187167 65085 187201 65113
rect 187229 65085 187263 65113
rect 187291 65085 192579 65113
rect 192607 65085 192641 65113
rect 192669 65085 202437 65113
rect 202465 65085 202499 65113
rect 202527 65085 202561 65113
rect 202589 65085 202623 65113
rect 202651 65085 207939 65113
rect 207967 65085 208001 65113
rect 208029 65085 217797 65113
rect 217825 65085 217859 65113
rect 217887 65085 217921 65113
rect 217949 65085 217983 65113
rect 218011 65085 223299 65113
rect 223327 65085 223361 65113
rect 223389 65085 233157 65113
rect 233185 65085 233219 65113
rect 233247 65085 233281 65113
rect 233309 65085 233343 65113
rect 233371 65085 238659 65113
rect 238687 65085 238721 65113
rect 238749 65085 248517 65113
rect 248545 65085 248579 65113
rect 248607 65085 248641 65113
rect 248669 65085 248703 65113
rect 248731 65085 254019 65113
rect 254047 65085 254081 65113
rect 254109 65085 263877 65113
rect 263905 65085 263939 65113
rect 263967 65085 264001 65113
rect 264029 65085 264063 65113
rect 264091 65085 269379 65113
rect 269407 65085 269441 65113
rect 269469 65085 279237 65113
rect 279265 65085 279299 65113
rect 279327 65085 279361 65113
rect 279389 65085 279423 65113
rect 279451 65085 284739 65113
rect 284767 65085 284801 65113
rect 284829 65085 294597 65113
rect 294625 65085 294659 65113
rect 294687 65085 294721 65113
rect 294749 65085 294783 65113
rect 294811 65085 298248 65113
rect 298276 65085 298310 65113
rect 298338 65085 298372 65113
rect 298400 65085 298434 65113
rect 298462 65085 298990 65113
rect -958 65051 298990 65085
rect -958 65023 -430 65051
rect -402 65023 -368 65051
rect -340 65023 -306 65051
rect -278 65023 -244 65051
rect -216 65023 2757 65051
rect 2785 65023 2819 65051
rect 2847 65023 2881 65051
rect 2909 65023 2943 65051
rect 2971 65023 8259 65051
rect 8287 65023 8321 65051
rect 8349 65023 18117 65051
rect 18145 65023 18179 65051
rect 18207 65023 18241 65051
rect 18269 65023 18303 65051
rect 18331 65023 23619 65051
rect 23647 65023 23681 65051
rect 23709 65023 33477 65051
rect 33505 65023 33539 65051
rect 33567 65023 33601 65051
rect 33629 65023 33663 65051
rect 33691 65023 38979 65051
rect 39007 65023 39041 65051
rect 39069 65023 48837 65051
rect 48865 65023 48899 65051
rect 48927 65023 48961 65051
rect 48989 65023 49023 65051
rect 49051 65023 54339 65051
rect 54367 65023 54401 65051
rect 54429 65023 64197 65051
rect 64225 65023 64259 65051
rect 64287 65023 64321 65051
rect 64349 65023 64383 65051
rect 64411 65023 69699 65051
rect 69727 65023 69761 65051
rect 69789 65023 79557 65051
rect 79585 65023 79619 65051
rect 79647 65023 79681 65051
rect 79709 65023 79743 65051
rect 79771 65023 85059 65051
rect 85087 65023 85121 65051
rect 85149 65023 94917 65051
rect 94945 65023 94979 65051
rect 95007 65023 95041 65051
rect 95069 65023 95103 65051
rect 95131 65023 100419 65051
rect 100447 65023 100481 65051
rect 100509 65023 110277 65051
rect 110305 65023 110339 65051
rect 110367 65023 110401 65051
rect 110429 65023 110463 65051
rect 110491 65023 115779 65051
rect 115807 65023 115841 65051
rect 115869 65023 125637 65051
rect 125665 65023 125699 65051
rect 125727 65023 125761 65051
rect 125789 65023 125823 65051
rect 125851 65023 131139 65051
rect 131167 65023 131201 65051
rect 131229 65023 140997 65051
rect 141025 65023 141059 65051
rect 141087 65023 141121 65051
rect 141149 65023 141183 65051
rect 141211 65023 146499 65051
rect 146527 65023 146561 65051
rect 146589 65023 156357 65051
rect 156385 65023 156419 65051
rect 156447 65023 156481 65051
rect 156509 65023 156543 65051
rect 156571 65023 161859 65051
rect 161887 65023 161921 65051
rect 161949 65023 171717 65051
rect 171745 65023 171779 65051
rect 171807 65023 171841 65051
rect 171869 65023 171903 65051
rect 171931 65023 177219 65051
rect 177247 65023 177281 65051
rect 177309 65023 187077 65051
rect 187105 65023 187139 65051
rect 187167 65023 187201 65051
rect 187229 65023 187263 65051
rect 187291 65023 192579 65051
rect 192607 65023 192641 65051
rect 192669 65023 202437 65051
rect 202465 65023 202499 65051
rect 202527 65023 202561 65051
rect 202589 65023 202623 65051
rect 202651 65023 207939 65051
rect 207967 65023 208001 65051
rect 208029 65023 217797 65051
rect 217825 65023 217859 65051
rect 217887 65023 217921 65051
rect 217949 65023 217983 65051
rect 218011 65023 223299 65051
rect 223327 65023 223361 65051
rect 223389 65023 233157 65051
rect 233185 65023 233219 65051
rect 233247 65023 233281 65051
rect 233309 65023 233343 65051
rect 233371 65023 238659 65051
rect 238687 65023 238721 65051
rect 238749 65023 248517 65051
rect 248545 65023 248579 65051
rect 248607 65023 248641 65051
rect 248669 65023 248703 65051
rect 248731 65023 254019 65051
rect 254047 65023 254081 65051
rect 254109 65023 263877 65051
rect 263905 65023 263939 65051
rect 263967 65023 264001 65051
rect 264029 65023 264063 65051
rect 264091 65023 269379 65051
rect 269407 65023 269441 65051
rect 269469 65023 279237 65051
rect 279265 65023 279299 65051
rect 279327 65023 279361 65051
rect 279389 65023 279423 65051
rect 279451 65023 284739 65051
rect 284767 65023 284801 65051
rect 284829 65023 294597 65051
rect 294625 65023 294659 65051
rect 294687 65023 294721 65051
rect 294749 65023 294783 65051
rect 294811 65023 298248 65051
rect 298276 65023 298310 65051
rect 298338 65023 298372 65051
rect 298400 65023 298434 65051
rect 298462 65023 298990 65051
rect -958 64989 298990 65023
rect -958 64961 -430 64989
rect -402 64961 -368 64989
rect -340 64961 -306 64989
rect -278 64961 -244 64989
rect -216 64961 2757 64989
rect 2785 64961 2819 64989
rect 2847 64961 2881 64989
rect 2909 64961 2943 64989
rect 2971 64961 8259 64989
rect 8287 64961 8321 64989
rect 8349 64961 18117 64989
rect 18145 64961 18179 64989
rect 18207 64961 18241 64989
rect 18269 64961 18303 64989
rect 18331 64961 23619 64989
rect 23647 64961 23681 64989
rect 23709 64961 33477 64989
rect 33505 64961 33539 64989
rect 33567 64961 33601 64989
rect 33629 64961 33663 64989
rect 33691 64961 38979 64989
rect 39007 64961 39041 64989
rect 39069 64961 48837 64989
rect 48865 64961 48899 64989
rect 48927 64961 48961 64989
rect 48989 64961 49023 64989
rect 49051 64961 54339 64989
rect 54367 64961 54401 64989
rect 54429 64961 64197 64989
rect 64225 64961 64259 64989
rect 64287 64961 64321 64989
rect 64349 64961 64383 64989
rect 64411 64961 69699 64989
rect 69727 64961 69761 64989
rect 69789 64961 79557 64989
rect 79585 64961 79619 64989
rect 79647 64961 79681 64989
rect 79709 64961 79743 64989
rect 79771 64961 85059 64989
rect 85087 64961 85121 64989
rect 85149 64961 94917 64989
rect 94945 64961 94979 64989
rect 95007 64961 95041 64989
rect 95069 64961 95103 64989
rect 95131 64961 100419 64989
rect 100447 64961 100481 64989
rect 100509 64961 110277 64989
rect 110305 64961 110339 64989
rect 110367 64961 110401 64989
rect 110429 64961 110463 64989
rect 110491 64961 115779 64989
rect 115807 64961 115841 64989
rect 115869 64961 125637 64989
rect 125665 64961 125699 64989
rect 125727 64961 125761 64989
rect 125789 64961 125823 64989
rect 125851 64961 131139 64989
rect 131167 64961 131201 64989
rect 131229 64961 140997 64989
rect 141025 64961 141059 64989
rect 141087 64961 141121 64989
rect 141149 64961 141183 64989
rect 141211 64961 146499 64989
rect 146527 64961 146561 64989
rect 146589 64961 156357 64989
rect 156385 64961 156419 64989
rect 156447 64961 156481 64989
rect 156509 64961 156543 64989
rect 156571 64961 161859 64989
rect 161887 64961 161921 64989
rect 161949 64961 171717 64989
rect 171745 64961 171779 64989
rect 171807 64961 171841 64989
rect 171869 64961 171903 64989
rect 171931 64961 177219 64989
rect 177247 64961 177281 64989
rect 177309 64961 187077 64989
rect 187105 64961 187139 64989
rect 187167 64961 187201 64989
rect 187229 64961 187263 64989
rect 187291 64961 192579 64989
rect 192607 64961 192641 64989
rect 192669 64961 202437 64989
rect 202465 64961 202499 64989
rect 202527 64961 202561 64989
rect 202589 64961 202623 64989
rect 202651 64961 207939 64989
rect 207967 64961 208001 64989
rect 208029 64961 217797 64989
rect 217825 64961 217859 64989
rect 217887 64961 217921 64989
rect 217949 64961 217983 64989
rect 218011 64961 223299 64989
rect 223327 64961 223361 64989
rect 223389 64961 233157 64989
rect 233185 64961 233219 64989
rect 233247 64961 233281 64989
rect 233309 64961 233343 64989
rect 233371 64961 238659 64989
rect 238687 64961 238721 64989
rect 238749 64961 248517 64989
rect 248545 64961 248579 64989
rect 248607 64961 248641 64989
rect 248669 64961 248703 64989
rect 248731 64961 254019 64989
rect 254047 64961 254081 64989
rect 254109 64961 263877 64989
rect 263905 64961 263939 64989
rect 263967 64961 264001 64989
rect 264029 64961 264063 64989
rect 264091 64961 269379 64989
rect 269407 64961 269441 64989
rect 269469 64961 279237 64989
rect 279265 64961 279299 64989
rect 279327 64961 279361 64989
rect 279389 64961 279423 64989
rect 279451 64961 284739 64989
rect 284767 64961 284801 64989
rect 284829 64961 294597 64989
rect 294625 64961 294659 64989
rect 294687 64961 294721 64989
rect 294749 64961 294783 64989
rect 294811 64961 298248 64989
rect 298276 64961 298310 64989
rect 298338 64961 298372 64989
rect 298400 64961 298434 64989
rect 298462 64961 298990 64989
rect -958 64913 298990 64961
rect -958 59175 298990 59223
rect -958 59147 -910 59175
rect -882 59147 -848 59175
rect -820 59147 -786 59175
rect -758 59147 -724 59175
rect -696 59147 4617 59175
rect 4645 59147 4679 59175
rect 4707 59147 4741 59175
rect 4769 59147 4803 59175
rect 4831 59147 15939 59175
rect 15967 59147 16001 59175
rect 16029 59147 19977 59175
rect 20005 59147 20039 59175
rect 20067 59147 20101 59175
rect 20129 59147 20163 59175
rect 20191 59147 31299 59175
rect 31327 59147 31361 59175
rect 31389 59147 35337 59175
rect 35365 59147 35399 59175
rect 35427 59147 35461 59175
rect 35489 59147 35523 59175
rect 35551 59147 46659 59175
rect 46687 59147 46721 59175
rect 46749 59147 50697 59175
rect 50725 59147 50759 59175
rect 50787 59147 50821 59175
rect 50849 59147 50883 59175
rect 50911 59147 62019 59175
rect 62047 59147 62081 59175
rect 62109 59147 66057 59175
rect 66085 59147 66119 59175
rect 66147 59147 66181 59175
rect 66209 59147 66243 59175
rect 66271 59147 77379 59175
rect 77407 59147 77441 59175
rect 77469 59147 81417 59175
rect 81445 59147 81479 59175
rect 81507 59147 81541 59175
rect 81569 59147 81603 59175
rect 81631 59147 92739 59175
rect 92767 59147 92801 59175
rect 92829 59147 96777 59175
rect 96805 59147 96839 59175
rect 96867 59147 96901 59175
rect 96929 59147 96963 59175
rect 96991 59147 108099 59175
rect 108127 59147 108161 59175
rect 108189 59147 112137 59175
rect 112165 59147 112199 59175
rect 112227 59147 112261 59175
rect 112289 59147 112323 59175
rect 112351 59147 123459 59175
rect 123487 59147 123521 59175
rect 123549 59147 127497 59175
rect 127525 59147 127559 59175
rect 127587 59147 127621 59175
rect 127649 59147 127683 59175
rect 127711 59147 138819 59175
rect 138847 59147 138881 59175
rect 138909 59147 142857 59175
rect 142885 59147 142919 59175
rect 142947 59147 142981 59175
rect 143009 59147 143043 59175
rect 143071 59147 154179 59175
rect 154207 59147 154241 59175
rect 154269 59147 158217 59175
rect 158245 59147 158279 59175
rect 158307 59147 158341 59175
rect 158369 59147 158403 59175
rect 158431 59147 169539 59175
rect 169567 59147 169601 59175
rect 169629 59147 173577 59175
rect 173605 59147 173639 59175
rect 173667 59147 173701 59175
rect 173729 59147 173763 59175
rect 173791 59147 184899 59175
rect 184927 59147 184961 59175
rect 184989 59147 188937 59175
rect 188965 59147 188999 59175
rect 189027 59147 189061 59175
rect 189089 59147 189123 59175
rect 189151 59147 200259 59175
rect 200287 59147 200321 59175
rect 200349 59147 204297 59175
rect 204325 59147 204359 59175
rect 204387 59147 204421 59175
rect 204449 59147 204483 59175
rect 204511 59147 215619 59175
rect 215647 59147 215681 59175
rect 215709 59147 219657 59175
rect 219685 59147 219719 59175
rect 219747 59147 219781 59175
rect 219809 59147 219843 59175
rect 219871 59147 230979 59175
rect 231007 59147 231041 59175
rect 231069 59147 235017 59175
rect 235045 59147 235079 59175
rect 235107 59147 235141 59175
rect 235169 59147 235203 59175
rect 235231 59147 246339 59175
rect 246367 59147 246401 59175
rect 246429 59147 250377 59175
rect 250405 59147 250439 59175
rect 250467 59147 250501 59175
rect 250529 59147 250563 59175
rect 250591 59147 261699 59175
rect 261727 59147 261761 59175
rect 261789 59147 265737 59175
rect 265765 59147 265799 59175
rect 265827 59147 265861 59175
rect 265889 59147 265923 59175
rect 265951 59147 277059 59175
rect 277087 59147 277121 59175
rect 277149 59147 281097 59175
rect 281125 59147 281159 59175
rect 281187 59147 281221 59175
rect 281249 59147 281283 59175
rect 281311 59147 296457 59175
rect 296485 59147 296519 59175
rect 296547 59147 296581 59175
rect 296609 59147 296643 59175
rect 296671 59147 298728 59175
rect 298756 59147 298790 59175
rect 298818 59147 298852 59175
rect 298880 59147 298914 59175
rect 298942 59147 298990 59175
rect -958 59113 298990 59147
rect -958 59085 -910 59113
rect -882 59085 -848 59113
rect -820 59085 -786 59113
rect -758 59085 -724 59113
rect -696 59085 4617 59113
rect 4645 59085 4679 59113
rect 4707 59085 4741 59113
rect 4769 59085 4803 59113
rect 4831 59085 15939 59113
rect 15967 59085 16001 59113
rect 16029 59085 19977 59113
rect 20005 59085 20039 59113
rect 20067 59085 20101 59113
rect 20129 59085 20163 59113
rect 20191 59085 31299 59113
rect 31327 59085 31361 59113
rect 31389 59085 35337 59113
rect 35365 59085 35399 59113
rect 35427 59085 35461 59113
rect 35489 59085 35523 59113
rect 35551 59085 46659 59113
rect 46687 59085 46721 59113
rect 46749 59085 50697 59113
rect 50725 59085 50759 59113
rect 50787 59085 50821 59113
rect 50849 59085 50883 59113
rect 50911 59085 62019 59113
rect 62047 59085 62081 59113
rect 62109 59085 66057 59113
rect 66085 59085 66119 59113
rect 66147 59085 66181 59113
rect 66209 59085 66243 59113
rect 66271 59085 77379 59113
rect 77407 59085 77441 59113
rect 77469 59085 81417 59113
rect 81445 59085 81479 59113
rect 81507 59085 81541 59113
rect 81569 59085 81603 59113
rect 81631 59085 92739 59113
rect 92767 59085 92801 59113
rect 92829 59085 96777 59113
rect 96805 59085 96839 59113
rect 96867 59085 96901 59113
rect 96929 59085 96963 59113
rect 96991 59085 108099 59113
rect 108127 59085 108161 59113
rect 108189 59085 112137 59113
rect 112165 59085 112199 59113
rect 112227 59085 112261 59113
rect 112289 59085 112323 59113
rect 112351 59085 123459 59113
rect 123487 59085 123521 59113
rect 123549 59085 127497 59113
rect 127525 59085 127559 59113
rect 127587 59085 127621 59113
rect 127649 59085 127683 59113
rect 127711 59085 138819 59113
rect 138847 59085 138881 59113
rect 138909 59085 142857 59113
rect 142885 59085 142919 59113
rect 142947 59085 142981 59113
rect 143009 59085 143043 59113
rect 143071 59085 154179 59113
rect 154207 59085 154241 59113
rect 154269 59085 158217 59113
rect 158245 59085 158279 59113
rect 158307 59085 158341 59113
rect 158369 59085 158403 59113
rect 158431 59085 169539 59113
rect 169567 59085 169601 59113
rect 169629 59085 173577 59113
rect 173605 59085 173639 59113
rect 173667 59085 173701 59113
rect 173729 59085 173763 59113
rect 173791 59085 184899 59113
rect 184927 59085 184961 59113
rect 184989 59085 188937 59113
rect 188965 59085 188999 59113
rect 189027 59085 189061 59113
rect 189089 59085 189123 59113
rect 189151 59085 200259 59113
rect 200287 59085 200321 59113
rect 200349 59085 204297 59113
rect 204325 59085 204359 59113
rect 204387 59085 204421 59113
rect 204449 59085 204483 59113
rect 204511 59085 215619 59113
rect 215647 59085 215681 59113
rect 215709 59085 219657 59113
rect 219685 59085 219719 59113
rect 219747 59085 219781 59113
rect 219809 59085 219843 59113
rect 219871 59085 230979 59113
rect 231007 59085 231041 59113
rect 231069 59085 235017 59113
rect 235045 59085 235079 59113
rect 235107 59085 235141 59113
rect 235169 59085 235203 59113
rect 235231 59085 246339 59113
rect 246367 59085 246401 59113
rect 246429 59085 250377 59113
rect 250405 59085 250439 59113
rect 250467 59085 250501 59113
rect 250529 59085 250563 59113
rect 250591 59085 261699 59113
rect 261727 59085 261761 59113
rect 261789 59085 265737 59113
rect 265765 59085 265799 59113
rect 265827 59085 265861 59113
rect 265889 59085 265923 59113
rect 265951 59085 277059 59113
rect 277087 59085 277121 59113
rect 277149 59085 281097 59113
rect 281125 59085 281159 59113
rect 281187 59085 281221 59113
rect 281249 59085 281283 59113
rect 281311 59085 296457 59113
rect 296485 59085 296519 59113
rect 296547 59085 296581 59113
rect 296609 59085 296643 59113
rect 296671 59085 298728 59113
rect 298756 59085 298790 59113
rect 298818 59085 298852 59113
rect 298880 59085 298914 59113
rect 298942 59085 298990 59113
rect -958 59051 298990 59085
rect -958 59023 -910 59051
rect -882 59023 -848 59051
rect -820 59023 -786 59051
rect -758 59023 -724 59051
rect -696 59023 4617 59051
rect 4645 59023 4679 59051
rect 4707 59023 4741 59051
rect 4769 59023 4803 59051
rect 4831 59023 15939 59051
rect 15967 59023 16001 59051
rect 16029 59023 19977 59051
rect 20005 59023 20039 59051
rect 20067 59023 20101 59051
rect 20129 59023 20163 59051
rect 20191 59023 31299 59051
rect 31327 59023 31361 59051
rect 31389 59023 35337 59051
rect 35365 59023 35399 59051
rect 35427 59023 35461 59051
rect 35489 59023 35523 59051
rect 35551 59023 46659 59051
rect 46687 59023 46721 59051
rect 46749 59023 50697 59051
rect 50725 59023 50759 59051
rect 50787 59023 50821 59051
rect 50849 59023 50883 59051
rect 50911 59023 62019 59051
rect 62047 59023 62081 59051
rect 62109 59023 66057 59051
rect 66085 59023 66119 59051
rect 66147 59023 66181 59051
rect 66209 59023 66243 59051
rect 66271 59023 77379 59051
rect 77407 59023 77441 59051
rect 77469 59023 81417 59051
rect 81445 59023 81479 59051
rect 81507 59023 81541 59051
rect 81569 59023 81603 59051
rect 81631 59023 92739 59051
rect 92767 59023 92801 59051
rect 92829 59023 96777 59051
rect 96805 59023 96839 59051
rect 96867 59023 96901 59051
rect 96929 59023 96963 59051
rect 96991 59023 108099 59051
rect 108127 59023 108161 59051
rect 108189 59023 112137 59051
rect 112165 59023 112199 59051
rect 112227 59023 112261 59051
rect 112289 59023 112323 59051
rect 112351 59023 123459 59051
rect 123487 59023 123521 59051
rect 123549 59023 127497 59051
rect 127525 59023 127559 59051
rect 127587 59023 127621 59051
rect 127649 59023 127683 59051
rect 127711 59023 138819 59051
rect 138847 59023 138881 59051
rect 138909 59023 142857 59051
rect 142885 59023 142919 59051
rect 142947 59023 142981 59051
rect 143009 59023 143043 59051
rect 143071 59023 154179 59051
rect 154207 59023 154241 59051
rect 154269 59023 158217 59051
rect 158245 59023 158279 59051
rect 158307 59023 158341 59051
rect 158369 59023 158403 59051
rect 158431 59023 169539 59051
rect 169567 59023 169601 59051
rect 169629 59023 173577 59051
rect 173605 59023 173639 59051
rect 173667 59023 173701 59051
rect 173729 59023 173763 59051
rect 173791 59023 184899 59051
rect 184927 59023 184961 59051
rect 184989 59023 188937 59051
rect 188965 59023 188999 59051
rect 189027 59023 189061 59051
rect 189089 59023 189123 59051
rect 189151 59023 200259 59051
rect 200287 59023 200321 59051
rect 200349 59023 204297 59051
rect 204325 59023 204359 59051
rect 204387 59023 204421 59051
rect 204449 59023 204483 59051
rect 204511 59023 215619 59051
rect 215647 59023 215681 59051
rect 215709 59023 219657 59051
rect 219685 59023 219719 59051
rect 219747 59023 219781 59051
rect 219809 59023 219843 59051
rect 219871 59023 230979 59051
rect 231007 59023 231041 59051
rect 231069 59023 235017 59051
rect 235045 59023 235079 59051
rect 235107 59023 235141 59051
rect 235169 59023 235203 59051
rect 235231 59023 246339 59051
rect 246367 59023 246401 59051
rect 246429 59023 250377 59051
rect 250405 59023 250439 59051
rect 250467 59023 250501 59051
rect 250529 59023 250563 59051
rect 250591 59023 261699 59051
rect 261727 59023 261761 59051
rect 261789 59023 265737 59051
rect 265765 59023 265799 59051
rect 265827 59023 265861 59051
rect 265889 59023 265923 59051
rect 265951 59023 277059 59051
rect 277087 59023 277121 59051
rect 277149 59023 281097 59051
rect 281125 59023 281159 59051
rect 281187 59023 281221 59051
rect 281249 59023 281283 59051
rect 281311 59023 296457 59051
rect 296485 59023 296519 59051
rect 296547 59023 296581 59051
rect 296609 59023 296643 59051
rect 296671 59023 298728 59051
rect 298756 59023 298790 59051
rect 298818 59023 298852 59051
rect 298880 59023 298914 59051
rect 298942 59023 298990 59051
rect -958 58989 298990 59023
rect -958 58961 -910 58989
rect -882 58961 -848 58989
rect -820 58961 -786 58989
rect -758 58961 -724 58989
rect -696 58961 4617 58989
rect 4645 58961 4679 58989
rect 4707 58961 4741 58989
rect 4769 58961 4803 58989
rect 4831 58961 15939 58989
rect 15967 58961 16001 58989
rect 16029 58961 19977 58989
rect 20005 58961 20039 58989
rect 20067 58961 20101 58989
rect 20129 58961 20163 58989
rect 20191 58961 31299 58989
rect 31327 58961 31361 58989
rect 31389 58961 35337 58989
rect 35365 58961 35399 58989
rect 35427 58961 35461 58989
rect 35489 58961 35523 58989
rect 35551 58961 46659 58989
rect 46687 58961 46721 58989
rect 46749 58961 50697 58989
rect 50725 58961 50759 58989
rect 50787 58961 50821 58989
rect 50849 58961 50883 58989
rect 50911 58961 62019 58989
rect 62047 58961 62081 58989
rect 62109 58961 66057 58989
rect 66085 58961 66119 58989
rect 66147 58961 66181 58989
rect 66209 58961 66243 58989
rect 66271 58961 77379 58989
rect 77407 58961 77441 58989
rect 77469 58961 81417 58989
rect 81445 58961 81479 58989
rect 81507 58961 81541 58989
rect 81569 58961 81603 58989
rect 81631 58961 92739 58989
rect 92767 58961 92801 58989
rect 92829 58961 96777 58989
rect 96805 58961 96839 58989
rect 96867 58961 96901 58989
rect 96929 58961 96963 58989
rect 96991 58961 108099 58989
rect 108127 58961 108161 58989
rect 108189 58961 112137 58989
rect 112165 58961 112199 58989
rect 112227 58961 112261 58989
rect 112289 58961 112323 58989
rect 112351 58961 123459 58989
rect 123487 58961 123521 58989
rect 123549 58961 127497 58989
rect 127525 58961 127559 58989
rect 127587 58961 127621 58989
rect 127649 58961 127683 58989
rect 127711 58961 138819 58989
rect 138847 58961 138881 58989
rect 138909 58961 142857 58989
rect 142885 58961 142919 58989
rect 142947 58961 142981 58989
rect 143009 58961 143043 58989
rect 143071 58961 154179 58989
rect 154207 58961 154241 58989
rect 154269 58961 158217 58989
rect 158245 58961 158279 58989
rect 158307 58961 158341 58989
rect 158369 58961 158403 58989
rect 158431 58961 169539 58989
rect 169567 58961 169601 58989
rect 169629 58961 173577 58989
rect 173605 58961 173639 58989
rect 173667 58961 173701 58989
rect 173729 58961 173763 58989
rect 173791 58961 184899 58989
rect 184927 58961 184961 58989
rect 184989 58961 188937 58989
rect 188965 58961 188999 58989
rect 189027 58961 189061 58989
rect 189089 58961 189123 58989
rect 189151 58961 200259 58989
rect 200287 58961 200321 58989
rect 200349 58961 204297 58989
rect 204325 58961 204359 58989
rect 204387 58961 204421 58989
rect 204449 58961 204483 58989
rect 204511 58961 215619 58989
rect 215647 58961 215681 58989
rect 215709 58961 219657 58989
rect 219685 58961 219719 58989
rect 219747 58961 219781 58989
rect 219809 58961 219843 58989
rect 219871 58961 230979 58989
rect 231007 58961 231041 58989
rect 231069 58961 235017 58989
rect 235045 58961 235079 58989
rect 235107 58961 235141 58989
rect 235169 58961 235203 58989
rect 235231 58961 246339 58989
rect 246367 58961 246401 58989
rect 246429 58961 250377 58989
rect 250405 58961 250439 58989
rect 250467 58961 250501 58989
rect 250529 58961 250563 58989
rect 250591 58961 261699 58989
rect 261727 58961 261761 58989
rect 261789 58961 265737 58989
rect 265765 58961 265799 58989
rect 265827 58961 265861 58989
rect 265889 58961 265923 58989
rect 265951 58961 277059 58989
rect 277087 58961 277121 58989
rect 277149 58961 281097 58989
rect 281125 58961 281159 58989
rect 281187 58961 281221 58989
rect 281249 58961 281283 58989
rect 281311 58961 296457 58989
rect 296485 58961 296519 58989
rect 296547 58961 296581 58989
rect 296609 58961 296643 58989
rect 296671 58961 298728 58989
rect 298756 58961 298790 58989
rect 298818 58961 298852 58989
rect 298880 58961 298914 58989
rect 298942 58961 298990 58989
rect -958 58913 298990 58961
rect -958 56175 298990 56223
rect -958 56147 -430 56175
rect -402 56147 -368 56175
rect -340 56147 -306 56175
rect -278 56147 -244 56175
rect -216 56147 2757 56175
rect 2785 56147 2819 56175
rect 2847 56147 2881 56175
rect 2909 56147 2943 56175
rect 2971 56147 8259 56175
rect 8287 56147 8321 56175
rect 8349 56147 18117 56175
rect 18145 56147 18179 56175
rect 18207 56147 18241 56175
rect 18269 56147 18303 56175
rect 18331 56147 23619 56175
rect 23647 56147 23681 56175
rect 23709 56147 33477 56175
rect 33505 56147 33539 56175
rect 33567 56147 33601 56175
rect 33629 56147 33663 56175
rect 33691 56147 38979 56175
rect 39007 56147 39041 56175
rect 39069 56147 48837 56175
rect 48865 56147 48899 56175
rect 48927 56147 48961 56175
rect 48989 56147 49023 56175
rect 49051 56147 54339 56175
rect 54367 56147 54401 56175
rect 54429 56147 64197 56175
rect 64225 56147 64259 56175
rect 64287 56147 64321 56175
rect 64349 56147 64383 56175
rect 64411 56147 69699 56175
rect 69727 56147 69761 56175
rect 69789 56147 79557 56175
rect 79585 56147 79619 56175
rect 79647 56147 79681 56175
rect 79709 56147 79743 56175
rect 79771 56147 85059 56175
rect 85087 56147 85121 56175
rect 85149 56147 94917 56175
rect 94945 56147 94979 56175
rect 95007 56147 95041 56175
rect 95069 56147 95103 56175
rect 95131 56147 100419 56175
rect 100447 56147 100481 56175
rect 100509 56147 110277 56175
rect 110305 56147 110339 56175
rect 110367 56147 110401 56175
rect 110429 56147 110463 56175
rect 110491 56147 115779 56175
rect 115807 56147 115841 56175
rect 115869 56147 125637 56175
rect 125665 56147 125699 56175
rect 125727 56147 125761 56175
rect 125789 56147 125823 56175
rect 125851 56147 131139 56175
rect 131167 56147 131201 56175
rect 131229 56147 140997 56175
rect 141025 56147 141059 56175
rect 141087 56147 141121 56175
rect 141149 56147 141183 56175
rect 141211 56147 146499 56175
rect 146527 56147 146561 56175
rect 146589 56147 156357 56175
rect 156385 56147 156419 56175
rect 156447 56147 156481 56175
rect 156509 56147 156543 56175
rect 156571 56147 161859 56175
rect 161887 56147 161921 56175
rect 161949 56147 171717 56175
rect 171745 56147 171779 56175
rect 171807 56147 171841 56175
rect 171869 56147 171903 56175
rect 171931 56147 177219 56175
rect 177247 56147 177281 56175
rect 177309 56147 187077 56175
rect 187105 56147 187139 56175
rect 187167 56147 187201 56175
rect 187229 56147 187263 56175
rect 187291 56147 192579 56175
rect 192607 56147 192641 56175
rect 192669 56147 202437 56175
rect 202465 56147 202499 56175
rect 202527 56147 202561 56175
rect 202589 56147 202623 56175
rect 202651 56147 207939 56175
rect 207967 56147 208001 56175
rect 208029 56147 217797 56175
rect 217825 56147 217859 56175
rect 217887 56147 217921 56175
rect 217949 56147 217983 56175
rect 218011 56147 223299 56175
rect 223327 56147 223361 56175
rect 223389 56147 233157 56175
rect 233185 56147 233219 56175
rect 233247 56147 233281 56175
rect 233309 56147 233343 56175
rect 233371 56147 238659 56175
rect 238687 56147 238721 56175
rect 238749 56147 248517 56175
rect 248545 56147 248579 56175
rect 248607 56147 248641 56175
rect 248669 56147 248703 56175
rect 248731 56147 254019 56175
rect 254047 56147 254081 56175
rect 254109 56147 263877 56175
rect 263905 56147 263939 56175
rect 263967 56147 264001 56175
rect 264029 56147 264063 56175
rect 264091 56147 269379 56175
rect 269407 56147 269441 56175
rect 269469 56147 279237 56175
rect 279265 56147 279299 56175
rect 279327 56147 279361 56175
rect 279389 56147 279423 56175
rect 279451 56147 284739 56175
rect 284767 56147 284801 56175
rect 284829 56147 294597 56175
rect 294625 56147 294659 56175
rect 294687 56147 294721 56175
rect 294749 56147 294783 56175
rect 294811 56147 298248 56175
rect 298276 56147 298310 56175
rect 298338 56147 298372 56175
rect 298400 56147 298434 56175
rect 298462 56147 298990 56175
rect -958 56113 298990 56147
rect -958 56085 -430 56113
rect -402 56085 -368 56113
rect -340 56085 -306 56113
rect -278 56085 -244 56113
rect -216 56085 2757 56113
rect 2785 56085 2819 56113
rect 2847 56085 2881 56113
rect 2909 56085 2943 56113
rect 2971 56085 8259 56113
rect 8287 56085 8321 56113
rect 8349 56085 18117 56113
rect 18145 56085 18179 56113
rect 18207 56085 18241 56113
rect 18269 56085 18303 56113
rect 18331 56085 23619 56113
rect 23647 56085 23681 56113
rect 23709 56085 33477 56113
rect 33505 56085 33539 56113
rect 33567 56085 33601 56113
rect 33629 56085 33663 56113
rect 33691 56085 38979 56113
rect 39007 56085 39041 56113
rect 39069 56085 48837 56113
rect 48865 56085 48899 56113
rect 48927 56085 48961 56113
rect 48989 56085 49023 56113
rect 49051 56085 54339 56113
rect 54367 56085 54401 56113
rect 54429 56085 64197 56113
rect 64225 56085 64259 56113
rect 64287 56085 64321 56113
rect 64349 56085 64383 56113
rect 64411 56085 69699 56113
rect 69727 56085 69761 56113
rect 69789 56085 79557 56113
rect 79585 56085 79619 56113
rect 79647 56085 79681 56113
rect 79709 56085 79743 56113
rect 79771 56085 85059 56113
rect 85087 56085 85121 56113
rect 85149 56085 94917 56113
rect 94945 56085 94979 56113
rect 95007 56085 95041 56113
rect 95069 56085 95103 56113
rect 95131 56085 100419 56113
rect 100447 56085 100481 56113
rect 100509 56085 110277 56113
rect 110305 56085 110339 56113
rect 110367 56085 110401 56113
rect 110429 56085 110463 56113
rect 110491 56085 115779 56113
rect 115807 56085 115841 56113
rect 115869 56085 125637 56113
rect 125665 56085 125699 56113
rect 125727 56085 125761 56113
rect 125789 56085 125823 56113
rect 125851 56085 131139 56113
rect 131167 56085 131201 56113
rect 131229 56085 140997 56113
rect 141025 56085 141059 56113
rect 141087 56085 141121 56113
rect 141149 56085 141183 56113
rect 141211 56085 146499 56113
rect 146527 56085 146561 56113
rect 146589 56085 156357 56113
rect 156385 56085 156419 56113
rect 156447 56085 156481 56113
rect 156509 56085 156543 56113
rect 156571 56085 161859 56113
rect 161887 56085 161921 56113
rect 161949 56085 171717 56113
rect 171745 56085 171779 56113
rect 171807 56085 171841 56113
rect 171869 56085 171903 56113
rect 171931 56085 177219 56113
rect 177247 56085 177281 56113
rect 177309 56085 187077 56113
rect 187105 56085 187139 56113
rect 187167 56085 187201 56113
rect 187229 56085 187263 56113
rect 187291 56085 192579 56113
rect 192607 56085 192641 56113
rect 192669 56085 202437 56113
rect 202465 56085 202499 56113
rect 202527 56085 202561 56113
rect 202589 56085 202623 56113
rect 202651 56085 207939 56113
rect 207967 56085 208001 56113
rect 208029 56085 217797 56113
rect 217825 56085 217859 56113
rect 217887 56085 217921 56113
rect 217949 56085 217983 56113
rect 218011 56085 223299 56113
rect 223327 56085 223361 56113
rect 223389 56085 233157 56113
rect 233185 56085 233219 56113
rect 233247 56085 233281 56113
rect 233309 56085 233343 56113
rect 233371 56085 238659 56113
rect 238687 56085 238721 56113
rect 238749 56085 248517 56113
rect 248545 56085 248579 56113
rect 248607 56085 248641 56113
rect 248669 56085 248703 56113
rect 248731 56085 254019 56113
rect 254047 56085 254081 56113
rect 254109 56085 263877 56113
rect 263905 56085 263939 56113
rect 263967 56085 264001 56113
rect 264029 56085 264063 56113
rect 264091 56085 269379 56113
rect 269407 56085 269441 56113
rect 269469 56085 279237 56113
rect 279265 56085 279299 56113
rect 279327 56085 279361 56113
rect 279389 56085 279423 56113
rect 279451 56085 284739 56113
rect 284767 56085 284801 56113
rect 284829 56085 294597 56113
rect 294625 56085 294659 56113
rect 294687 56085 294721 56113
rect 294749 56085 294783 56113
rect 294811 56085 298248 56113
rect 298276 56085 298310 56113
rect 298338 56085 298372 56113
rect 298400 56085 298434 56113
rect 298462 56085 298990 56113
rect -958 56051 298990 56085
rect -958 56023 -430 56051
rect -402 56023 -368 56051
rect -340 56023 -306 56051
rect -278 56023 -244 56051
rect -216 56023 2757 56051
rect 2785 56023 2819 56051
rect 2847 56023 2881 56051
rect 2909 56023 2943 56051
rect 2971 56023 8259 56051
rect 8287 56023 8321 56051
rect 8349 56023 18117 56051
rect 18145 56023 18179 56051
rect 18207 56023 18241 56051
rect 18269 56023 18303 56051
rect 18331 56023 23619 56051
rect 23647 56023 23681 56051
rect 23709 56023 33477 56051
rect 33505 56023 33539 56051
rect 33567 56023 33601 56051
rect 33629 56023 33663 56051
rect 33691 56023 38979 56051
rect 39007 56023 39041 56051
rect 39069 56023 48837 56051
rect 48865 56023 48899 56051
rect 48927 56023 48961 56051
rect 48989 56023 49023 56051
rect 49051 56023 54339 56051
rect 54367 56023 54401 56051
rect 54429 56023 64197 56051
rect 64225 56023 64259 56051
rect 64287 56023 64321 56051
rect 64349 56023 64383 56051
rect 64411 56023 69699 56051
rect 69727 56023 69761 56051
rect 69789 56023 79557 56051
rect 79585 56023 79619 56051
rect 79647 56023 79681 56051
rect 79709 56023 79743 56051
rect 79771 56023 85059 56051
rect 85087 56023 85121 56051
rect 85149 56023 94917 56051
rect 94945 56023 94979 56051
rect 95007 56023 95041 56051
rect 95069 56023 95103 56051
rect 95131 56023 100419 56051
rect 100447 56023 100481 56051
rect 100509 56023 110277 56051
rect 110305 56023 110339 56051
rect 110367 56023 110401 56051
rect 110429 56023 110463 56051
rect 110491 56023 115779 56051
rect 115807 56023 115841 56051
rect 115869 56023 125637 56051
rect 125665 56023 125699 56051
rect 125727 56023 125761 56051
rect 125789 56023 125823 56051
rect 125851 56023 131139 56051
rect 131167 56023 131201 56051
rect 131229 56023 140997 56051
rect 141025 56023 141059 56051
rect 141087 56023 141121 56051
rect 141149 56023 141183 56051
rect 141211 56023 146499 56051
rect 146527 56023 146561 56051
rect 146589 56023 156357 56051
rect 156385 56023 156419 56051
rect 156447 56023 156481 56051
rect 156509 56023 156543 56051
rect 156571 56023 161859 56051
rect 161887 56023 161921 56051
rect 161949 56023 171717 56051
rect 171745 56023 171779 56051
rect 171807 56023 171841 56051
rect 171869 56023 171903 56051
rect 171931 56023 177219 56051
rect 177247 56023 177281 56051
rect 177309 56023 187077 56051
rect 187105 56023 187139 56051
rect 187167 56023 187201 56051
rect 187229 56023 187263 56051
rect 187291 56023 192579 56051
rect 192607 56023 192641 56051
rect 192669 56023 202437 56051
rect 202465 56023 202499 56051
rect 202527 56023 202561 56051
rect 202589 56023 202623 56051
rect 202651 56023 207939 56051
rect 207967 56023 208001 56051
rect 208029 56023 217797 56051
rect 217825 56023 217859 56051
rect 217887 56023 217921 56051
rect 217949 56023 217983 56051
rect 218011 56023 223299 56051
rect 223327 56023 223361 56051
rect 223389 56023 233157 56051
rect 233185 56023 233219 56051
rect 233247 56023 233281 56051
rect 233309 56023 233343 56051
rect 233371 56023 238659 56051
rect 238687 56023 238721 56051
rect 238749 56023 248517 56051
rect 248545 56023 248579 56051
rect 248607 56023 248641 56051
rect 248669 56023 248703 56051
rect 248731 56023 254019 56051
rect 254047 56023 254081 56051
rect 254109 56023 263877 56051
rect 263905 56023 263939 56051
rect 263967 56023 264001 56051
rect 264029 56023 264063 56051
rect 264091 56023 269379 56051
rect 269407 56023 269441 56051
rect 269469 56023 279237 56051
rect 279265 56023 279299 56051
rect 279327 56023 279361 56051
rect 279389 56023 279423 56051
rect 279451 56023 284739 56051
rect 284767 56023 284801 56051
rect 284829 56023 294597 56051
rect 294625 56023 294659 56051
rect 294687 56023 294721 56051
rect 294749 56023 294783 56051
rect 294811 56023 298248 56051
rect 298276 56023 298310 56051
rect 298338 56023 298372 56051
rect 298400 56023 298434 56051
rect 298462 56023 298990 56051
rect -958 55989 298990 56023
rect -958 55961 -430 55989
rect -402 55961 -368 55989
rect -340 55961 -306 55989
rect -278 55961 -244 55989
rect -216 55961 2757 55989
rect 2785 55961 2819 55989
rect 2847 55961 2881 55989
rect 2909 55961 2943 55989
rect 2971 55961 8259 55989
rect 8287 55961 8321 55989
rect 8349 55961 18117 55989
rect 18145 55961 18179 55989
rect 18207 55961 18241 55989
rect 18269 55961 18303 55989
rect 18331 55961 23619 55989
rect 23647 55961 23681 55989
rect 23709 55961 33477 55989
rect 33505 55961 33539 55989
rect 33567 55961 33601 55989
rect 33629 55961 33663 55989
rect 33691 55961 38979 55989
rect 39007 55961 39041 55989
rect 39069 55961 48837 55989
rect 48865 55961 48899 55989
rect 48927 55961 48961 55989
rect 48989 55961 49023 55989
rect 49051 55961 54339 55989
rect 54367 55961 54401 55989
rect 54429 55961 64197 55989
rect 64225 55961 64259 55989
rect 64287 55961 64321 55989
rect 64349 55961 64383 55989
rect 64411 55961 69699 55989
rect 69727 55961 69761 55989
rect 69789 55961 79557 55989
rect 79585 55961 79619 55989
rect 79647 55961 79681 55989
rect 79709 55961 79743 55989
rect 79771 55961 85059 55989
rect 85087 55961 85121 55989
rect 85149 55961 94917 55989
rect 94945 55961 94979 55989
rect 95007 55961 95041 55989
rect 95069 55961 95103 55989
rect 95131 55961 100419 55989
rect 100447 55961 100481 55989
rect 100509 55961 110277 55989
rect 110305 55961 110339 55989
rect 110367 55961 110401 55989
rect 110429 55961 110463 55989
rect 110491 55961 115779 55989
rect 115807 55961 115841 55989
rect 115869 55961 125637 55989
rect 125665 55961 125699 55989
rect 125727 55961 125761 55989
rect 125789 55961 125823 55989
rect 125851 55961 131139 55989
rect 131167 55961 131201 55989
rect 131229 55961 140997 55989
rect 141025 55961 141059 55989
rect 141087 55961 141121 55989
rect 141149 55961 141183 55989
rect 141211 55961 146499 55989
rect 146527 55961 146561 55989
rect 146589 55961 156357 55989
rect 156385 55961 156419 55989
rect 156447 55961 156481 55989
rect 156509 55961 156543 55989
rect 156571 55961 161859 55989
rect 161887 55961 161921 55989
rect 161949 55961 171717 55989
rect 171745 55961 171779 55989
rect 171807 55961 171841 55989
rect 171869 55961 171903 55989
rect 171931 55961 177219 55989
rect 177247 55961 177281 55989
rect 177309 55961 187077 55989
rect 187105 55961 187139 55989
rect 187167 55961 187201 55989
rect 187229 55961 187263 55989
rect 187291 55961 192579 55989
rect 192607 55961 192641 55989
rect 192669 55961 202437 55989
rect 202465 55961 202499 55989
rect 202527 55961 202561 55989
rect 202589 55961 202623 55989
rect 202651 55961 207939 55989
rect 207967 55961 208001 55989
rect 208029 55961 217797 55989
rect 217825 55961 217859 55989
rect 217887 55961 217921 55989
rect 217949 55961 217983 55989
rect 218011 55961 223299 55989
rect 223327 55961 223361 55989
rect 223389 55961 233157 55989
rect 233185 55961 233219 55989
rect 233247 55961 233281 55989
rect 233309 55961 233343 55989
rect 233371 55961 238659 55989
rect 238687 55961 238721 55989
rect 238749 55961 248517 55989
rect 248545 55961 248579 55989
rect 248607 55961 248641 55989
rect 248669 55961 248703 55989
rect 248731 55961 254019 55989
rect 254047 55961 254081 55989
rect 254109 55961 263877 55989
rect 263905 55961 263939 55989
rect 263967 55961 264001 55989
rect 264029 55961 264063 55989
rect 264091 55961 269379 55989
rect 269407 55961 269441 55989
rect 269469 55961 279237 55989
rect 279265 55961 279299 55989
rect 279327 55961 279361 55989
rect 279389 55961 279423 55989
rect 279451 55961 284739 55989
rect 284767 55961 284801 55989
rect 284829 55961 294597 55989
rect 294625 55961 294659 55989
rect 294687 55961 294721 55989
rect 294749 55961 294783 55989
rect 294811 55961 298248 55989
rect 298276 55961 298310 55989
rect 298338 55961 298372 55989
rect 298400 55961 298434 55989
rect 298462 55961 298990 55989
rect -958 55913 298990 55961
rect -958 50175 298990 50223
rect -958 50147 -910 50175
rect -882 50147 -848 50175
rect -820 50147 -786 50175
rect -758 50147 -724 50175
rect -696 50147 4617 50175
rect 4645 50147 4679 50175
rect 4707 50147 4741 50175
rect 4769 50147 4803 50175
rect 4831 50147 15939 50175
rect 15967 50147 16001 50175
rect 16029 50147 19977 50175
rect 20005 50147 20039 50175
rect 20067 50147 20101 50175
rect 20129 50147 20163 50175
rect 20191 50147 31299 50175
rect 31327 50147 31361 50175
rect 31389 50147 35337 50175
rect 35365 50147 35399 50175
rect 35427 50147 35461 50175
rect 35489 50147 35523 50175
rect 35551 50147 46659 50175
rect 46687 50147 46721 50175
rect 46749 50147 50697 50175
rect 50725 50147 50759 50175
rect 50787 50147 50821 50175
rect 50849 50147 50883 50175
rect 50911 50147 62019 50175
rect 62047 50147 62081 50175
rect 62109 50147 66057 50175
rect 66085 50147 66119 50175
rect 66147 50147 66181 50175
rect 66209 50147 66243 50175
rect 66271 50147 77379 50175
rect 77407 50147 77441 50175
rect 77469 50147 81417 50175
rect 81445 50147 81479 50175
rect 81507 50147 81541 50175
rect 81569 50147 81603 50175
rect 81631 50147 92739 50175
rect 92767 50147 92801 50175
rect 92829 50147 96777 50175
rect 96805 50147 96839 50175
rect 96867 50147 96901 50175
rect 96929 50147 96963 50175
rect 96991 50147 108099 50175
rect 108127 50147 108161 50175
rect 108189 50147 112137 50175
rect 112165 50147 112199 50175
rect 112227 50147 112261 50175
rect 112289 50147 112323 50175
rect 112351 50147 123459 50175
rect 123487 50147 123521 50175
rect 123549 50147 127497 50175
rect 127525 50147 127559 50175
rect 127587 50147 127621 50175
rect 127649 50147 127683 50175
rect 127711 50147 138819 50175
rect 138847 50147 138881 50175
rect 138909 50147 142857 50175
rect 142885 50147 142919 50175
rect 142947 50147 142981 50175
rect 143009 50147 143043 50175
rect 143071 50147 154179 50175
rect 154207 50147 154241 50175
rect 154269 50147 158217 50175
rect 158245 50147 158279 50175
rect 158307 50147 158341 50175
rect 158369 50147 158403 50175
rect 158431 50147 169539 50175
rect 169567 50147 169601 50175
rect 169629 50147 173577 50175
rect 173605 50147 173639 50175
rect 173667 50147 173701 50175
rect 173729 50147 173763 50175
rect 173791 50147 184899 50175
rect 184927 50147 184961 50175
rect 184989 50147 188937 50175
rect 188965 50147 188999 50175
rect 189027 50147 189061 50175
rect 189089 50147 189123 50175
rect 189151 50147 200259 50175
rect 200287 50147 200321 50175
rect 200349 50147 204297 50175
rect 204325 50147 204359 50175
rect 204387 50147 204421 50175
rect 204449 50147 204483 50175
rect 204511 50147 215619 50175
rect 215647 50147 215681 50175
rect 215709 50147 219657 50175
rect 219685 50147 219719 50175
rect 219747 50147 219781 50175
rect 219809 50147 219843 50175
rect 219871 50147 230979 50175
rect 231007 50147 231041 50175
rect 231069 50147 235017 50175
rect 235045 50147 235079 50175
rect 235107 50147 235141 50175
rect 235169 50147 235203 50175
rect 235231 50147 246339 50175
rect 246367 50147 246401 50175
rect 246429 50147 250377 50175
rect 250405 50147 250439 50175
rect 250467 50147 250501 50175
rect 250529 50147 250563 50175
rect 250591 50147 261699 50175
rect 261727 50147 261761 50175
rect 261789 50147 265737 50175
rect 265765 50147 265799 50175
rect 265827 50147 265861 50175
rect 265889 50147 265923 50175
rect 265951 50147 277059 50175
rect 277087 50147 277121 50175
rect 277149 50147 281097 50175
rect 281125 50147 281159 50175
rect 281187 50147 281221 50175
rect 281249 50147 281283 50175
rect 281311 50147 296457 50175
rect 296485 50147 296519 50175
rect 296547 50147 296581 50175
rect 296609 50147 296643 50175
rect 296671 50147 298728 50175
rect 298756 50147 298790 50175
rect 298818 50147 298852 50175
rect 298880 50147 298914 50175
rect 298942 50147 298990 50175
rect -958 50113 298990 50147
rect -958 50085 -910 50113
rect -882 50085 -848 50113
rect -820 50085 -786 50113
rect -758 50085 -724 50113
rect -696 50085 4617 50113
rect 4645 50085 4679 50113
rect 4707 50085 4741 50113
rect 4769 50085 4803 50113
rect 4831 50085 15939 50113
rect 15967 50085 16001 50113
rect 16029 50085 19977 50113
rect 20005 50085 20039 50113
rect 20067 50085 20101 50113
rect 20129 50085 20163 50113
rect 20191 50085 31299 50113
rect 31327 50085 31361 50113
rect 31389 50085 35337 50113
rect 35365 50085 35399 50113
rect 35427 50085 35461 50113
rect 35489 50085 35523 50113
rect 35551 50085 46659 50113
rect 46687 50085 46721 50113
rect 46749 50085 50697 50113
rect 50725 50085 50759 50113
rect 50787 50085 50821 50113
rect 50849 50085 50883 50113
rect 50911 50085 62019 50113
rect 62047 50085 62081 50113
rect 62109 50085 66057 50113
rect 66085 50085 66119 50113
rect 66147 50085 66181 50113
rect 66209 50085 66243 50113
rect 66271 50085 77379 50113
rect 77407 50085 77441 50113
rect 77469 50085 81417 50113
rect 81445 50085 81479 50113
rect 81507 50085 81541 50113
rect 81569 50085 81603 50113
rect 81631 50085 92739 50113
rect 92767 50085 92801 50113
rect 92829 50085 96777 50113
rect 96805 50085 96839 50113
rect 96867 50085 96901 50113
rect 96929 50085 96963 50113
rect 96991 50085 108099 50113
rect 108127 50085 108161 50113
rect 108189 50085 112137 50113
rect 112165 50085 112199 50113
rect 112227 50085 112261 50113
rect 112289 50085 112323 50113
rect 112351 50085 123459 50113
rect 123487 50085 123521 50113
rect 123549 50085 127497 50113
rect 127525 50085 127559 50113
rect 127587 50085 127621 50113
rect 127649 50085 127683 50113
rect 127711 50085 138819 50113
rect 138847 50085 138881 50113
rect 138909 50085 142857 50113
rect 142885 50085 142919 50113
rect 142947 50085 142981 50113
rect 143009 50085 143043 50113
rect 143071 50085 154179 50113
rect 154207 50085 154241 50113
rect 154269 50085 158217 50113
rect 158245 50085 158279 50113
rect 158307 50085 158341 50113
rect 158369 50085 158403 50113
rect 158431 50085 169539 50113
rect 169567 50085 169601 50113
rect 169629 50085 173577 50113
rect 173605 50085 173639 50113
rect 173667 50085 173701 50113
rect 173729 50085 173763 50113
rect 173791 50085 184899 50113
rect 184927 50085 184961 50113
rect 184989 50085 188937 50113
rect 188965 50085 188999 50113
rect 189027 50085 189061 50113
rect 189089 50085 189123 50113
rect 189151 50085 200259 50113
rect 200287 50085 200321 50113
rect 200349 50085 204297 50113
rect 204325 50085 204359 50113
rect 204387 50085 204421 50113
rect 204449 50085 204483 50113
rect 204511 50085 215619 50113
rect 215647 50085 215681 50113
rect 215709 50085 219657 50113
rect 219685 50085 219719 50113
rect 219747 50085 219781 50113
rect 219809 50085 219843 50113
rect 219871 50085 230979 50113
rect 231007 50085 231041 50113
rect 231069 50085 235017 50113
rect 235045 50085 235079 50113
rect 235107 50085 235141 50113
rect 235169 50085 235203 50113
rect 235231 50085 246339 50113
rect 246367 50085 246401 50113
rect 246429 50085 250377 50113
rect 250405 50085 250439 50113
rect 250467 50085 250501 50113
rect 250529 50085 250563 50113
rect 250591 50085 261699 50113
rect 261727 50085 261761 50113
rect 261789 50085 265737 50113
rect 265765 50085 265799 50113
rect 265827 50085 265861 50113
rect 265889 50085 265923 50113
rect 265951 50085 277059 50113
rect 277087 50085 277121 50113
rect 277149 50085 281097 50113
rect 281125 50085 281159 50113
rect 281187 50085 281221 50113
rect 281249 50085 281283 50113
rect 281311 50085 296457 50113
rect 296485 50085 296519 50113
rect 296547 50085 296581 50113
rect 296609 50085 296643 50113
rect 296671 50085 298728 50113
rect 298756 50085 298790 50113
rect 298818 50085 298852 50113
rect 298880 50085 298914 50113
rect 298942 50085 298990 50113
rect -958 50051 298990 50085
rect -958 50023 -910 50051
rect -882 50023 -848 50051
rect -820 50023 -786 50051
rect -758 50023 -724 50051
rect -696 50023 4617 50051
rect 4645 50023 4679 50051
rect 4707 50023 4741 50051
rect 4769 50023 4803 50051
rect 4831 50023 15939 50051
rect 15967 50023 16001 50051
rect 16029 50023 19977 50051
rect 20005 50023 20039 50051
rect 20067 50023 20101 50051
rect 20129 50023 20163 50051
rect 20191 50023 31299 50051
rect 31327 50023 31361 50051
rect 31389 50023 35337 50051
rect 35365 50023 35399 50051
rect 35427 50023 35461 50051
rect 35489 50023 35523 50051
rect 35551 50023 46659 50051
rect 46687 50023 46721 50051
rect 46749 50023 50697 50051
rect 50725 50023 50759 50051
rect 50787 50023 50821 50051
rect 50849 50023 50883 50051
rect 50911 50023 62019 50051
rect 62047 50023 62081 50051
rect 62109 50023 66057 50051
rect 66085 50023 66119 50051
rect 66147 50023 66181 50051
rect 66209 50023 66243 50051
rect 66271 50023 77379 50051
rect 77407 50023 77441 50051
rect 77469 50023 81417 50051
rect 81445 50023 81479 50051
rect 81507 50023 81541 50051
rect 81569 50023 81603 50051
rect 81631 50023 92739 50051
rect 92767 50023 92801 50051
rect 92829 50023 96777 50051
rect 96805 50023 96839 50051
rect 96867 50023 96901 50051
rect 96929 50023 96963 50051
rect 96991 50023 108099 50051
rect 108127 50023 108161 50051
rect 108189 50023 112137 50051
rect 112165 50023 112199 50051
rect 112227 50023 112261 50051
rect 112289 50023 112323 50051
rect 112351 50023 123459 50051
rect 123487 50023 123521 50051
rect 123549 50023 127497 50051
rect 127525 50023 127559 50051
rect 127587 50023 127621 50051
rect 127649 50023 127683 50051
rect 127711 50023 138819 50051
rect 138847 50023 138881 50051
rect 138909 50023 142857 50051
rect 142885 50023 142919 50051
rect 142947 50023 142981 50051
rect 143009 50023 143043 50051
rect 143071 50023 154179 50051
rect 154207 50023 154241 50051
rect 154269 50023 158217 50051
rect 158245 50023 158279 50051
rect 158307 50023 158341 50051
rect 158369 50023 158403 50051
rect 158431 50023 169539 50051
rect 169567 50023 169601 50051
rect 169629 50023 173577 50051
rect 173605 50023 173639 50051
rect 173667 50023 173701 50051
rect 173729 50023 173763 50051
rect 173791 50023 184899 50051
rect 184927 50023 184961 50051
rect 184989 50023 188937 50051
rect 188965 50023 188999 50051
rect 189027 50023 189061 50051
rect 189089 50023 189123 50051
rect 189151 50023 200259 50051
rect 200287 50023 200321 50051
rect 200349 50023 204297 50051
rect 204325 50023 204359 50051
rect 204387 50023 204421 50051
rect 204449 50023 204483 50051
rect 204511 50023 215619 50051
rect 215647 50023 215681 50051
rect 215709 50023 219657 50051
rect 219685 50023 219719 50051
rect 219747 50023 219781 50051
rect 219809 50023 219843 50051
rect 219871 50023 230979 50051
rect 231007 50023 231041 50051
rect 231069 50023 235017 50051
rect 235045 50023 235079 50051
rect 235107 50023 235141 50051
rect 235169 50023 235203 50051
rect 235231 50023 246339 50051
rect 246367 50023 246401 50051
rect 246429 50023 250377 50051
rect 250405 50023 250439 50051
rect 250467 50023 250501 50051
rect 250529 50023 250563 50051
rect 250591 50023 261699 50051
rect 261727 50023 261761 50051
rect 261789 50023 265737 50051
rect 265765 50023 265799 50051
rect 265827 50023 265861 50051
rect 265889 50023 265923 50051
rect 265951 50023 277059 50051
rect 277087 50023 277121 50051
rect 277149 50023 281097 50051
rect 281125 50023 281159 50051
rect 281187 50023 281221 50051
rect 281249 50023 281283 50051
rect 281311 50023 296457 50051
rect 296485 50023 296519 50051
rect 296547 50023 296581 50051
rect 296609 50023 296643 50051
rect 296671 50023 298728 50051
rect 298756 50023 298790 50051
rect 298818 50023 298852 50051
rect 298880 50023 298914 50051
rect 298942 50023 298990 50051
rect -958 49989 298990 50023
rect -958 49961 -910 49989
rect -882 49961 -848 49989
rect -820 49961 -786 49989
rect -758 49961 -724 49989
rect -696 49961 4617 49989
rect 4645 49961 4679 49989
rect 4707 49961 4741 49989
rect 4769 49961 4803 49989
rect 4831 49961 15939 49989
rect 15967 49961 16001 49989
rect 16029 49961 19977 49989
rect 20005 49961 20039 49989
rect 20067 49961 20101 49989
rect 20129 49961 20163 49989
rect 20191 49961 31299 49989
rect 31327 49961 31361 49989
rect 31389 49961 35337 49989
rect 35365 49961 35399 49989
rect 35427 49961 35461 49989
rect 35489 49961 35523 49989
rect 35551 49961 46659 49989
rect 46687 49961 46721 49989
rect 46749 49961 50697 49989
rect 50725 49961 50759 49989
rect 50787 49961 50821 49989
rect 50849 49961 50883 49989
rect 50911 49961 62019 49989
rect 62047 49961 62081 49989
rect 62109 49961 66057 49989
rect 66085 49961 66119 49989
rect 66147 49961 66181 49989
rect 66209 49961 66243 49989
rect 66271 49961 77379 49989
rect 77407 49961 77441 49989
rect 77469 49961 81417 49989
rect 81445 49961 81479 49989
rect 81507 49961 81541 49989
rect 81569 49961 81603 49989
rect 81631 49961 92739 49989
rect 92767 49961 92801 49989
rect 92829 49961 96777 49989
rect 96805 49961 96839 49989
rect 96867 49961 96901 49989
rect 96929 49961 96963 49989
rect 96991 49961 108099 49989
rect 108127 49961 108161 49989
rect 108189 49961 112137 49989
rect 112165 49961 112199 49989
rect 112227 49961 112261 49989
rect 112289 49961 112323 49989
rect 112351 49961 123459 49989
rect 123487 49961 123521 49989
rect 123549 49961 127497 49989
rect 127525 49961 127559 49989
rect 127587 49961 127621 49989
rect 127649 49961 127683 49989
rect 127711 49961 138819 49989
rect 138847 49961 138881 49989
rect 138909 49961 142857 49989
rect 142885 49961 142919 49989
rect 142947 49961 142981 49989
rect 143009 49961 143043 49989
rect 143071 49961 154179 49989
rect 154207 49961 154241 49989
rect 154269 49961 158217 49989
rect 158245 49961 158279 49989
rect 158307 49961 158341 49989
rect 158369 49961 158403 49989
rect 158431 49961 169539 49989
rect 169567 49961 169601 49989
rect 169629 49961 173577 49989
rect 173605 49961 173639 49989
rect 173667 49961 173701 49989
rect 173729 49961 173763 49989
rect 173791 49961 184899 49989
rect 184927 49961 184961 49989
rect 184989 49961 188937 49989
rect 188965 49961 188999 49989
rect 189027 49961 189061 49989
rect 189089 49961 189123 49989
rect 189151 49961 200259 49989
rect 200287 49961 200321 49989
rect 200349 49961 204297 49989
rect 204325 49961 204359 49989
rect 204387 49961 204421 49989
rect 204449 49961 204483 49989
rect 204511 49961 215619 49989
rect 215647 49961 215681 49989
rect 215709 49961 219657 49989
rect 219685 49961 219719 49989
rect 219747 49961 219781 49989
rect 219809 49961 219843 49989
rect 219871 49961 230979 49989
rect 231007 49961 231041 49989
rect 231069 49961 235017 49989
rect 235045 49961 235079 49989
rect 235107 49961 235141 49989
rect 235169 49961 235203 49989
rect 235231 49961 246339 49989
rect 246367 49961 246401 49989
rect 246429 49961 250377 49989
rect 250405 49961 250439 49989
rect 250467 49961 250501 49989
rect 250529 49961 250563 49989
rect 250591 49961 261699 49989
rect 261727 49961 261761 49989
rect 261789 49961 265737 49989
rect 265765 49961 265799 49989
rect 265827 49961 265861 49989
rect 265889 49961 265923 49989
rect 265951 49961 277059 49989
rect 277087 49961 277121 49989
rect 277149 49961 281097 49989
rect 281125 49961 281159 49989
rect 281187 49961 281221 49989
rect 281249 49961 281283 49989
rect 281311 49961 296457 49989
rect 296485 49961 296519 49989
rect 296547 49961 296581 49989
rect 296609 49961 296643 49989
rect 296671 49961 298728 49989
rect 298756 49961 298790 49989
rect 298818 49961 298852 49989
rect 298880 49961 298914 49989
rect 298942 49961 298990 49989
rect -958 49913 298990 49961
rect -958 47175 298990 47223
rect -958 47147 -430 47175
rect -402 47147 -368 47175
rect -340 47147 -306 47175
rect -278 47147 -244 47175
rect -216 47147 2757 47175
rect 2785 47147 2819 47175
rect 2847 47147 2881 47175
rect 2909 47147 2943 47175
rect 2971 47147 8259 47175
rect 8287 47147 8321 47175
rect 8349 47147 18117 47175
rect 18145 47147 18179 47175
rect 18207 47147 18241 47175
rect 18269 47147 18303 47175
rect 18331 47147 23619 47175
rect 23647 47147 23681 47175
rect 23709 47147 33477 47175
rect 33505 47147 33539 47175
rect 33567 47147 33601 47175
rect 33629 47147 33663 47175
rect 33691 47147 38979 47175
rect 39007 47147 39041 47175
rect 39069 47147 48837 47175
rect 48865 47147 48899 47175
rect 48927 47147 48961 47175
rect 48989 47147 49023 47175
rect 49051 47147 54339 47175
rect 54367 47147 54401 47175
rect 54429 47147 64197 47175
rect 64225 47147 64259 47175
rect 64287 47147 64321 47175
rect 64349 47147 64383 47175
rect 64411 47147 69699 47175
rect 69727 47147 69761 47175
rect 69789 47147 79557 47175
rect 79585 47147 79619 47175
rect 79647 47147 79681 47175
rect 79709 47147 79743 47175
rect 79771 47147 85059 47175
rect 85087 47147 85121 47175
rect 85149 47147 94917 47175
rect 94945 47147 94979 47175
rect 95007 47147 95041 47175
rect 95069 47147 95103 47175
rect 95131 47147 100419 47175
rect 100447 47147 100481 47175
rect 100509 47147 110277 47175
rect 110305 47147 110339 47175
rect 110367 47147 110401 47175
rect 110429 47147 110463 47175
rect 110491 47147 115779 47175
rect 115807 47147 115841 47175
rect 115869 47147 125637 47175
rect 125665 47147 125699 47175
rect 125727 47147 125761 47175
rect 125789 47147 125823 47175
rect 125851 47147 131139 47175
rect 131167 47147 131201 47175
rect 131229 47147 140997 47175
rect 141025 47147 141059 47175
rect 141087 47147 141121 47175
rect 141149 47147 141183 47175
rect 141211 47147 146499 47175
rect 146527 47147 146561 47175
rect 146589 47147 156357 47175
rect 156385 47147 156419 47175
rect 156447 47147 156481 47175
rect 156509 47147 156543 47175
rect 156571 47147 161859 47175
rect 161887 47147 161921 47175
rect 161949 47147 171717 47175
rect 171745 47147 171779 47175
rect 171807 47147 171841 47175
rect 171869 47147 171903 47175
rect 171931 47147 177219 47175
rect 177247 47147 177281 47175
rect 177309 47147 187077 47175
rect 187105 47147 187139 47175
rect 187167 47147 187201 47175
rect 187229 47147 187263 47175
rect 187291 47147 192579 47175
rect 192607 47147 192641 47175
rect 192669 47147 202437 47175
rect 202465 47147 202499 47175
rect 202527 47147 202561 47175
rect 202589 47147 202623 47175
rect 202651 47147 207939 47175
rect 207967 47147 208001 47175
rect 208029 47147 217797 47175
rect 217825 47147 217859 47175
rect 217887 47147 217921 47175
rect 217949 47147 217983 47175
rect 218011 47147 223299 47175
rect 223327 47147 223361 47175
rect 223389 47147 233157 47175
rect 233185 47147 233219 47175
rect 233247 47147 233281 47175
rect 233309 47147 233343 47175
rect 233371 47147 238659 47175
rect 238687 47147 238721 47175
rect 238749 47147 248517 47175
rect 248545 47147 248579 47175
rect 248607 47147 248641 47175
rect 248669 47147 248703 47175
rect 248731 47147 254019 47175
rect 254047 47147 254081 47175
rect 254109 47147 263877 47175
rect 263905 47147 263939 47175
rect 263967 47147 264001 47175
rect 264029 47147 264063 47175
rect 264091 47147 269379 47175
rect 269407 47147 269441 47175
rect 269469 47147 279237 47175
rect 279265 47147 279299 47175
rect 279327 47147 279361 47175
rect 279389 47147 279423 47175
rect 279451 47147 284739 47175
rect 284767 47147 284801 47175
rect 284829 47147 294597 47175
rect 294625 47147 294659 47175
rect 294687 47147 294721 47175
rect 294749 47147 294783 47175
rect 294811 47147 298248 47175
rect 298276 47147 298310 47175
rect 298338 47147 298372 47175
rect 298400 47147 298434 47175
rect 298462 47147 298990 47175
rect -958 47113 298990 47147
rect -958 47085 -430 47113
rect -402 47085 -368 47113
rect -340 47085 -306 47113
rect -278 47085 -244 47113
rect -216 47085 2757 47113
rect 2785 47085 2819 47113
rect 2847 47085 2881 47113
rect 2909 47085 2943 47113
rect 2971 47085 8259 47113
rect 8287 47085 8321 47113
rect 8349 47085 18117 47113
rect 18145 47085 18179 47113
rect 18207 47085 18241 47113
rect 18269 47085 18303 47113
rect 18331 47085 23619 47113
rect 23647 47085 23681 47113
rect 23709 47085 33477 47113
rect 33505 47085 33539 47113
rect 33567 47085 33601 47113
rect 33629 47085 33663 47113
rect 33691 47085 38979 47113
rect 39007 47085 39041 47113
rect 39069 47085 48837 47113
rect 48865 47085 48899 47113
rect 48927 47085 48961 47113
rect 48989 47085 49023 47113
rect 49051 47085 54339 47113
rect 54367 47085 54401 47113
rect 54429 47085 64197 47113
rect 64225 47085 64259 47113
rect 64287 47085 64321 47113
rect 64349 47085 64383 47113
rect 64411 47085 69699 47113
rect 69727 47085 69761 47113
rect 69789 47085 79557 47113
rect 79585 47085 79619 47113
rect 79647 47085 79681 47113
rect 79709 47085 79743 47113
rect 79771 47085 85059 47113
rect 85087 47085 85121 47113
rect 85149 47085 94917 47113
rect 94945 47085 94979 47113
rect 95007 47085 95041 47113
rect 95069 47085 95103 47113
rect 95131 47085 100419 47113
rect 100447 47085 100481 47113
rect 100509 47085 110277 47113
rect 110305 47085 110339 47113
rect 110367 47085 110401 47113
rect 110429 47085 110463 47113
rect 110491 47085 115779 47113
rect 115807 47085 115841 47113
rect 115869 47085 125637 47113
rect 125665 47085 125699 47113
rect 125727 47085 125761 47113
rect 125789 47085 125823 47113
rect 125851 47085 131139 47113
rect 131167 47085 131201 47113
rect 131229 47085 140997 47113
rect 141025 47085 141059 47113
rect 141087 47085 141121 47113
rect 141149 47085 141183 47113
rect 141211 47085 146499 47113
rect 146527 47085 146561 47113
rect 146589 47085 156357 47113
rect 156385 47085 156419 47113
rect 156447 47085 156481 47113
rect 156509 47085 156543 47113
rect 156571 47085 161859 47113
rect 161887 47085 161921 47113
rect 161949 47085 171717 47113
rect 171745 47085 171779 47113
rect 171807 47085 171841 47113
rect 171869 47085 171903 47113
rect 171931 47085 177219 47113
rect 177247 47085 177281 47113
rect 177309 47085 187077 47113
rect 187105 47085 187139 47113
rect 187167 47085 187201 47113
rect 187229 47085 187263 47113
rect 187291 47085 192579 47113
rect 192607 47085 192641 47113
rect 192669 47085 202437 47113
rect 202465 47085 202499 47113
rect 202527 47085 202561 47113
rect 202589 47085 202623 47113
rect 202651 47085 207939 47113
rect 207967 47085 208001 47113
rect 208029 47085 217797 47113
rect 217825 47085 217859 47113
rect 217887 47085 217921 47113
rect 217949 47085 217983 47113
rect 218011 47085 223299 47113
rect 223327 47085 223361 47113
rect 223389 47085 233157 47113
rect 233185 47085 233219 47113
rect 233247 47085 233281 47113
rect 233309 47085 233343 47113
rect 233371 47085 238659 47113
rect 238687 47085 238721 47113
rect 238749 47085 248517 47113
rect 248545 47085 248579 47113
rect 248607 47085 248641 47113
rect 248669 47085 248703 47113
rect 248731 47085 254019 47113
rect 254047 47085 254081 47113
rect 254109 47085 263877 47113
rect 263905 47085 263939 47113
rect 263967 47085 264001 47113
rect 264029 47085 264063 47113
rect 264091 47085 269379 47113
rect 269407 47085 269441 47113
rect 269469 47085 279237 47113
rect 279265 47085 279299 47113
rect 279327 47085 279361 47113
rect 279389 47085 279423 47113
rect 279451 47085 284739 47113
rect 284767 47085 284801 47113
rect 284829 47085 294597 47113
rect 294625 47085 294659 47113
rect 294687 47085 294721 47113
rect 294749 47085 294783 47113
rect 294811 47085 298248 47113
rect 298276 47085 298310 47113
rect 298338 47085 298372 47113
rect 298400 47085 298434 47113
rect 298462 47085 298990 47113
rect -958 47051 298990 47085
rect -958 47023 -430 47051
rect -402 47023 -368 47051
rect -340 47023 -306 47051
rect -278 47023 -244 47051
rect -216 47023 2757 47051
rect 2785 47023 2819 47051
rect 2847 47023 2881 47051
rect 2909 47023 2943 47051
rect 2971 47023 8259 47051
rect 8287 47023 8321 47051
rect 8349 47023 18117 47051
rect 18145 47023 18179 47051
rect 18207 47023 18241 47051
rect 18269 47023 18303 47051
rect 18331 47023 23619 47051
rect 23647 47023 23681 47051
rect 23709 47023 33477 47051
rect 33505 47023 33539 47051
rect 33567 47023 33601 47051
rect 33629 47023 33663 47051
rect 33691 47023 38979 47051
rect 39007 47023 39041 47051
rect 39069 47023 48837 47051
rect 48865 47023 48899 47051
rect 48927 47023 48961 47051
rect 48989 47023 49023 47051
rect 49051 47023 54339 47051
rect 54367 47023 54401 47051
rect 54429 47023 64197 47051
rect 64225 47023 64259 47051
rect 64287 47023 64321 47051
rect 64349 47023 64383 47051
rect 64411 47023 69699 47051
rect 69727 47023 69761 47051
rect 69789 47023 79557 47051
rect 79585 47023 79619 47051
rect 79647 47023 79681 47051
rect 79709 47023 79743 47051
rect 79771 47023 85059 47051
rect 85087 47023 85121 47051
rect 85149 47023 94917 47051
rect 94945 47023 94979 47051
rect 95007 47023 95041 47051
rect 95069 47023 95103 47051
rect 95131 47023 100419 47051
rect 100447 47023 100481 47051
rect 100509 47023 110277 47051
rect 110305 47023 110339 47051
rect 110367 47023 110401 47051
rect 110429 47023 110463 47051
rect 110491 47023 115779 47051
rect 115807 47023 115841 47051
rect 115869 47023 125637 47051
rect 125665 47023 125699 47051
rect 125727 47023 125761 47051
rect 125789 47023 125823 47051
rect 125851 47023 131139 47051
rect 131167 47023 131201 47051
rect 131229 47023 140997 47051
rect 141025 47023 141059 47051
rect 141087 47023 141121 47051
rect 141149 47023 141183 47051
rect 141211 47023 146499 47051
rect 146527 47023 146561 47051
rect 146589 47023 156357 47051
rect 156385 47023 156419 47051
rect 156447 47023 156481 47051
rect 156509 47023 156543 47051
rect 156571 47023 161859 47051
rect 161887 47023 161921 47051
rect 161949 47023 171717 47051
rect 171745 47023 171779 47051
rect 171807 47023 171841 47051
rect 171869 47023 171903 47051
rect 171931 47023 177219 47051
rect 177247 47023 177281 47051
rect 177309 47023 187077 47051
rect 187105 47023 187139 47051
rect 187167 47023 187201 47051
rect 187229 47023 187263 47051
rect 187291 47023 192579 47051
rect 192607 47023 192641 47051
rect 192669 47023 202437 47051
rect 202465 47023 202499 47051
rect 202527 47023 202561 47051
rect 202589 47023 202623 47051
rect 202651 47023 207939 47051
rect 207967 47023 208001 47051
rect 208029 47023 217797 47051
rect 217825 47023 217859 47051
rect 217887 47023 217921 47051
rect 217949 47023 217983 47051
rect 218011 47023 223299 47051
rect 223327 47023 223361 47051
rect 223389 47023 233157 47051
rect 233185 47023 233219 47051
rect 233247 47023 233281 47051
rect 233309 47023 233343 47051
rect 233371 47023 238659 47051
rect 238687 47023 238721 47051
rect 238749 47023 248517 47051
rect 248545 47023 248579 47051
rect 248607 47023 248641 47051
rect 248669 47023 248703 47051
rect 248731 47023 254019 47051
rect 254047 47023 254081 47051
rect 254109 47023 263877 47051
rect 263905 47023 263939 47051
rect 263967 47023 264001 47051
rect 264029 47023 264063 47051
rect 264091 47023 269379 47051
rect 269407 47023 269441 47051
rect 269469 47023 279237 47051
rect 279265 47023 279299 47051
rect 279327 47023 279361 47051
rect 279389 47023 279423 47051
rect 279451 47023 284739 47051
rect 284767 47023 284801 47051
rect 284829 47023 294597 47051
rect 294625 47023 294659 47051
rect 294687 47023 294721 47051
rect 294749 47023 294783 47051
rect 294811 47023 298248 47051
rect 298276 47023 298310 47051
rect 298338 47023 298372 47051
rect 298400 47023 298434 47051
rect 298462 47023 298990 47051
rect -958 46989 298990 47023
rect -958 46961 -430 46989
rect -402 46961 -368 46989
rect -340 46961 -306 46989
rect -278 46961 -244 46989
rect -216 46961 2757 46989
rect 2785 46961 2819 46989
rect 2847 46961 2881 46989
rect 2909 46961 2943 46989
rect 2971 46961 8259 46989
rect 8287 46961 8321 46989
rect 8349 46961 18117 46989
rect 18145 46961 18179 46989
rect 18207 46961 18241 46989
rect 18269 46961 18303 46989
rect 18331 46961 23619 46989
rect 23647 46961 23681 46989
rect 23709 46961 33477 46989
rect 33505 46961 33539 46989
rect 33567 46961 33601 46989
rect 33629 46961 33663 46989
rect 33691 46961 38979 46989
rect 39007 46961 39041 46989
rect 39069 46961 48837 46989
rect 48865 46961 48899 46989
rect 48927 46961 48961 46989
rect 48989 46961 49023 46989
rect 49051 46961 54339 46989
rect 54367 46961 54401 46989
rect 54429 46961 64197 46989
rect 64225 46961 64259 46989
rect 64287 46961 64321 46989
rect 64349 46961 64383 46989
rect 64411 46961 69699 46989
rect 69727 46961 69761 46989
rect 69789 46961 79557 46989
rect 79585 46961 79619 46989
rect 79647 46961 79681 46989
rect 79709 46961 79743 46989
rect 79771 46961 85059 46989
rect 85087 46961 85121 46989
rect 85149 46961 94917 46989
rect 94945 46961 94979 46989
rect 95007 46961 95041 46989
rect 95069 46961 95103 46989
rect 95131 46961 100419 46989
rect 100447 46961 100481 46989
rect 100509 46961 110277 46989
rect 110305 46961 110339 46989
rect 110367 46961 110401 46989
rect 110429 46961 110463 46989
rect 110491 46961 115779 46989
rect 115807 46961 115841 46989
rect 115869 46961 125637 46989
rect 125665 46961 125699 46989
rect 125727 46961 125761 46989
rect 125789 46961 125823 46989
rect 125851 46961 131139 46989
rect 131167 46961 131201 46989
rect 131229 46961 140997 46989
rect 141025 46961 141059 46989
rect 141087 46961 141121 46989
rect 141149 46961 141183 46989
rect 141211 46961 146499 46989
rect 146527 46961 146561 46989
rect 146589 46961 156357 46989
rect 156385 46961 156419 46989
rect 156447 46961 156481 46989
rect 156509 46961 156543 46989
rect 156571 46961 161859 46989
rect 161887 46961 161921 46989
rect 161949 46961 171717 46989
rect 171745 46961 171779 46989
rect 171807 46961 171841 46989
rect 171869 46961 171903 46989
rect 171931 46961 177219 46989
rect 177247 46961 177281 46989
rect 177309 46961 187077 46989
rect 187105 46961 187139 46989
rect 187167 46961 187201 46989
rect 187229 46961 187263 46989
rect 187291 46961 192579 46989
rect 192607 46961 192641 46989
rect 192669 46961 202437 46989
rect 202465 46961 202499 46989
rect 202527 46961 202561 46989
rect 202589 46961 202623 46989
rect 202651 46961 207939 46989
rect 207967 46961 208001 46989
rect 208029 46961 217797 46989
rect 217825 46961 217859 46989
rect 217887 46961 217921 46989
rect 217949 46961 217983 46989
rect 218011 46961 223299 46989
rect 223327 46961 223361 46989
rect 223389 46961 233157 46989
rect 233185 46961 233219 46989
rect 233247 46961 233281 46989
rect 233309 46961 233343 46989
rect 233371 46961 238659 46989
rect 238687 46961 238721 46989
rect 238749 46961 248517 46989
rect 248545 46961 248579 46989
rect 248607 46961 248641 46989
rect 248669 46961 248703 46989
rect 248731 46961 254019 46989
rect 254047 46961 254081 46989
rect 254109 46961 263877 46989
rect 263905 46961 263939 46989
rect 263967 46961 264001 46989
rect 264029 46961 264063 46989
rect 264091 46961 269379 46989
rect 269407 46961 269441 46989
rect 269469 46961 279237 46989
rect 279265 46961 279299 46989
rect 279327 46961 279361 46989
rect 279389 46961 279423 46989
rect 279451 46961 284739 46989
rect 284767 46961 284801 46989
rect 284829 46961 294597 46989
rect 294625 46961 294659 46989
rect 294687 46961 294721 46989
rect 294749 46961 294783 46989
rect 294811 46961 298248 46989
rect 298276 46961 298310 46989
rect 298338 46961 298372 46989
rect 298400 46961 298434 46989
rect 298462 46961 298990 46989
rect -958 46913 298990 46961
rect -958 41175 298990 41223
rect -958 41147 -910 41175
rect -882 41147 -848 41175
rect -820 41147 -786 41175
rect -758 41147 -724 41175
rect -696 41147 4617 41175
rect 4645 41147 4679 41175
rect 4707 41147 4741 41175
rect 4769 41147 4803 41175
rect 4831 41147 15939 41175
rect 15967 41147 16001 41175
rect 16029 41147 19977 41175
rect 20005 41147 20039 41175
rect 20067 41147 20101 41175
rect 20129 41147 20163 41175
rect 20191 41147 31299 41175
rect 31327 41147 31361 41175
rect 31389 41147 35337 41175
rect 35365 41147 35399 41175
rect 35427 41147 35461 41175
rect 35489 41147 35523 41175
rect 35551 41147 46659 41175
rect 46687 41147 46721 41175
rect 46749 41147 50697 41175
rect 50725 41147 50759 41175
rect 50787 41147 50821 41175
rect 50849 41147 50883 41175
rect 50911 41147 62019 41175
rect 62047 41147 62081 41175
rect 62109 41147 66057 41175
rect 66085 41147 66119 41175
rect 66147 41147 66181 41175
rect 66209 41147 66243 41175
rect 66271 41147 77379 41175
rect 77407 41147 77441 41175
rect 77469 41147 81417 41175
rect 81445 41147 81479 41175
rect 81507 41147 81541 41175
rect 81569 41147 81603 41175
rect 81631 41147 92739 41175
rect 92767 41147 92801 41175
rect 92829 41147 96777 41175
rect 96805 41147 96839 41175
rect 96867 41147 96901 41175
rect 96929 41147 96963 41175
rect 96991 41147 108099 41175
rect 108127 41147 108161 41175
rect 108189 41147 112137 41175
rect 112165 41147 112199 41175
rect 112227 41147 112261 41175
rect 112289 41147 112323 41175
rect 112351 41147 123459 41175
rect 123487 41147 123521 41175
rect 123549 41147 127497 41175
rect 127525 41147 127559 41175
rect 127587 41147 127621 41175
rect 127649 41147 127683 41175
rect 127711 41147 138819 41175
rect 138847 41147 138881 41175
rect 138909 41147 142857 41175
rect 142885 41147 142919 41175
rect 142947 41147 142981 41175
rect 143009 41147 143043 41175
rect 143071 41147 154179 41175
rect 154207 41147 154241 41175
rect 154269 41147 158217 41175
rect 158245 41147 158279 41175
rect 158307 41147 158341 41175
rect 158369 41147 158403 41175
rect 158431 41147 169539 41175
rect 169567 41147 169601 41175
rect 169629 41147 173577 41175
rect 173605 41147 173639 41175
rect 173667 41147 173701 41175
rect 173729 41147 173763 41175
rect 173791 41147 184899 41175
rect 184927 41147 184961 41175
rect 184989 41147 188937 41175
rect 188965 41147 188999 41175
rect 189027 41147 189061 41175
rect 189089 41147 189123 41175
rect 189151 41147 200259 41175
rect 200287 41147 200321 41175
rect 200349 41147 204297 41175
rect 204325 41147 204359 41175
rect 204387 41147 204421 41175
rect 204449 41147 204483 41175
rect 204511 41147 215619 41175
rect 215647 41147 215681 41175
rect 215709 41147 219657 41175
rect 219685 41147 219719 41175
rect 219747 41147 219781 41175
rect 219809 41147 219843 41175
rect 219871 41147 230979 41175
rect 231007 41147 231041 41175
rect 231069 41147 235017 41175
rect 235045 41147 235079 41175
rect 235107 41147 235141 41175
rect 235169 41147 235203 41175
rect 235231 41147 246339 41175
rect 246367 41147 246401 41175
rect 246429 41147 250377 41175
rect 250405 41147 250439 41175
rect 250467 41147 250501 41175
rect 250529 41147 250563 41175
rect 250591 41147 261699 41175
rect 261727 41147 261761 41175
rect 261789 41147 265737 41175
rect 265765 41147 265799 41175
rect 265827 41147 265861 41175
rect 265889 41147 265923 41175
rect 265951 41147 277059 41175
rect 277087 41147 277121 41175
rect 277149 41147 281097 41175
rect 281125 41147 281159 41175
rect 281187 41147 281221 41175
rect 281249 41147 281283 41175
rect 281311 41147 296457 41175
rect 296485 41147 296519 41175
rect 296547 41147 296581 41175
rect 296609 41147 296643 41175
rect 296671 41147 298728 41175
rect 298756 41147 298790 41175
rect 298818 41147 298852 41175
rect 298880 41147 298914 41175
rect 298942 41147 298990 41175
rect -958 41113 298990 41147
rect -958 41085 -910 41113
rect -882 41085 -848 41113
rect -820 41085 -786 41113
rect -758 41085 -724 41113
rect -696 41085 4617 41113
rect 4645 41085 4679 41113
rect 4707 41085 4741 41113
rect 4769 41085 4803 41113
rect 4831 41085 15939 41113
rect 15967 41085 16001 41113
rect 16029 41085 19977 41113
rect 20005 41085 20039 41113
rect 20067 41085 20101 41113
rect 20129 41085 20163 41113
rect 20191 41085 31299 41113
rect 31327 41085 31361 41113
rect 31389 41085 35337 41113
rect 35365 41085 35399 41113
rect 35427 41085 35461 41113
rect 35489 41085 35523 41113
rect 35551 41085 46659 41113
rect 46687 41085 46721 41113
rect 46749 41085 50697 41113
rect 50725 41085 50759 41113
rect 50787 41085 50821 41113
rect 50849 41085 50883 41113
rect 50911 41085 62019 41113
rect 62047 41085 62081 41113
rect 62109 41085 66057 41113
rect 66085 41085 66119 41113
rect 66147 41085 66181 41113
rect 66209 41085 66243 41113
rect 66271 41085 77379 41113
rect 77407 41085 77441 41113
rect 77469 41085 81417 41113
rect 81445 41085 81479 41113
rect 81507 41085 81541 41113
rect 81569 41085 81603 41113
rect 81631 41085 92739 41113
rect 92767 41085 92801 41113
rect 92829 41085 96777 41113
rect 96805 41085 96839 41113
rect 96867 41085 96901 41113
rect 96929 41085 96963 41113
rect 96991 41085 108099 41113
rect 108127 41085 108161 41113
rect 108189 41085 112137 41113
rect 112165 41085 112199 41113
rect 112227 41085 112261 41113
rect 112289 41085 112323 41113
rect 112351 41085 123459 41113
rect 123487 41085 123521 41113
rect 123549 41085 127497 41113
rect 127525 41085 127559 41113
rect 127587 41085 127621 41113
rect 127649 41085 127683 41113
rect 127711 41085 138819 41113
rect 138847 41085 138881 41113
rect 138909 41085 142857 41113
rect 142885 41085 142919 41113
rect 142947 41085 142981 41113
rect 143009 41085 143043 41113
rect 143071 41085 154179 41113
rect 154207 41085 154241 41113
rect 154269 41085 158217 41113
rect 158245 41085 158279 41113
rect 158307 41085 158341 41113
rect 158369 41085 158403 41113
rect 158431 41085 169539 41113
rect 169567 41085 169601 41113
rect 169629 41085 173577 41113
rect 173605 41085 173639 41113
rect 173667 41085 173701 41113
rect 173729 41085 173763 41113
rect 173791 41085 184899 41113
rect 184927 41085 184961 41113
rect 184989 41085 188937 41113
rect 188965 41085 188999 41113
rect 189027 41085 189061 41113
rect 189089 41085 189123 41113
rect 189151 41085 200259 41113
rect 200287 41085 200321 41113
rect 200349 41085 204297 41113
rect 204325 41085 204359 41113
rect 204387 41085 204421 41113
rect 204449 41085 204483 41113
rect 204511 41085 215619 41113
rect 215647 41085 215681 41113
rect 215709 41085 219657 41113
rect 219685 41085 219719 41113
rect 219747 41085 219781 41113
rect 219809 41085 219843 41113
rect 219871 41085 230979 41113
rect 231007 41085 231041 41113
rect 231069 41085 235017 41113
rect 235045 41085 235079 41113
rect 235107 41085 235141 41113
rect 235169 41085 235203 41113
rect 235231 41085 246339 41113
rect 246367 41085 246401 41113
rect 246429 41085 250377 41113
rect 250405 41085 250439 41113
rect 250467 41085 250501 41113
rect 250529 41085 250563 41113
rect 250591 41085 261699 41113
rect 261727 41085 261761 41113
rect 261789 41085 265737 41113
rect 265765 41085 265799 41113
rect 265827 41085 265861 41113
rect 265889 41085 265923 41113
rect 265951 41085 277059 41113
rect 277087 41085 277121 41113
rect 277149 41085 281097 41113
rect 281125 41085 281159 41113
rect 281187 41085 281221 41113
rect 281249 41085 281283 41113
rect 281311 41085 296457 41113
rect 296485 41085 296519 41113
rect 296547 41085 296581 41113
rect 296609 41085 296643 41113
rect 296671 41085 298728 41113
rect 298756 41085 298790 41113
rect 298818 41085 298852 41113
rect 298880 41085 298914 41113
rect 298942 41085 298990 41113
rect -958 41051 298990 41085
rect -958 41023 -910 41051
rect -882 41023 -848 41051
rect -820 41023 -786 41051
rect -758 41023 -724 41051
rect -696 41023 4617 41051
rect 4645 41023 4679 41051
rect 4707 41023 4741 41051
rect 4769 41023 4803 41051
rect 4831 41023 15939 41051
rect 15967 41023 16001 41051
rect 16029 41023 19977 41051
rect 20005 41023 20039 41051
rect 20067 41023 20101 41051
rect 20129 41023 20163 41051
rect 20191 41023 31299 41051
rect 31327 41023 31361 41051
rect 31389 41023 35337 41051
rect 35365 41023 35399 41051
rect 35427 41023 35461 41051
rect 35489 41023 35523 41051
rect 35551 41023 46659 41051
rect 46687 41023 46721 41051
rect 46749 41023 50697 41051
rect 50725 41023 50759 41051
rect 50787 41023 50821 41051
rect 50849 41023 50883 41051
rect 50911 41023 62019 41051
rect 62047 41023 62081 41051
rect 62109 41023 66057 41051
rect 66085 41023 66119 41051
rect 66147 41023 66181 41051
rect 66209 41023 66243 41051
rect 66271 41023 77379 41051
rect 77407 41023 77441 41051
rect 77469 41023 81417 41051
rect 81445 41023 81479 41051
rect 81507 41023 81541 41051
rect 81569 41023 81603 41051
rect 81631 41023 92739 41051
rect 92767 41023 92801 41051
rect 92829 41023 96777 41051
rect 96805 41023 96839 41051
rect 96867 41023 96901 41051
rect 96929 41023 96963 41051
rect 96991 41023 108099 41051
rect 108127 41023 108161 41051
rect 108189 41023 112137 41051
rect 112165 41023 112199 41051
rect 112227 41023 112261 41051
rect 112289 41023 112323 41051
rect 112351 41023 123459 41051
rect 123487 41023 123521 41051
rect 123549 41023 127497 41051
rect 127525 41023 127559 41051
rect 127587 41023 127621 41051
rect 127649 41023 127683 41051
rect 127711 41023 138819 41051
rect 138847 41023 138881 41051
rect 138909 41023 142857 41051
rect 142885 41023 142919 41051
rect 142947 41023 142981 41051
rect 143009 41023 143043 41051
rect 143071 41023 154179 41051
rect 154207 41023 154241 41051
rect 154269 41023 158217 41051
rect 158245 41023 158279 41051
rect 158307 41023 158341 41051
rect 158369 41023 158403 41051
rect 158431 41023 169539 41051
rect 169567 41023 169601 41051
rect 169629 41023 173577 41051
rect 173605 41023 173639 41051
rect 173667 41023 173701 41051
rect 173729 41023 173763 41051
rect 173791 41023 184899 41051
rect 184927 41023 184961 41051
rect 184989 41023 188937 41051
rect 188965 41023 188999 41051
rect 189027 41023 189061 41051
rect 189089 41023 189123 41051
rect 189151 41023 200259 41051
rect 200287 41023 200321 41051
rect 200349 41023 204297 41051
rect 204325 41023 204359 41051
rect 204387 41023 204421 41051
rect 204449 41023 204483 41051
rect 204511 41023 215619 41051
rect 215647 41023 215681 41051
rect 215709 41023 219657 41051
rect 219685 41023 219719 41051
rect 219747 41023 219781 41051
rect 219809 41023 219843 41051
rect 219871 41023 230979 41051
rect 231007 41023 231041 41051
rect 231069 41023 235017 41051
rect 235045 41023 235079 41051
rect 235107 41023 235141 41051
rect 235169 41023 235203 41051
rect 235231 41023 246339 41051
rect 246367 41023 246401 41051
rect 246429 41023 250377 41051
rect 250405 41023 250439 41051
rect 250467 41023 250501 41051
rect 250529 41023 250563 41051
rect 250591 41023 261699 41051
rect 261727 41023 261761 41051
rect 261789 41023 265737 41051
rect 265765 41023 265799 41051
rect 265827 41023 265861 41051
rect 265889 41023 265923 41051
rect 265951 41023 277059 41051
rect 277087 41023 277121 41051
rect 277149 41023 281097 41051
rect 281125 41023 281159 41051
rect 281187 41023 281221 41051
rect 281249 41023 281283 41051
rect 281311 41023 296457 41051
rect 296485 41023 296519 41051
rect 296547 41023 296581 41051
rect 296609 41023 296643 41051
rect 296671 41023 298728 41051
rect 298756 41023 298790 41051
rect 298818 41023 298852 41051
rect 298880 41023 298914 41051
rect 298942 41023 298990 41051
rect -958 40989 298990 41023
rect -958 40961 -910 40989
rect -882 40961 -848 40989
rect -820 40961 -786 40989
rect -758 40961 -724 40989
rect -696 40961 4617 40989
rect 4645 40961 4679 40989
rect 4707 40961 4741 40989
rect 4769 40961 4803 40989
rect 4831 40961 15939 40989
rect 15967 40961 16001 40989
rect 16029 40961 19977 40989
rect 20005 40961 20039 40989
rect 20067 40961 20101 40989
rect 20129 40961 20163 40989
rect 20191 40961 31299 40989
rect 31327 40961 31361 40989
rect 31389 40961 35337 40989
rect 35365 40961 35399 40989
rect 35427 40961 35461 40989
rect 35489 40961 35523 40989
rect 35551 40961 46659 40989
rect 46687 40961 46721 40989
rect 46749 40961 50697 40989
rect 50725 40961 50759 40989
rect 50787 40961 50821 40989
rect 50849 40961 50883 40989
rect 50911 40961 62019 40989
rect 62047 40961 62081 40989
rect 62109 40961 66057 40989
rect 66085 40961 66119 40989
rect 66147 40961 66181 40989
rect 66209 40961 66243 40989
rect 66271 40961 77379 40989
rect 77407 40961 77441 40989
rect 77469 40961 81417 40989
rect 81445 40961 81479 40989
rect 81507 40961 81541 40989
rect 81569 40961 81603 40989
rect 81631 40961 92739 40989
rect 92767 40961 92801 40989
rect 92829 40961 96777 40989
rect 96805 40961 96839 40989
rect 96867 40961 96901 40989
rect 96929 40961 96963 40989
rect 96991 40961 108099 40989
rect 108127 40961 108161 40989
rect 108189 40961 112137 40989
rect 112165 40961 112199 40989
rect 112227 40961 112261 40989
rect 112289 40961 112323 40989
rect 112351 40961 123459 40989
rect 123487 40961 123521 40989
rect 123549 40961 127497 40989
rect 127525 40961 127559 40989
rect 127587 40961 127621 40989
rect 127649 40961 127683 40989
rect 127711 40961 138819 40989
rect 138847 40961 138881 40989
rect 138909 40961 142857 40989
rect 142885 40961 142919 40989
rect 142947 40961 142981 40989
rect 143009 40961 143043 40989
rect 143071 40961 154179 40989
rect 154207 40961 154241 40989
rect 154269 40961 158217 40989
rect 158245 40961 158279 40989
rect 158307 40961 158341 40989
rect 158369 40961 158403 40989
rect 158431 40961 169539 40989
rect 169567 40961 169601 40989
rect 169629 40961 173577 40989
rect 173605 40961 173639 40989
rect 173667 40961 173701 40989
rect 173729 40961 173763 40989
rect 173791 40961 184899 40989
rect 184927 40961 184961 40989
rect 184989 40961 188937 40989
rect 188965 40961 188999 40989
rect 189027 40961 189061 40989
rect 189089 40961 189123 40989
rect 189151 40961 200259 40989
rect 200287 40961 200321 40989
rect 200349 40961 204297 40989
rect 204325 40961 204359 40989
rect 204387 40961 204421 40989
rect 204449 40961 204483 40989
rect 204511 40961 215619 40989
rect 215647 40961 215681 40989
rect 215709 40961 219657 40989
rect 219685 40961 219719 40989
rect 219747 40961 219781 40989
rect 219809 40961 219843 40989
rect 219871 40961 230979 40989
rect 231007 40961 231041 40989
rect 231069 40961 235017 40989
rect 235045 40961 235079 40989
rect 235107 40961 235141 40989
rect 235169 40961 235203 40989
rect 235231 40961 246339 40989
rect 246367 40961 246401 40989
rect 246429 40961 250377 40989
rect 250405 40961 250439 40989
rect 250467 40961 250501 40989
rect 250529 40961 250563 40989
rect 250591 40961 261699 40989
rect 261727 40961 261761 40989
rect 261789 40961 265737 40989
rect 265765 40961 265799 40989
rect 265827 40961 265861 40989
rect 265889 40961 265923 40989
rect 265951 40961 277059 40989
rect 277087 40961 277121 40989
rect 277149 40961 281097 40989
rect 281125 40961 281159 40989
rect 281187 40961 281221 40989
rect 281249 40961 281283 40989
rect 281311 40961 296457 40989
rect 296485 40961 296519 40989
rect 296547 40961 296581 40989
rect 296609 40961 296643 40989
rect 296671 40961 298728 40989
rect 298756 40961 298790 40989
rect 298818 40961 298852 40989
rect 298880 40961 298914 40989
rect 298942 40961 298990 40989
rect -958 40913 298990 40961
rect -958 38175 298990 38223
rect -958 38147 -430 38175
rect -402 38147 -368 38175
rect -340 38147 -306 38175
rect -278 38147 -244 38175
rect -216 38147 2757 38175
rect 2785 38147 2819 38175
rect 2847 38147 2881 38175
rect 2909 38147 2943 38175
rect 2971 38147 8259 38175
rect 8287 38147 8321 38175
rect 8349 38147 18117 38175
rect 18145 38147 18179 38175
rect 18207 38147 18241 38175
rect 18269 38147 18303 38175
rect 18331 38147 23619 38175
rect 23647 38147 23681 38175
rect 23709 38147 33477 38175
rect 33505 38147 33539 38175
rect 33567 38147 33601 38175
rect 33629 38147 33663 38175
rect 33691 38147 38979 38175
rect 39007 38147 39041 38175
rect 39069 38147 48837 38175
rect 48865 38147 48899 38175
rect 48927 38147 48961 38175
rect 48989 38147 49023 38175
rect 49051 38147 54339 38175
rect 54367 38147 54401 38175
rect 54429 38147 64197 38175
rect 64225 38147 64259 38175
rect 64287 38147 64321 38175
rect 64349 38147 64383 38175
rect 64411 38147 69699 38175
rect 69727 38147 69761 38175
rect 69789 38147 79557 38175
rect 79585 38147 79619 38175
rect 79647 38147 79681 38175
rect 79709 38147 79743 38175
rect 79771 38147 85059 38175
rect 85087 38147 85121 38175
rect 85149 38147 94917 38175
rect 94945 38147 94979 38175
rect 95007 38147 95041 38175
rect 95069 38147 95103 38175
rect 95131 38147 100419 38175
rect 100447 38147 100481 38175
rect 100509 38147 110277 38175
rect 110305 38147 110339 38175
rect 110367 38147 110401 38175
rect 110429 38147 110463 38175
rect 110491 38147 115779 38175
rect 115807 38147 115841 38175
rect 115869 38147 125637 38175
rect 125665 38147 125699 38175
rect 125727 38147 125761 38175
rect 125789 38147 125823 38175
rect 125851 38147 131139 38175
rect 131167 38147 131201 38175
rect 131229 38147 140997 38175
rect 141025 38147 141059 38175
rect 141087 38147 141121 38175
rect 141149 38147 141183 38175
rect 141211 38147 146499 38175
rect 146527 38147 146561 38175
rect 146589 38147 156357 38175
rect 156385 38147 156419 38175
rect 156447 38147 156481 38175
rect 156509 38147 156543 38175
rect 156571 38147 161859 38175
rect 161887 38147 161921 38175
rect 161949 38147 171717 38175
rect 171745 38147 171779 38175
rect 171807 38147 171841 38175
rect 171869 38147 171903 38175
rect 171931 38147 177219 38175
rect 177247 38147 177281 38175
rect 177309 38147 187077 38175
rect 187105 38147 187139 38175
rect 187167 38147 187201 38175
rect 187229 38147 187263 38175
rect 187291 38147 192579 38175
rect 192607 38147 192641 38175
rect 192669 38147 202437 38175
rect 202465 38147 202499 38175
rect 202527 38147 202561 38175
rect 202589 38147 202623 38175
rect 202651 38147 207939 38175
rect 207967 38147 208001 38175
rect 208029 38147 217797 38175
rect 217825 38147 217859 38175
rect 217887 38147 217921 38175
rect 217949 38147 217983 38175
rect 218011 38147 223299 38175
rect 223327 38147 223361 38175
rect 223389 38147 233157 38175
rect 233185 38147 233219 38175
rect 233247 38147 233281 38175
rect 233309 38147 233343 38175
rect 233371 38147 238659 38175
rect 238687 38147 238721 38175
rect 238749 38147 248517 38175
rect 248545 38147 248579 38175
rect 248607 38147 248641 38175
rect 248669 38147 248703 38175
rect 248731 38147 254019 38175
rect 254047 38147 254081 38175
rect 254109 38147 263877 38175
rect 263905 38147 263939 38175
rect 263967 38147 264001 38175
rect 264029 38147 264063 38175
rect 264091 38147 269379 38175
rect 269407 38147 269441 38175
rect 269469 38147 279237 38175
rect 279265 38147 279299 38175
rect 279327 38147 279361 38175
rect 279389 38147 279423 38175
rect 279451 38147 284739 38175
rect 284767 38147 284801 38175
rect 284829 38147 294597 38175
rect 294625 38147 294659 38175
rect 294687 38147 294721 38175
rect 294749 38147 294783 38175
rect 294811 38147 298248 38175
rect 298276 38147 298310 38175
rect 298338 38147 298372 38175
rect 298400 38147 298434 38175
rect 298462 38147 298990 38175
rect -958 38113 298990 38147
rect -958 38085 -430 38113
rect -402 38085 -368 38113
rect -340 38085 -306 38113
rect -278 38085 -244 38113
rect -216 38085 2757 38113
rect 2785 38085 2819 38113
rect 2847 38085 2881 38113
rect 2909 38085 2943 38113
rect 2971 38085 8259 38113
rect 8287 38085 8321 38113
rect 8349 38085 18117 38113
rect 18145 38085 18179 38113
rect 18207 38085 18241 38113
rect 18269 38085 18303 38113
rect 18331 38085 23619 38113
rect 23647 38085 23681 38113
rect 23709 38085 33477 38113
rect 33505 38085 33539 38113
rect 33567 38085 33601 38113
rect 33629 38085 33663 38113
rect 33691 38085 38979 38113
rect 39007 38085 39041 38113
rect 39069 38085 48837 38113
rect 48865 38085 48899 38113
rect 48927 38085 48961 38113
rect 48989 38085 49023 38113
rect 49051 38085 54339 38113
rect 54367 38085 54401 38113
rect 54429 38085 64197 38113
rect 64225 38085 64259 38113
rect 64287 38085 64321 38113
rect 64349 38085 64383 38113
rect 64411 38085 69699 38113
rect 69727 38085 69761 38113
rect 69789 38085 79557 38113
rect 79585 38085 79619 38113
rect 79647 38085 79681 38113
rect 79709 38085 79743 38113
rect 79771 38085 85059 38113
rect 85087 38085 85121 38113
rect 85149 38085 94917 38113
rect 94945 38085 94979 38113
rect 95007 38085 95041 38113
rect 95069 38085 95103 38113
rect 95131 38085 100419 38113
rect 100447 38085 100481 38113
rect 100509 38085 110277 38113
rect 110305 38085 110339 38113
rect 110367 38085 110401 38113
rect 110429 38085 110463 38113
rect 110491 38085 115779 38113
rect 115807 38085 115841 38113
rect 115869 38085 125637 38113
rect 125665 38085 125699 38113
rect 125727 38085 125761 38113
rect 125789 38085 125823 38113
rect 125851 38085 131139 38113
rect 131167 38085 131201 38113
rect 131229 38085 140997 38113
rect 141025 38085 141059 38113
rect 141087 38085 141121 38113
rect 141149 38085 141183 38113
rect 141211 38085 146499 38113
rect 146527 38085 146561 38113
rect 146589 38085 156357 38113
rect 156385 38085 156419 38113
rect 156447 38085 156481 38113
rect 156509 38085 156543 38113
rect 156571 38085 161859 38113
rect 161887 38085 161921 38113
rect 161949 38085 171717 38113
rect 171745 38085 171779 38113
rect 171807 38085 171841 38113
rect 171869 38085 171903 38113
rect 171931 38085 177219 38113
rect 177247 38085 177281 38113
rect 177309 38085 187077 38113
rect 187105 38085 187139 38113
rect 187167 38085 187201 38113
rect 187229 38085 187263 38113
rect 187291 38085 192579 38113
rect 192607 38085 192641 38113
rect 192669 38085 202437 38113
rect 202465 38085 202499 38113
rect 202527 38085 202561 38113
rect 202589 38085 202623 38113
rect 202651 38085 207939 38113
rect 207967 38085 208001 38113
rect 208029 38085 217797 38113
rect 217825 38085 217859 38113
rect 217887 38085 217921 38113
rect 217949 38085 217983 38113
rect 218011 38085 223299 38113
rect 223327 38085 223361 38113
rect 223389 38085 233157 38113
rect 233185 38085 233219 38113
rect 233247 38085 233281 38113
rect 233309 38085 233343 38113
rect 233371 38085 238659 38113
rect 238687 38085 238721 38113
rect 238749 38085 248517 38113
rect 248545 38085 248579 38113
rect 248607 38085 248641 38113
rect 248669 38085 248703 38113
rect 248731 38085 254019 38113
rect 254047 38085 254081 38113
rect 254109 38085 263877 38113
rect 263905 38085 263939 38113
rect 263967 38085 264001 38113
rect 264029 38085 264063 38113
rect 264091 38085 269379 38113
rect 269407 38085 269441 38113
rect 269469 38085 279237 38113
rect 279265 38085 279299 38113
rect 279327 38085 279361 38113
rect 279389 38085 279423 38113
rect 279451 38085 284739 38113
rect 284767 38085 284801 38113
rect 284829 38085 294597 38113
rect 294625 38085 294659 38113
rect 294687 38085 294721 38113
rect 294749 38085 294783 38113
rect 294811 38085 298248 38113
rect 298276 38085 298310 38113
rect 298338 38085 298372 38113
rect 298400 38085 298434 38113
rect 298462 38085 298990 38113
rect -958 38051 298990 38085
rect -958 38023 -430 38051
rect -402 38023 -368 38051
rect -340 38023 -306 38051
rect -278 38023 -244 38051
rect -216 38023 2757 38051
rect 2785 38023 2819 38051
rect 2847 38023 2881 38051
rect 2909 38023 2943 38051
rect 2971 38023 8259 38051
rect 8287 38023 8321 38051
rect 8349 38023 18117 38051
rect 18145 38023 18179 38051
rect 18207 38023 18241 38051
rect 18269 38023 18303 38051
rect 18331 38023 23619 38051
rect 23647 38023 23681 38051
rect 23709 38023 33477 38051
rect 33505 38023 33539 38051
rect 33567 38023 33601 38051
rect 33629 38023 33663 38051
rect 33691 38023 38979 38051
rect 39007 38023 39041 38051
rect 39069 38023 48837 38051
rect 48865 38023 48899 38051
rect 48927 38023 48961 38051
rect 48989 38023 49023 38051
rect 49051 38023 54339 38051
rect 54367 38023 54401 38051
rect 54429 38023 64197 38051
rect 64225 38023 64259 38051
rect 64287 38023 64321 38051
rect 64349 38023 64383 38051
rect 64411 38023 69699 38051
rect 69727 38023 69761 38051
rect 69789 38023 79557 38051
rect 79585 38023 79619 38051
rect 79647 38023 79681 38051
rect 79709 38023 79743 38051
rect 79771 38023 85059 38051
rect 85087 38023 85121 38051
rect 85149 38023 94917 38051
rect 94945 38023 94979 38051
rect 95007 38023 95041 38051
rect 95069 38023 95103 38051
rect 95131 38023 100419 38051
rect 100447 38023 100481 38051
rect 100509 38023 110277 38051
rect 110305 38023 110339 38051
rect 110367 38023 110401 38051
rect 110429 38023 110463 38051
rect 110491 38023 115779 38051
rect 115807 38023 115841 38051
rect 115869 38023 125637 38051
rect 125665 38023 125699 38051
rect 125727 38023 125761 38051
rect 125789 38023 125823 38051
rect 125851 38023 131139 38051
rect 131167 38023 131201 38051
rect 131229 38023 140997 38051
rect 141025 38023 141059 38051
rect 141087 38023 141121 38051
rect 141149 38023 141183 38051
rect 141211 38023 146499 38051
rect 146527 38023 146561 38051
rect 146589 38023 156357 38051
rect 156385 38023 156419 38051
rect 156447 38023 156481 38051
rect 156509 38023 156543 38051
rect 156571 38023 161859 38051
rect 161887 38023 161921 38051
rect 161949 38023 171717 38051
rect 171745 38023 171779 38051
rect 171807 38023 171841 38051
rect 171869 38023 171903 38051
rect 171931 38023 177219 38051
rect 177247 38023 177281 38051
rect 177309 38023 187077 38051
rect 187105 38023 187139 38051
rect 187167 38023 187201 38051
rect 187229 38023 187263 38051
rect 187291 38023 192579 38051
rect 192607 38023 192641 38051
rect 192669 38023 202437 38051
rect 202465 38023 202499 38051
rect 202527 38023 202561 38051
rect 202589 38023 202623 38051
rect 202651 38023 207939 38051
rect 207967 38023 208001 38051
rect 208029 38023 217797 38051
rect 217825 38023 217859 38051
rect 217887 38023 217921 38051
rect 217949 38023 217983 38051
rect 218011 38023 223299 38051
rect 223327 38023 223361 38051
rect 223389 38023 233157 38051
rect 233185 38023 233219 38051
rect 233247 38023 233281 38051
rect 233309 38023 233343 38051
rect 233371 38023 238659 38051
rect 238687 38023 238721 38051
rect 238749 38023 248517 38051
rect 248545 38023 248579 38051
rect 248607 38023 248641 38051
rect 248669 38023 248703 38051
rect 248731 38023 254019 38051
rect 254047 38023 254081 38051
rect 254109 38023 263877 38051
rect 263905 38023 263939 38051
rect 263967 38023 264001 38051
rect 264029 38023 264063 38051
rect 264091 38023 269379 38051
rect 269407 38023 269441 38051
rect 269469 38023 279237 38051
rect 279265 38023 279299 38051
rect 279327 38023 279361 38051
rect 279389 38023 279423 38051
rect 279451 38023 284739 38051
rect 284767 38023 284801 38051
rect 284829 38023 294597 38051
rect 294625 38023 294659 38051
rect 294687 38023 294721 38051
rect 294749 38023 294783 38051
rect 294811 38023 298248 38051
rect 298276 38023 298310 38051
rect 298338 38023 298372 38051
rect 298400 38023 298434 38051
rect 298462 38023 298990 38051
rect -958 37989 298990 38023
rect -958 37961 -430 37989
rect -402 37961 -368 37989
rect -340 37961 -306 37989
rect -278 37961 -244 37989
rect -216 37961 2757 37989
rect 2785 37961 2819 37989
rect 2847 37961 2881 37989
rect 2909 37961 2943 37989
rect 2971 37961 8259 37989
rect 8287 37961 8321 37989
rect 8349 37961 18117 37989
rect 18145 37961 18179 37989
rect 18207 37961 18241 37989
rect 18269 37961 18303 37989
rect 18331 37961 23619 37989
rect 23647 37961 23681 37989
rect 23709 37961 33477 37989
rect 33505 37961 33539 37989
rect 33567 37961 33601 37989
rect 33629 37961 33663 37989
rect 33691 37961 38979 37989
rect 39007 37961 39041 37989
rect 39069 37961 48837 37989
rect 48865 37961 48899 37989
rect 48927 37961 48961 37989
rect 48989 37961 49023 37989
rect 49051 37961 54339 37989
rect 54367 37961 54401 37989
rect 54429 37961 64197 37989
rect 64225 37961 64259 37989
rect 64287 37961 64321 37989
rect 64349 37961 64383 37989
rect 64411 37961 69699 37989
rect 69727 37961 69761 37989
rect 69789 37961 79557 37989
rect 79585 37961 79619 37989
rect 79647 37961 79681 37989
rect 79709 37961 79743 37989
rect 79771 37961 85059 37989
rect 85087 37961 85121 37989
rect 85149 37961 94917 37989
rect 94945 37961 94979 37989
rect 95007 37961 95041 37989
rect 95069 37961 95103 37989
rect 95131 37961 100419 37989
rect 100447 37961 100481 37989
rect 100509 37961 110277 37989
rect 110305 37961 110339 37989
rect 110367 37961 110401 37989
rect 110429 37961 110463 37989
rect 110491 37961 115779 37989
rect 115807 37961 115841 37989
rect 115869 37961 125637 37989
rect 125665 37961 125699 37989
rect 125727 37961 125761 37989
rect 125789 37961 125823 37989
rect 125851 37961 131139 37989
rect 131167 37961 131201 37989
rect 131229 37961 140997 37989
rect 141025 37961 141059 37989
rect 141087 37961 141121 37989
rect 141149 37961 141183 37989
rect 141211 37961 146499 37989
rect 146527 37961 146561 37989
rect 146589 37961 156357 37989
rect 156385 37961 156419 37989
rect 156447 37961 156481 37989
rect 156509 37961 156543 37989
rect 156571 37961 161859 37989
rect 161887 37961 161921 37989
rect 161949 37961 171717 37989
rect 171745 37961 171779 37989
rect 171807 37961 171841 37989
rect 171869 37961 171903 37989
rect 171931 37961 177219 37989
rect 177247 37961 177281 37989
rect 177309 37961 187077 37989
rect 187105 37961 187139 37989
rect 187167 37961 187201 37989
rect 187229 37961 187263 37989
rect 187291 37961 192579 37989
rect 192607 37961 192641 37989
rect 192669 37961 202437 37989
rect 202465 37961 202499 37989
rect 202527 37961 202561 37989
rect 202589 37961 202623 37989
rect 202651 37961 207939 37989
rect 207967 37961 208001 37989
rect 208029 37961 217797 37989
rect 217825 37961 217859 37989
rect 217887 37961 217921 37989
rect 217949 37961 217983 37989
rect 218011 37961 223299 37989
rect 223327 37961 223361 37989
rect 223389 37961 233157 37989
rect 233185 37961 233219 37989
rect 233247 37961 233281 37989
rect 233309 37961 233343 37989
rect 233371 37961 238659 37989
rect 238687 37961 238721 37989
rect 238749 37961 248517 37989
rect 248545 37961 248579 37989
rect 248607 37961 248641 37989
rect 248669 37961 248703 37989
rect 248731 37961 254019 37989
rect 254047 37961 254081 37989
rect 254109 37961 263877 37989
rect 263905 37961 263939 37989
rect 263967 37961 264001 37989
rect 264029 37961 264063 37989
rect 264091 37961 269379 37989
rect 269407 37961 269441 37989
rect 269469 37961 279237 37989
rect 279265 37961 279299 37989
rect 279327 37961 279361 37989
rect 279389 37961 279423 37989
rect 279451 37961 284739 37989
rect 284767 37961 284801 37989
rect 284829 37961 294597 37989
rect 294625 37961 294659 37989
rect 294687 37961 294721 37989
rect 294749 37961 294783 37989
rect 294811 37961 298248 37989
rect 298276 37961 298310 37989
rect 298338 37961 298372 37989
rect 298400 37961 298434 37989
rect 298462 37961 298990 37989
rect -958 37913 298990 37961
rect -958 32175 298990 32223
rect -958 32147 -910 32175
rect -882 32147 -848 32175
rect -820 32147 -786 32175
rect -758 32147 -724 32175
rect -696 32147 4617 32175
rect 4645 32147 4679 32175
rect 4707 32147 4741 32175
rect 4769 32147 4803 32175
rect 4831 32147 15939 32175
rect 15967 32147 16001 32175
rect 16029 32147 19977 32175
rect 20005 32147 20039 32175
rect 20067 32147 20101 32175
rect 20129 32147 20163 32175
rect 20191 32147 31299 32175
rect 31327 32147 31361 32175
rect 31389 32147 35337 32175
rect 35365 32147 35399 32175
rect 35427 32147 35461 32175
rect 35489 32147 35523 32175
rect 35551 32147 46659 32175
rect 46687 32147 46721 32175
rect 46749 32147 50697 32175
rect 50725 32147 50759 32175
rect 50787 32147 50821 32175
rect 50849 32147 50883 32175
rect 50911 32147 62019 32175
rect 62047 32147 62081 32175
rect 62109 32147 66057 32175
rect 66085 32147 66119 32175
rect 66147 32147 66181 32175
rect 66209 32147 66243 32175
rect 66271 32147 77379 32175
rect 77407 32147 77441 32175
rect 77469 32147 81417 32175
rect 81445 32147 81479 32175
rect 81507 32147 81541 32175
rect 81569 32147 81603 32175
rect 81631 32147 92739 32175
rect 92767 32147 92801 32175
rect 92829 32147 96777 32175
rect 96805 32147 96839 32175
rect 96867 32147 96901 32175
rect 96929 32147 96963 32175
rect 96991 32147 108099 32175
rect 108127 32147 108161 32175
rect 108189 32147 112137 32175
rect 112165 32147 112199 32175
rect 112227 32147 112261 32175
rect 112289 32147 112323 32175
rect 112351 32147 123459 32175
rect 123487 32147 123521 32175
rect 123549 32147 127497 32175
rect 127525 32147 127559 32175
rect 127587 32147 127621 32175
rect 127649 32147 127683 32175
rect 127711 32147 138819 32175
rect 138847 32147 138881 32175
rect 138909 32147 142857 32175
rect 142885 32147 142919 32175
rect 142947 32147 142981 32175
rect 143009 32147 143043 32175
rect 143071 32147 154179 32175
rect 154207 32147 154241 32175
rect 154269 32147 158217 32175
rect 158245 32147 158279 32175
rect 158307 32147 158341 32175
rect 158369 32147 158403 32175
rect 158431 32147 169539 32175
rect 169567 32147 169601 32175
rect 169629 32147 173577 32175
rect 173605 32147 173639 32175
rect 173667 32147 173701 32175
rect 173729 32147 173763 32175
rect 173791 32147 184899 32175
rect 184927 32147 184961 32175
rect 184989 32147 188937 32175
rect 188965 32147 188999 32175
rect 189027 32147 189061 32175
rect 189089 32147 189123 32175
rect 189151 32147 200259 32175
rect 200287 32147 200321 32175
rect 200349 32147 204297 32175
rect 204325 32147 204359 32175
rect 204387 32147 204421 32175
rect 204449 32147 204483 32175
rect 204511 32147 215619 32175
rect 215647 32147 215681 32175
rect 215709 32147 219657 32175
rect 219685 32147 219719 32175
rect 219747 32147 219781 32175
rect 219809 32147 219843 32175
rect 219871 32147 230979 32175
rect 231007 32147 231041 32175
rect 231069 32147 235017 32175
rect 235045 32147 235079 32175
rect 235107 32147 235141 32175
rect 235169 32147 235203 32175
rect 235231 32147 246339 32175
rect 246367 32147 246401 32175
rect 246429 32147 250377 32175
rect 250405 32147 250439 32175
rect 250467 32147 250501 32175
rect 250529 32147 250563 32175
rect 250591 32147 261699 32175
rect 261727 32147 261761 32175
rect 261789 32147 265737 32175
rect 265765 32147 265799 32175
rect 265827 32147 265861 32175
rect 265889 32147 265923 32175
rect 265951 32147 277059 32175
rect 277087 32147 277121 32175
rect 277149 32147 281097 32175
rect 281125 32147 281159 32175
rect 281187 32147 281221 32175
rect 281249 32147 281283 32175
rect 281311 32147 296457 32175
rect 296485 32147 296519 32175
rect 296547 32147 296581 32175
rect 296609 32147 296643 32175
rect 296671 32147 298728 32175
rect 298756 32147 298790 32175
rect 298818 32147 298852 32175
rect 298880 32147 298914 32175
rect 298942 32147 298990 32175
rect -958 32113 298990 32147
rect -958 32085 -910 32113
rect -882 32085 -848 32113
rect -820 32085 -786 32113
rect -758 32085 -724 32113
rect -696 32085 4617 32113
rect 4645 32085 4679 32113
rect 4707 32085 4741 32113
rect 4769 32085 4803 32113
rect 4831 32085 15939 32113
rect 15967 32085 16001 32113
rect 16029 32085 19977 32113
rect 20005 32085 20039 32113
rect 20067 32085 20101 32113
rect 20129 32085 20163 32113
rect 20191 32085 31299 32113
rect 31327 32085 31361 32113
rect 31389 32085 35337 32113
rect 35365 32085 35399 32113
rect 35427 32085 35461 32113
rect 35489 32085 35523 32113
rect 35551 32085 46659 32113
rect 46687 32085 46721 32113
rect 46749 32085 50697 32113
rect 50725 32085 50759 32113
rect 50787 32085 50821 32113
rect 50849 32085 50883 32113
rect 50911 32085 62019 32113
rect 62047 32085 62081 32113
rect 62109 32085 66057 32113
rect 66085 32085 66119 32113
rect 66147 32085 66181 32113
rect 66209 32085 66243 32113
rect 66271 32085 77379 32113
rect 77407 32085 77441 32113
rect 77469 32085 81417 32113
rect 81445 32085 81479 32113
rect 81507 32085 81541 32113
rect 81569 32085 81603 32113
rect 81631 32085 92739 32113
rect 92767 32085 92801 32113
rect 92829 32085 96777 32113
rect 96805 32085 96839 32113
rect 96867 32085 96901 32113
rect 96929 32085 96963 32113
rect 96991 32085 108099 32113
rect 108127 32085 108161 32113
rect 108189 32085 112137 32113
rect 112165 32085 112199 32113
rect 112227 32085 112261 32113
rect 112289 32085 112323 32113
rect 112351 32085 123459 32113
rect 123487 32085 123521 32113
rect 123549 32085 127497 32113
rect 127525 32085 127559 32113
rect 127587 32085 127621 32113
rect 127649 32085 127683 32113
rect 127711 32085 138819 32113
rect 138847 32085 138881 32113
rect 138909 32085 142857 32113
rect 142885 32085 142919 32113
rect 142947 32085 142981 32113
rect 143009 32085 143043 32113
rect 143071 32085 154179 32113
rect 154207 32085 154241 32113
rect 154269 32085 158217 32113
rect 158245 32085 158279 32113
rect 158307 32085 158341 32113
rect 158369 32085 158403 32113
rect 158431 32085 169539 32113
rect 169567 32085 169601 32113
rect 169629 32085 173577 32113
rect 173605 32085 173639 32113
rect 173667 32085 173701 32113
rect 173729 32085 173763 32113
rect 173791 32085 184899 32113
rect 184927 32085 184961 32113
rect 184989 32085 188937 32113
rect 188965 32085 188999 32113
rect 189027 32085 189061 32113
rect 189089 32085 189123 32113
rect 189151 32085 200259 32113
rect 200287 32085 200321 32113
rect 200349 32085 204297 32113
rect 204325 32085 204359 32113
rect 204387 32085 204421 32113
rect 204449 32085 204483 32113
rect 204511 32085 215619 32113
rect 215647 32085 215681 32113
rect 215709 32085 219657 32113
rect 219685 32085 219719 32113
rect 219747 32085 219781 32113
rect 219809 32085 219843 32113
rect 219871 32085 230979 32113
rect 231007 32085 231041 32113
rect 231069 32085 235017 32113
rect 235045 32085 235079 32113
rect 235107 32085 235141 32113
rect 235169 32085 235203 32113
rect 235231 32085 246339 32113
rect 246367 32085 246401 32113
rect 246429 32085 250377 32113
rect 250405 32085 250439 32113
rect 250467 32085 250501 32113
rect 250529 32085 250563 32113
rect 250591 32085 261699 32113
rect 261727 32085 261761 32113
rect 261789 32085 265737 32113
rect 265765 32085 265799 32113
rect 265827 32085 265861 32113
rect 265889 32085 265923 32113
rect 265951 32085 277059 32113
rect 277087 32085 277121 32113
rect 277149 32085 281097 32113
rect 281125 32085 281159 32113
rect 281187 32085 281221 32113
rect 281249 32085 281283 32113
rect 281311 32085 296457 32113
rect 296485 32085 296519 32113
rect 296547 32085 296581 32113
rect 296609 32085 296643 32113
rect 296671 32085 298728 32113
rect 298756 32085 298790 32113
rect 298818 32085 298852 32113
rect 298880 32085 298914 32113
rect 298942 32085 298990 32113
rect -958 32051 298990 32085
rect -958 32023 -910 32051
rect -882 32023 -848 32051
rect -820 32023 -786 32051
rect -758 32023 -724 32051
rect -696 32023 4617 32051
rect 4645 32023 4679 32051
rect 4707 32023 4741 32051
rect 4769 32023 4803 32051
rect 4831 32023 15939 32051
rect 15967 32023 16001 32051
rect 16029 32023 19977 32051
rect 20005 32023 20039 32051
rect 20067 32023 20101 32051
rect 20129 32023 20163 32051
rect 20191 32023 31299 32051
rect 31327 32023 31361 32051
rect 31389 32023 35337 32051
rect 35365 32023 35399 32051
rect 35427 32023 35461 32051
rect 35489 32023 35523 32051
rect 35551 32023 46659 32051
rect 46687 32023 46721 32051
rect 46749 32023 50697 32051
rect 50725 32023 50759 32051
rect 50787 32023 50821 32051
rect 50849 32023 50883 32051
rect 50911 32023 62019 32051
rect 62047 32023 62081 32051
rect 62109 32023 66057 32051
rect 66085 32023 66119 32051
rect 66147 32023 66181 32051
rect 66209 32023 66243 32051
rect 66271 32023 77379 32051
rect 77407 32023 77441 32051
rect 77469 32023 81417 32051
rect 81445 32023 81479 32051
rect 81507 32023 81541 32051
rect 81569 32023 81603 32051
rect 81631 32023 92739 32051
rect 92767 32023 92801 32051
rect 92829 32023 96777 32051
rect 96805 32023 96839 32051
rect 96867 32023 96901 32051
rect 96929 32023 96963 32051
rect 96991 32023 108099 32051
rect 108127 32023 108161 32051
rect 108189 32023 112137 32051
rect 112165 32023 112199 32051
rect 112227 32023 112261 32051
rect 112289 32023 112323 32051
rect 112351 32023 123459 32051
rect 123487 32023 123521 32051
rect 123549 32023 127497 32051
rect 127525 32023 127559 32051
rect 127587 32023 127621 32051
rect 127649 32023 127683 32051
rect 127711 32023 138819 32051
rect 138847 32023 138881 32051
rect 138909 32023 142857 32051
rect 142885 32023 142919 32051
rect 142947 32023 142981 32051
rect 143009 32023 143043 32051
rect 143071 32023 154179 32051
rect 154207 32023 154241 32051
rect 154269 32023 158217 32051
rect 158245 32023 158279 32051
rect 158307 32023 158341 32051
rect 158369 32023 158403 32051
rect 158431 32023 169539 32051
rect 169567 32023 169601 32051
rect 169629 32023 173577 32051
rect 173605 32023 173639 32051
rect 173667 32023 173701 32051
rect 173729 32023 173763 32051
rect 173791 32023 184899 32051
rect 184927 32023 184961 32051
rect 184989 32023 188937 32051
rect 188965 32023 188999 32051
rect 189027 32023 189061 32051
rect 189089 32023 189123 32051
rect 189151 32023 200259 32051
rect 200287 32023 200321 32051
rect 200349 32023 204297 32051
rect 204325 32023 204359 32051
rect 204387 32023 204421 32051
rect 204449 32023 204483 32051
rect 204511 32023 215619 32051
rect 215647 32023 215681 32051
rect 215709 32023 219657 32051
rect 219685 32023 219719 32051
rect 219747 32023 219781 32051
rect 219809 32023 219843 32051
rect 219871 32023 230979 32051
rect 231007 32023 231041 32051
rect 231069 32023 235017 32051
rect 235045 32023 235079 32051
rect 235107 32023 235141 32051
rect 235169 32023 235203 32051
rect 235231 32023 246339 32051
rect 246367 32023 246401 32051
rect 246429 32023 250377 32051
rect 250405 32023 250439 32051
rect 250467 32023 250501 32051
rect 250529 32023 250563 32051
rect 250591 32023 261699 32051
rect 261727 32023 261761 32051
rect 261789 32023 265737 32051
rect 265765 32023 265799 32051
rect 265827 32023 265861 32051
rect 265889 32023 265923 32051
rect 265951 32023 277059 32051
rect 277087 32023 277121 32051
rect 277149 32023 281097 32051
rect 281125 32023 281159 32051
rect 281187 32023 281221 32051
rect 281249 32023 281283 32051
rect 281311 32023 296457 32051
rect 296485 32023 296519 32051
rect 296547 32023 296581 32051
rect 296609 32023 296643 32051
rect 296671 32023 298728 32051
rect 298756 32023 298790 32051
rect 298818 32023 298852 32051
rect 298880 32023 298914 32051
rect 298942 32023 298990 32051
rect -958 31989 298990 32023
rect -958 31961 -910 31989
rect -882 31961 -848 31989
rect -820 31961 -786 31989
rect -758 31961 -724 31989
rect -696 31961 4617 31989
rect 4645 31961 4679 31989
rect 4707 31961 4741 31989
rect 4769 31961 4803 31989
rect 4831 31961 15939 31989
rect 15967 31961 16001 31989
rect 16029 31961 19977 31989
rect 20005 31961 20039 31989
rect 20067 31961 20101 31989
rect 20129 31961 20163 31989
rect 20191 31961 31299 31989
rect 31327 31961 31361 31989
rect 31389 31961 35337 31989
rect 35365 31961 35399 31989
rect 35427 31961 35461 31989
rect 35489 31961 35523 31989
rect 35551 31961 46659 31989
rect 46687 31961 46721 31989
rect 46749 31961 50697 31989
rect 50725 31961 50759 31989
rect 50787 31961 50821 31989
rect 50849 31961 50883 31989
rect 50911 31961 62019 31989
rect 62047 31961 62081 31989
rect 62109 31961 66057 31989
rect 66085 31961 66119 31989
rect 66147 31961 66181 31989
rect 66209 31961 66243 31989
rect 66271 31961 77379 31989
rect 77407 31961 77441 31989
rect 77469 31961 81417 31989
rect 81445 31961 81479 31989
rect 81507 31961 81541 31989
rect 81569 31961 81603 31989
rect 81631 31961 92739 31989
rect 92767 31961 92801 31989
rect 92829 31961 96777 31989
rect 96805 31961 96839 31989
rect 96867 31961 96901 31989
rect 96929 31961 96963 31989
rect 96991 31961 108099 31989
rect 108127 31961 108161 31989
rect 108189 31961 112137 31989
rect 112165 31961 112199 31989
rect 112227 31961 112261 31989
rect 112289 31961 112323 31989
rect 112351 31961 123459 31989
rect 123487 31961 123521 31989
rect 123549 31961 127497 31989
rect 127525 31961 127559 31989
rect 127587 31961 127621 31989
rect 127649 31961 127683 31989
rect 127711 31961 138819 31989
rect 138847 31961 138881 31989
rect 138909 31961 142857 31989
rect 142885 31961 142919 31989
rect 142947 31961 142981 31989
rect 143009 31961 143043 31989
rect 143071 31961 154179 31989
rect 154207 31961 154241 31989
rect 154269 31961 158217 31989
rect 158245 31961 158279 31989
rect 158307 31961 158341 31989
rect 158369 31961 158403 31989
rect 158431 31961 169539 31989
rect 169567 31961 169601 31989
rect 169629 31961 173577 31989
rect 173605 31961 173639 31989
rect 173667 31961 173701 31989
rect 173729 31961 173763 31989
rect 173791 31961 184899 31989
rect 184927 31961 184961 31989
rect 184989 31961 188937 31989
rect 188965 31961 188999 31989
rect 189027 31961 189061 31989
rect 189089 31961 189123 31989
rect 189151 31961 200259 31989
rect 200287 31961 200321 31989
rect 200349 31961 204297 31989
rect 204325 31961 204359 31989
rect 204387 31961 204421 31989
rect 204449 31961 204483 31989
rect 204511 31961 215619 31989
rect 215647 31961 215681 31989
rect 215709 31961 219657 31989
rect 219685 31961 219719 31989
rect 219747 31961 219781 31989
rect 219809 31961 219843 31989
rect 219871 31961 230979 31989
rect 231007 31961 231041 31989
rect 231069 31961 235017 31989
rect 235045 31961 235079 31989
rect 235107 31961 235141 31989
rect 235169 31961 235203 31989
rect 235231 31961 246339 31989
rect 246367 31961 246401 31989
rect 246429 31961 250377 31989
rect 250405 31961 250439 31989
rect 250467 31961 250501 31989
rect 250529 31961 250563 31989
rect 250591 31961 261699 31989
rect 261727 31961 261761 31989
rect 261789 31961 265737 31989
rect 265765 31961 265799 31989
rect 265827 31961 265861 31989
rect 265889 31961 265923 31989
rect 265951 31961 277059 31989
rect 277087 31961 277121 31989
rect 277149 31961 281097 31989
rect 281125 31961 281159 31989
rect 281187 31961 281221 31989
rect 281249 31961 281283 31989
rect 281311 31961 296457 31989
rect 296485 31961 296519 31989
rect 296547 31961 296581 31989
rect 296609 31961 296643 31989
rect 296671 31961 298728 31989
rect 298756 31961 298790 31989
rect 298818 31961 298852 31989
rect 298880 31961 298914 31989
rect 298942 31961 298990 31989
rect -958 31913 298990 31961
rect -958 29175 298990 29223
rect -958 29147 -430 29175
rect -402 29147 -368 29175
rect -340 29147 -306 29175
rect -278 29147 -244 29175
rect -216 29147 2757 29175
rect 2785 29147 2819 29175
rect 2847 29147 2881 29175
rect 2909 29147 2943 29175
rect 2971 29147 8259 29175
rect 8287 29147 8321 29175
rect 8349 29147 18117 29175
rect 18145 29147 18179 29175
rect 18207 29147 18241 29175
rect 18269 29147 18303 29175
rect 18331 29147 23619 29175
rect 23647 29147 23681 29175
rect 23709 29147 33477 29175
rect 33505 29147 33539 29175
rect 33567 29147 33601 29175
rect 33629 29147 33663 29175
rect 33691 29147 38979 29175
rect 39007 29147 39041 29175
rect 39069 29147 48837 29175
rect 48865 29147 48899 29175
rect 48927 29147 48961 29175
rect 48989 29147 49023 29175
rect 49051 29147 54339 29175
rect 54367 29147 54401 29175
rect 54429 29147 64197 29175
rect 64225 29147 64259 29175
rect 64287 29147 64321 29175
rect 64349 29147 64383 29175
rect 64411 29147 69699 29175
rect 69727 29147 69761 29175
rect 69789 29147 79557 29175
rect 79585 29147 79619 29175
rect 79647 29147 79681 29175
rect 79709 29147 79743 29175
rect 79771 29147 85059 29175
rect 85087 29147 85121 29175
rect 85149 29147 94917 29175
rect 94945 29147 94979 29175
rect 95007 29147 95041 29175
rect 95069 29147 95103 29175
rect 95131 29147 100419 29175
rect 100447 29147 100481 29175
rect 100509 29147 110277 29175
rect 110305 29147 110339 29175
rect 110367 29147 110401 29175
rect 110429 29147 110463 29175
rect 110491 29147 115779 29175
rect 115807 29147 115841 29175
rect 115869 29147 125637 29175
rect 125665 29147 125699 29175
rect 125727 29147 125761 29175
rect 125789 29147 125823 29175
rect 125851 29147 131139 29175
rect 131167 29147 131201 29175
rect 131229 29147 140997 29175
rect 141025 29147 141059 29175
rect 141087 29147 141121 29175
rect 141149 29147 141183 29175
rect 141211 29147 146499 29175
rect 146527 29147 146561 29175
rect 146589 29147 156357 29175
rect 156385 29147 156419 29175
rect 156447 29147 156481 29175
rect 156509 29147 156543 29175
rect 156571 29147 161859 29175
rect 161887 29147 161921 29175
rect 161949 29147 171717 29175
rect 171745 29147 171779 29175
rect 171807 29147 171841 29175
rect 171869 29147 171903 29175
rect 171931 29147 177219 29175
rect 177247 29147 177281 29175
rect 177309 29147 187077 29175
rect 187105 29147 187139 29175
rect 187167 29147 187201 29175
rect 187229 29147 187263 29175
rect 187291 29147 192579 29175
rect 192607 29147 192641 29175
rect 192669 29147 202437 29175
rect 202465 29147 202499 29175
rect 202527 29147 202561 29175
rect 202589 29147 202623 29175
rect 202651 29147 207939 29175
rect 207967 29147 208001 29175
rect 208029 29147 217797 29175
rect 217825 29147 217859 29175
rect 217887 29147 217921 29175
rect 217949 29147 217983 29175
rect 218011 29147 223299 29175
rect 223327 29147 223361 29175
rect 223389 29147 233157 29175
rect 233185 29147 233219 29175
rect 233247 29147 233281 29175
rect 233309 29147 233343 29175
rect 233371 29147 238659 29175
rect 238687 29147 238721 29175
rect 238749 29147 248517 29175
rect 248545 29147 248579 29175
rect 248607 29147 248641 29175
rect 248669 29147 248703 29175
rect 248731 29147 254019 29175
rect 254047 29147 254081 29175
rect 254109 29147 263877 29175
rect 263905 29147 263939 29175
rect 263967 29147 264001 29175
rect 264029 29147 264063 29175
rect 264091 29147 269379 29175
rect 269407 29147 269441 29175
rect 269469 29147 279237 29175
rect 279265 29147 279299 29175
rect 279327 29147 279361 29175
rect 279389 29147 279423 29175
rect 279451 29147 284739 29175
rect 284767 29147 284801 29175
rect 284829 29147 294597 29175
rect 294625 29147 294659 29175
rect 294687 29147 294721 29175
rect 294749 29147 294783 29175
rect 294811 29147 298248 29175
rect 298276 29147 298310 29175
rect 298338 29147 298372 29175
rect 298400 29147 298434 29175
rect 298462 29147 298990 29175
rect -958 29113 298990 29147
rect -958 29085 -430 29113
rect -402 29085 -368 29113
rect -340 29085 -306 29113
rect -278 29085 -244 29113
rect -216 29085 2757 29113
rect 2785 29085 2819 29113
rect 2847 29085 2881 29113
rect 2909 29085 2943 29113
rect 2971 29085 8259 29113
rect 8287 29085 8321 29113
rect 8349 29085 18117 29113
rect 18145 29085 18179 29113
rect 18207 29085 18241 29113
rect 18269 29085 18303 29113
rect 18331 29085 23619 29113
rect 23647 29085 23681 29113
rect 23709 29085 33477 29113
rect 33505 29085 33539 29113
rect 33567 29085 33601 29113
rect 33629 29085 33663 29113
rect 33691 29085 38979 29113
rect 39007 29085 39041 29113
rect 39069 29085 48837 29113
rect 48865 29085 48899 29113
rect 48927 29085 48961 29113
rect 48989 29085 49023 29113
rect 49051 29085 54339 29113
rect 54367 29085 54401 29113
rect 54429 29085 64197 29113
rect 64225 29085 64259 29113
rect 64287 29085 64321 29113
rect 64349 29085 64383 29113
rect 64411 29085 69699 29113
rect 69727 29085 69761 29113
rect 69789 29085 79557 29113
rect 79585 29085 79619 29113
rect 79647 29085 79681 29113
rect 79709 29085 79743 29113
rect 79771 29085 85059 29113
rect 85087 29085 85121 29113
rect 85149 29085 94917 29113
rect 94945 29085 94979 29113
rect 95007 29085 95041 29113
rect 95069 29085 95103 29113
rect 95131 29085 100419 29113
rect 100447 29085 100481 29113
rect 100509 29085 110277 29113
rect 110305 29085 110339 29113
rect 110367 29085 110401 29113
rect 110429 29085 110463 29113
rect 110491 29085 115779 29113
rect 115807 29085 115841 29113
rect 115869 29085 125637 29113
rect 125665 29085 125699 29113
rect 125727 29085 125761 29113
rect 125789 29085 125823 29113
rect 125851 29085 131139 29113
rect 131167 29085 131201 29113
rect 131229 29085 140997 29113
rect 141025 29085 141059 29113
rect 141087 29085 141121 29113
rect 141149 29085 141183 29113
rect 141211 29085 146499 29113
rect 146527 29085 146561 29113
rect 146589 29085 156357 29113
rect 156385 29085 156419 29113
rect 156447 29085 156481 29113
rect 156509 29085 156543 29113
rect 156571 29085 161859 29113
rect 161887 29085 161921 29113
rect 161949 29085 171717 29113
rect 171745 29085 171779 29113
rect 171807 29085 171841 29113
rect 171869 29085 171903 29113
rect 171931 29085 177219 29113
rect 177247 29085 177281 29113
rect 177309 29085 187077 29113
rect 187105 29085 187139 29113
rect 187167 29085 187201 29113
rect 187229 29085 187263 29113
rect 187291 29085 192579 29113
rect 192607 29085 192641 29113
rect 192669 29085 202437 29113
rect 202465 29085 202499 29113
rect 202527 29085 202561 29113
rect 202589 29085 202623 29113
rect 202651 29085 207939 29113
rect 207967 29085 208001 29113
rect 208029 29085 217797 29113
rect 217825 29085 217859 29113
rect 217887 29085 217921 29113
rect 217949 29085 217983 29113
rect 218011 29085 223299 29113
rect 223327 29085 223361 29113
rect 223389 29085 233157 29113
rect 233185 29085 233219 29113
rect 233247 29085 233281 29113
rect 233309 29085 233343 29113
rect 233371 29085 238659 29113
rect 238687 29085 238721 29113
rect 238749 29085 248517 29113
rect 248545 29085 248579 29113
rect 248607 29085 248641 29113
rect 248669 29085 248703 29113
rect 248731 29085 254019 29113
rect 254047 29085 254081 29113
rect 254109 29085 263877 29113
rect 263905 29085 263939 29113
rect 263967 29085 264001 29113
rect 264029 29085 264063 29113
rect 264091 29085 269379 29113
rect 269407 29085 269441 29113
rect 269469 29085 279237 29113
rect 279265 29085 279299 29113
rect 279327 29085 279361 29113
rect 279389 29085 279423 29113
rect 279451 29085 284739 29113
rect 284767 29085 284801 29113
rect 284829 29085 294597 29113
rect 294625 29085 294659 29113
rect 294687 29085 294721 29113
rect 294749 29085 294783 29113
rect 294811 29085 298248 29113
rect 298276 29085 298310 29113
rect 298338 29085 298372 29113
rect 298400 29085 298434 29113
rect 298462 29085 298990 29113
rect -958 29051 298990 29085
rect -958 29023 -430 29051
rect -402 29023 -368 29051
rect -340 29023 -306 29051
rect -278 29023 -244 29051
rect -216 29023 2757 29051
rect 2785 29023 2819 29051
rect 2847 29023 2881 29051
rect 2909 29023 2943 29051
rect 2971 29023 8259 29051
rect 8287 29023 8321 29051
rect 8349 29023 18117 29051
rect 18145 29023 18179 29051
rect 18207 29023 18241 29051
rect 18269 29023 18303 29051
rect 18331 29023 23619 29051
rect 23647 29023 23681 29051
rect 23709 29023 33477 29051
rect 33505 29023 33539 29051
rect 33567 29023 33601 29051
rect 33629 29023 33663 29051
rect 33691 29023 38979 29051
rect 39007 29023 39041 29051
rect 39069 29023 48837 29051
rect 48865 29023 48899 29051
rect 48927 29023 48961 29051
rect 48989 29023 49023 29051
rect 49051 29023 54339 29051
rect 54367 29023 54401 29051
rect 54429 29023 64197 29051
rect 64225 29023 64259 29051
rect 64287 29023 64321 29051
rect 64349 29023 64383 29051
rect 64411 29023 69699 29051
rect 69727 29023 69761 29051
rect 69789 29023 79557 29051
rect 79585 29023 79619 29051
rect 79647 29023 79681 29051
rect 79709 29023 79743 29051
rect 79771 29023 85059 29051
rect 85087 29023 85121 29051
rect 85149 29023 94917 29051
rect 94945 29023 94979 29051
rect 95007 29023 95041 29051
rect 95069 29023 95103 29051
rect 95131 29023 100419 29051
rect 100447 29023 100481 29051
rect 100509 29023 110277 29051
rect 110305 29023 110339 29051
rect 110367 29023 110401 29051
rect 110429 29023 110463 29051
rect 110491 29023 115779 29051
rect 115807 29023 115841 29051
rect 115869 29023 125637 29051
rect 125665 29023 125699 29051
rect 125727 29023 125761 29051
rect 125789 29023 125823 29051
rect 125851 29023 131139 29051
rect 131167 29023 131201 29051
rect 131229 29023 140997 29051
rect 141025 29023 141059 29051
rect 141087 29023 141121 29051
rect 141149 29023 141183 29051
rect 141211 29023 146499 29051
rect 146527 29023 146561 29051
rect 146589 29023 156357 29051
rect 156385 29023 156419 29051
rect 156447 29023 156481 29051
rect 156509 29023 156543 29051
rect 156571 29023 161859 29051
rect 161887 29023 161921 29051
rect 161949 29023 171717 29051
rect 171745 29023 171779 29051
rect 171807 29023 171841 29051
rect 171869 29023 171903 29051
rect 171931 29023 177219 29051
rect 177247 29023 177281 29051
rect 177309 29023 187077 29051
rect 187105 29023 187139 29051
rect 187167 29023 187201 29051
rect 187229 29023 187263 29051
rect 187291 29023 192579 29051
rect 192607 29023 192641 29051
rect 192669 29023 202437 29051
rect 202465 29023 202499 29051
rect 202527 29023 202561 29051
rect 202589 29023 202623 29051
rect 202651 29023 207939 29051
rect 207967 29023 208001 29051
rect 208029 29023 217797 29051
rect 217825 29023 217859 29051
rect 217887 29023 217921 29051
rect 217949 29023 217983 29051
rect 218011 29023 223299 29051
rect 223327 29023 223361 29051
rect 223389 29023 233157 29051
rect 233185 29023 233219 29051
rect 233247 29023 233281 29051
rect 233309 29023 233343 29051
rect 233371 29023 238659 29051
rect 238687 29023 238721 29051
rect 238749 29023 248517 29051
rect 248545 29023 248579 29051
rect 248607 29023 248641 29051
rect 248669 29023 248703 29051
rect 248731 29023 254019 29051
rect 254047 29023 254081 29051
rect 254109 29023 263877 29051
rect 263905 29023 263939 29051
rect 263967 29023 264001 29051
rect 264029 29023 264063 29051
rect 264091 29023 269379 29051
rect 269407 29023 269441 29051
rect 269469 29023 279237 29051
rect 279265 29023 279299 29051
rect 279327 29023 279361 29051
rect 279389 29023 279423 29051
rect 279451 29023 284739 29051
rect 284767 29023 284801 29051
rect 284829 29023 294597 29051
rect 294625 29023 294659 29051
rect 294687 29023 294721 29051
rect 294749 29023 294783 29051
rect 294811 29023 298248 29051
rect 298276 29023 298310 29051
rect 298338 29023 298372 29051
rect 298400 29023 298434 29051
rect 298462 29023 298990 29051
rect -958 28989 298990 29023
rect -958 28961 -430 28989
rect -402 28961 -368 28989
rect -340 28961 -306 28989
rect -278 28961 -244 28989
rect -216 28961 2757 28989
rect 2785 28961 2819 28989
rect 2847 28961 2881 28989
rect 2909 28961 2943 28989
rect 2971 28961 8259 28989
rect 8287 28961 8321 28989
rect 8349 28961 18117 28989
rect 18145 28961 18179 28989
rect 18207 28961 18241 28989
rect 18269 28961 18303 28989
rect 18331 28961 23619 28989
rect 23647 28961 23681 28989
rect 23709 28961 33477 28989
rect 33505 28961 33539 28989
rect 33567 28961 33601 28989
rect 33629 28961 33663 28989
rect 33691 28961 38979 28989
rect 39007 28961 39041 28989
rect 39069 28961 48837 28989
rect 48865 28961 48899 28989
rect 48927 28961 48961 28989
rect 48989 28961 49023 28989
rect 49051 28961 54339 28989
rect 54367 28961 54401 28989
rect 54429 28961 64197 28989
rect 64225 28961 64259 28989
rect 64287 28961 64321 28989
rect 64349 28961 64383 28989
rect 64411 28961 69699 28989
rect 69727 28961 69761 28989
rect 69789 28961 79557 28989
rect 79585 28961 79619 28989
rect 79647 28961 79681 28989
rect 79709 28961 79743 28989
rect 79771 28961 85059 28989
rect 85087 28961 85121 28989
rect 85149 28961 94917 28989
rect 94945 28961 94979 28989
rect 95007 28961 95041 28989
rect 95069 28961 95103 28989
rect 95131 28961 100419 28989
rect 100447 28961 100481 28989
rect 100509 28961 110277 28989
rect 110305 28961 110339 28989
rect 110367 28961 110401 28989
rect 110429 28961 110463 28989
rect 110491 28961 115779 28989
rect 115807 28961 115841 28989
rect 115869 28961 125637 28989
rect 125665 28961 125699 28989
rect 125727 28961 125761 28989
rect 125789 28961 125823 28989
rect 125851 28961 131139 28989
rect 131167 28961 131201 28989
rect 131229 28961 140997 28989
rect 141025 28961 141059 28989
rect 141087 28961 141121 28989
rect 141149 28961 141183 28989
rect 141211 28961 146499 28989
rect 146527 28961 146561 28989
rect 146589 28961 156357 28989
rect 156385 28961 156419 28989
rect 156447 28961 156481 28989
rect 156509 28961 156543 28989
rect 156571 28961 161859 28989
rect 161887 28961 161921 28989
rect 161949 28961 171717 28989
rect 171745 28961 171779 28989
rect 171807 28961 171841 28989
rect 171869 28961 171903 28989
rect 171931 28961 177219 28989
rect 177247 28961 177281 28989
rect 177309 28961 187077 28989
rect 187105 28961 187139 28989
rect 187167 28961 187201 28989
rect 187229 28961 187263 28989
rect 187291 28961 192579 28989
rect 192607 28961 192641 28989
rect 192669 28961 202437 28989
rect 202465 28961 202499 28989
rect 202527 28961 202561 28989
rect 202589 28961 202623 28989
rect 202651 28961 207939 28989
rect 207967 28961 208001 28989
rect 208029 28961 217797 28989
rect 217825 28961 217859 28989
rect 217887 28961 217921 28989
rect 217949 28961 217983 28989
rect 218011 28961 223299 28989
rect 223327 28961 223361 28989
rect 223389 28961 233157 28989
rect 233185 28961 233219 28989
rect 233247 28961 233281 28989
rect 233309 28961 233343 28989
rect 233371 28961 238659 28989
rect 238687 28961 238721 28989
rect 238749 28961 248517 28989
rect 248545 28961 248579 28989
rect 248607 28961 248641 28989
rect 248669 28961 248703 28989
rect 248731 28961 254019 28989
rect 254047 28961 254081 28989
rect 254109 28961 263877 28989
rect 263905 28961 263939 28989
rect 263967 28961 264001 28989
rect 264029 28961 264063 28989
rect 264091 28961 269379 28989
rect 269407 28961 269441 28989
rect 269469 28961 279237 28989
rect 279265 28961 279299 28989
rect 279327 28961 279361 28989
rect 279389 28961 279423 28989
rect 279451 28961 284739 28989
rect 284767 28961 284801 28989
rect 284829 28961 294597 28989
rect 294625 28961 294659 28989
rect 294687 28961 294721 28989
rect 294749 28961 294783 28989
rect 294811 28961 298248 28989
rect 298276 28961 298310 28989
rect 298338 28961 298372 28989
rect 298400 28961 298434 28989
rect 298462 28961 298990 28989
rect -958 28913 298990 28961
rect -958 23175 298990 23223
rect -958 23147 -910 23175
rect -882 23147 -848 23175
rect -820 23147 -786 23175
rect -758 23147 -724 23175
rect -696 23147 4617 23175
rect 4645 23147 4679 23175
rect 4707 23147 4741 23175
rect 4769 23147 4803 23175
rect 4831 23147 15939 23175
rect 15967 23147 16001 23175
rect 16029 23147 19977 23175
rect 20005 23147 20039 23175
rect 20067 23147 20101 23175
rect 20129 23147 20163 23175
rect 20191 23147 31299 23175
rect 31327 23147 31361 23175
rect 31389 23147 35337 23175
rect 35365 23147 35399 23175
rect 35427 23147 35461 23175
rect 35489 23147 35523 23175
rect 35551 23147 46659 23175
rect 46687 23147 46721 23175
rect 46749 23147 50697 23175
rect 50725 23147 50759 23175
rect 50787 23147 50821 23175
rect 50849 23147 50883 23175
rect 50911 23147 62019 23175
rect 62047 23147 62081 23175
rect 62109 23147 66057 23175
rect 66085 23147 66119 23175
rect 66147 23147 66181 23175
rect 66209 23147 66243 23175
rect 66271 23147 77379 23175
rect 77407 23147 77441 23175
rect 77469 23147 81417 23175
rect 81445 23147 81479 23175
rect 81507 23147 81541 23175
rect 81569 23147 81603 23175
rect 81631 23147 92739 23175
rect 92767 23147 92801 23175
rect 92829 23147 96777 23175
rect 96805 23147 96839 23175
rect 96867 23147 96901 23175
rect 96929 23147 96963 23175
rect 96991 23147 108099 23175
rect 108127 23147 108161 23175
rect 108189 23147 112137 23175
rect 112165 23147 112199 23175
rect 112227 23147 112261 23175
rect 112289 23147 112323 23175
rect 112351 23147 123459 23175
rect 123487 23147 123521 23175
rect 123549 23147 127497 23175
rect 127525 23147 127559 23175
rect 127587 23147 127621 23175
rect 127649 23147 127683 23175
rect 127711 23147 138819 23175
rect 138847 23147 138881 23175
rect 138909 23147 142857 23175
rect 142885 23147 142919 23175
rect 142947 23147 142981 23175
rect 143009 23147 143043 23175
rect 143071 23147 154179 23175
rect 154207 23147 154241 23175
rect 154269 23147 158217 23175
rect 158245 23147 158279 23175
rect 158307 23147 158341 23175
rect 158369 23147 158403 23175
rect 158431 23147 169539 23175
rect 169567 23147 169601 23175
rect 169629 23147 173577 23175
rect 173605 23147 173639 23175
rect 173667 23147 173701 23175
rect 173729 23147 173763 23175
rect 173791 23147 184899 23175
rect 184927 23147 184961 23175
rect 184989 23147 188937 23175
rect 188965 23147 188999 23175
rect 189027 23147 189061 23175
rect 189089 23147 189123 23175
rect 189151 23147 200259 23175
rect 200287 23147 200321 23175
rect 200349 23147 204297 23175
rect 204325 23147 204359 23175
rect 204387 23147 204421 23175
rect 204449 23147 204483 23175
rect 204511 23147 215619 23175
rect 215647 23147 215681 23175
rect 215709 23147 219657 23175
rect 219685 23147 219719 23175
rect 219747 23147 219781 23175
rect 219809 23147 219843 23175
rect 219871 23147 230979 23175
rect 231007 23147 231041 23175
rect 231069 23147 235017 23175
rect 235045 23147 235079 23175
rect 235107 23147 235141 23175
rect 235169 23147 235203 23175
rect 235231 23147 246339 23175
rect 246367 23147 246401 23175
rect 246429 23147 250377 23175
rect 250405 23147 250439 23175
rect 250467 23147 250501 23175
rect 250529 23147 250563 23175
rect 250591 23147 261699 23175
rect 261727 23147 261761 23175
rect 261789 23147 265737 23175
rect 265765 23147 265799 23175
rect 265827 23147 265861 23175
rect 265889 23147 265923 23175
rect 265951 23147 277059 23175
rect 277087 23147 277121 23175
rect 277149 23147 281097 23175
rect 281125 23147 281159 23175
rect 281187 23147 281221 23175
rect 281249 23147 281283 23175
rect 281311 23147 296457 23175
rect 296485 23147 296519 23175
rect 296547 23147 296581 23175
rect 296609 23147 296643 23175
rect 296671 23147 298728 23175
rect 298756 23147 298790 23175
rect 298818 23147 298852 23175
rect 298880 23147 298914 23175
rect 298942 23147 298990 23175
rect -958 23113 298990 23147
rect -958 23085 -910 23113
rect -882 23085 -848 23113
rect -820 23085 -786 23113
rect -758 23085 -724 23113
rect -696 23085 4617 23113
rect 4645 23085 4679 23113
rect 4707 23085 4741 23113
rect 4769 23085 4803 23113
rect 4831 23085 15939 23113
rect 15967 23085 16001 23113
rect 16029 23085 19977 23113
rect 20005 23085 20039 23113
rect 20067 23085 20101 23113
rect 20129 23085 20163 23113
rect 20191 23085 31299 23113
rect 31327 23085 31361 23113
rect 31389 23085 35337 23113
rect 35365 23085 35399 23113
rect 35427 23085 35461 23113
rect 35489 23085 35523 23113
rect 35551 23085 46659 23113
rect 46687 23085 46721 23113
rect 46749 23085 50697 23113
rect 50725 23085 50759 23113
rect 50787 23085 50821 23113
rect 50849 23085 50883 23113
rect 50911 23085 62019 23113
rect 62047 23085 62081 23113
rect 62109 23085 66057 23113
rect 66085 23085 66119 23113
rect 66147 23085 66181 23113
rect 66209 23085 66243 23113
rect 66271 23085 77379 23113
rect 77407 23085 77441 23113
rect 77469 23085 81417 23113
rect 81445 23085 81479 23113
rect 81507 23085 81541 23113
rect 81569 23085 81603 23113
rect 81631 23085 92739 23113
rect 92767 23085 92801 23113
rect 92829 23085 96777 23113
rect 96805 23085 96839 23113
rect 96867 23085 96901 23113
rect 96929 23085 96963 23113
rect 96991 23085 108099 23113
rect 108127 23085 108161 23113
rect 108189 23085 112137 23113
rect 112165 23085 112199 23113
rect 112227 23085 112261 23113
rect 112289 23085 112323 23113
rect 112351 23085 123459 23113
rect 123487 23085 123521 23113
rect 123549 23085 127497 23113
rect 127525 23085 127559 23113
rect 127587 23085 127621 23113
rect 127649 23085 127683 23113
rect 127711 23085 138819 23113
rect 138847 23085 138881 23113
rect 138909 23085 142857 23113
rect 142885 23085 142919 23113
rect 142947 23085 142981 23113
rect 143009 23085 143043 23113
rect 143071 23085 154179 23113
rect 154207 23085 154241 23113
rect 154269 23085 158217 23113
rect 158245 23085 158279 23113
rect 158307 23085 158341 23113
rect 158369 23085 158403 23113
rect 158431 23085 169539 23113
rect 169567 23085 169601 23113
rect 169629 23085 173577 23113
rect 173605 23085 173639 23113
rect 173667 23085 173701 23113
rect 173729 23085 173763 23113
rect 173791 23085 184899 23113
rect 184927 23085 184961 23113
rect 184989 23085 188937 23113
rect 188965 23085 188999 23113
rect 189027 23085 189061 23113
rect 189089 23085 189123 23113
rect 189151 23085 200259 23113
rect 200287 23085 200321 23113
rect 200349 23085 204297 23113
rect 204325 23085 204359 23113
rect 204387 23085 204421 23113
rect 204449 23085 204483 23113
rect 204511 23085 215619 23113
rect 215647 23085 215681 23113
rect 215709 23085 219657 23113
rect 219685 23085 219719 23113
rect 219747 23085 219781 23113
rect 219809 23085 219843 23113
rect 219871 23085 230979 23113
rect 231007 23085 231041 23113
rect 231069 23085 235017 23113
rect 235045 23085 235079 23113
rect 235107 23085 235141 23113
rect 235169 23085 235203 23113
rect 235231 23085 246339 23113
rect 246367 23085 246401 23113
rect 246429 23085 250377 23113
rect 250405 23085 250439 23113
rect 250467 23085 250501 23113
rect 250529 23085 250563 23113
rect 250591 23085 261699 23113
rect 261727 23085 261761 23113
rect 261789 23085 265737 23113
rect 265765 23085 265799 23113
rect 265827 23085 265861 23113
rect 265889 23085 265923 23113
rect 265951 23085 277059 23113
rect 277087 23085 277121 23113
rect 277149 23085 281097 23113
rect 281125 23085 281159 23113
rect 281187 23085 281221 23113
rect 281249 23085 281283 23113
rect 281311 23085 296457 23113
rect 296485 23085 296519 23113
rect 296547 23085 296581 23113
rect 296609 23085 296643 23113
rect 296671 23085 298728 23113
rect 298756 23085 298790 23113
rect 298818 23085 298852 23113
rect 298880 23085 298914 23113
rect 298942 23085 298990 23113
rect -958 23051 298990 23085
rect -958 23023 -910 23051
rect -882 23023 -848 23051
rect -820 23023 -786 23051
rect -758 23023 -724 23051
rect -696 23023 4617 23051
rect 4645 23023 4679 23051
rect 4707 23023 4741 23051
rect 4769 23023 4803 23051
rect 4831 23023 15939 23051
rect 15967 23023 16001 23051
rect 16029 23023 19977 23051
rect 20005 23023 20039 23051
rect 20067 23023 20101 23051
rect 20129 23023 20163 23051
rect 20191 23023 31299 23051
rect 31327 23023 31361 23051
rect 31389 23023 35337 23051
rect 35365 23023 35399 23051
rect 35427 23023 35461 23051
rect 35489 23023 35523 23051
rect 35551 23023 46659 23051
rect 46687 23023 46721 23051
rect 46749 23023 50697 23051
rect 50725 23023 50759 23051
rect 50787 23023 50821 23051
rect 50849 23023 50883 23051
rect 50911 23023 62019 23051
rect 62047 23023 62081 23051
rect 62109 23023 66057 23051
rect 66085 23023 66119 23051
rect 66147 23023 66181 23051
rect 66209 23023 66243 23051
rect 66271 23023 77379 23051
rect 77407 23023 77441 23051
rect 77469 23023 81417 23051
rect 81445 23023 81479 23051
rect 81507 23023 81541 23051
rect 81569 23023 81603 23051
rect 81631 23023 92739 23051
rect 92767 23023 92801 23051
rect 92829 23023 96777 23051
rect 96805 23023 96839 23051
rect 96867 23023 96901 23051
rect 96929 23023 96963 23051
rect 96991 23023 108099 23051
rect 108127 23023 108161 23051
rect 108189 23023 112137 23051
rect 112165 23023 112199 23051
rect 112227 23023 112261 23051
rect 112289 23023 112323 23051
rect 112351 23023 123459 23051
rect 123487 23023 123521 23051
rect 123549 23023 127497 23051
rect 127525 23023 127559 23051
rect 127587 23023 127621 23051
rect 127649 23023 127683 23051
rect 127711 23023 138819 23051
rect 138847 23023 138881 23051
rect 138909 23023 142857 23051
rect 142885 23023 142919 23051
rect 142947 23023 142981 23051
rect 143009 23023 143043 23051
rect 143071 23023 154179 23051
rect 154207 23023 154241 23051
rect 154269 23023 158217 23051
rect 158245 23023 158279 23051
rect 158307 23023 158341 23051
rect 158369 23023 158403 23051
rect 158431 23023 169539 23051
rect 169567 23023 169601 23051
rect 169629 23023 173577 23051
rect 173605 23023 173639 23051
rect 173667 23023 173701 23051
rect 173729 23023 173763 23051
rect 173791 23023 184899 23051
rect 184927 23023 184961 23051
rect 184989 23023 188937 23051
rect 188965 23023 188999 23051
rect 189027 23023 189061 23051
rect 189089 23023 189123 23051
rect 189151 23023 200259 23051
rect 200287 23023 200321 23051
rect 200349 23023 204297 23051
rect 204325 23023 204359 23051
rect 204387 23023 204421 23051
rect 204449 23023 204483 23051
rect 204511 23023 215619 23051
rect 215647 23023 215681 23051
rect 215709 23023 219657 23051
rect 219685 23023 219719 23051
rect 219747 23023 219781 23051
rect 219809 23023 219843 23051
rect 219871 23023 230979 23051
rect 231007 23023 231041 23051
rect 231069 23023 235017 23051
rect 235045 23023 235079 23051
rect 235107 23023 235141 23051
rect 235169 23023 235203 23051
rect 235231 23023 246339 23051
rect 246367 23023 246401 23051
rect 246429 23023 250377 23051
rect 250405 23023 250439 23051
rect 250467 23023 250501 23051
rect 250529 23023 250563 23051
rect 250591 23023 261699 23051
rect 261727 23023 261761 23051
rect 261789 23023 265737 23051
rect 265765 23023 265799 23051
rect 265827 23023 265861 23051
rect 265889 23023 265923 23051
rect 265951 23023 277059 23051
rect 277087 23023 277121 23051
rect 277149 23023 281097 23051
rect 281125 23023 281159 23051
rect 281187 23023 281221 23051
rect 281249 23023 281283 23051
rect 281311 23023 296457 23051
rect 296485 23023 296519 23051
rect 296547 23023 296581 23051
rect 296609 23023 296643 23051
rect 296671 23023 298728 23051
rect 298756 23023 298790 23051
rect 298818 23023 298852 23051
rect 298880 23023 298914 23051
rect 298942 23023 298990 23051
rect -958 22989 298990 23023
rect -958 22961 -910 22989
rect -882 22961 -848 22989
rect -820 22961 -786 22989
rect -758 22961 -724 22989
rect -696 22961 4617 22989
rect 4645 22961 4679 22989
rect 4707 22961 4741 22989
rect 4769 22961 4803 22989
rect 4831 22961 15939 22989
rect 15967 22961 16001 22989
rect 16029 22961 19977 22989
rect 20005 22961 20039 22989
rect 20067 22961 20101 22989
rect 20129 22961 20163 22989
rect 20191 22961 31299 22989
rect 31327 22961 31361 22989
rect 31389 22961 35337 22989
rect 35365 22961 35399 22989
rect 35427 22961 35461 22989
rect 35489 22961 35523 22989
rect 35551 22961 46659 22989
rect 46687 22961 46721 22989
rect 46749 22961 50697 22989
rect 50725 22961 50759 22989
rect 50787 22961 50821 22989
rect 50849 22961 50883 22989
rect 50911 22961 62019 22989
rect 62047 22961 62081 22989
rect 62109 22961 66057 22989
rect 66085 22961 66119 22989
rect 66147 22961 66181 22989
rect 66209 22961 66243 22989
rect 66271 22961 77379 22989
rect 77407 22961 77441 22989
rect 77469 22961 81417 22989
rect 81445 22961 81479 22989
rect 81507 22961 81541 22989
rect 81569 22961 81603 22989
rect 81631 22961 92739 22989
rect 92767 22961 92801 22989
rect 92829 22961 96777 22989
rect 96805 22961 96839 22989
rect 96867 22961 96901 22989
rect 96929 22961 96963 22989
rect 96991 22961 108099 22989
rect 108127 22961 108161 22989
rect 108189 22961 112137 22989
rect 112165 22961 112199 22989
rect 112227 22961 112261 22989
rect 112289 22961 112323 22989
rect 112351 22961 123459 22989
rect 123487 22961 123521 22989
rect 123549 22961 127497 22989
rect 127525 22961 127559 22989
rect 127587 22961 127621 22989
rect 127649 22961 127683 22989
rect 127711 22961 138819 22989
rect 138847 22961 138881 22989
rect 138909 22961 142857 22989
rect 142885 22961 142919 22989
rect 142947 22961 142981 22989
rect 143009 22961 143043 22989
rect 143071 22961 154179 22989
rect 154207 22961 154241 22989
rect 154269 22961 158217 22989
rect 158245 22961 158279 22989
rect 158307 22961 158341 22989
rect 158369 22961 158403 22989
rect 158431 22961 169539 22989
rect 169567 22961 169601 22989
rect 169629 22961 173577 22989
rect 173605 22961 173639 22989
rect 173667 22961 173701 22989
rect 173729 22961 173763 22989
rect 173791 22961 184899 22989
rect 184927 22961 184961 22989
rect 184989 22961 188937 22989
rect 188965 22961 188999 22989
rect 189027 22961 189061 22989
rect 189089 22961 189123 22989
rect 189151 22961 200259 22989
rect 200287 22961 200321 22989
rect 200349 22961 204297 22989
rect 204325 22961 204359 22989
rect 204387 22961 204421 22989
rect 204449 22961 204483 22989
rect 204511 22961 215619 22989
rect 215647 22961 215681 22989
rect 215709 22961 219657 22989
rect 219685 22961 219719 22989
rect 219747 22961 219781 22989
rect 219809 22961 219843 22989
rect 219871 22961 230979 22989
rect 231007 22961 231041 22989
rect 231069 22961 235017 22989
rect 235045 22961 235079 22989
rect 235107 22961 235141 22989
rect 235169 22961 235203 22989
rect 235231 22961 246339 22989
rect 246367 22961 246401 22989
rect 246429 22961 250377 22989
rect 250405 22961 250439 22989
rect 250467 22961 250501 22989
rect 250529 22961 250563 22989
rect 250591 22961 261699 22989
rect 261727 22961 261761 22989
rect 261789 22961 265737 22989
rect 265765 22961 265799 22989
rect 265827 22961 265861 22989
rect 265889 22961 265923 22989
rect 265951 22961 277059 22989
rect 277087 22961 277121 22989
rect 277149 22961 281097 22989
rect 281125 22961 281159 22989
rect 281187 22961 281221 22989
rect 281249 22961 281283 22989
rect 281311 22961 296457 22989
rect 296485 22961 296519 22989
rect 296547 22961 296581 22989
rect 296609 22961 296643 22989
rect 296671 22961 298728 22989
rect 298756 22961 298790 22989
rect 298818 22961 298852 22989
rect 298880 22961 298914 22989
rect 298942 22961 298990 22989
rect -958 22913 298990 22961
rect -958 20175 298990 20223
rect -958 20147 -430 20175
rect -402 20147 -368 20175
rect -340 20147 -306 20175
rect -278 20147 -244 20175
rect -216 20147 2757 20175
rect 2785 20147 2819 20175
rect 2847 20147 2881 20175
rect 2909 20147 2943 20175
rect 2971 20147 8259 20175
rect 8287 20147 8321 20175
rect 8349 20147 18117 20175
rect 18145 20147 18179 20175
rect 18207 20147 18241 20175
rect 18269 20147 18303 20175
rect 18331 20147 23619 20175
rect 23647 20147 23681 20175
rect 23709 20147 33477 20175
rect 33505 20147 33539 20175
rect 33567 20147 33601 20175
rect 33629 20147 33663 20175
rect 33691 20147 38979 20175
rect 39007 20147 39041 20175
rect 39069 20147 48837 20175
rect 48865 20147 48899 20175
rect 48927 20147 48961 20175
rect 48989 20147 49023 20175
rect 49051 20147 54339 20175
rect 54367 20147 54401 20175
rect 54429 20147 64197 20175
rect 64225 20147 64259 20175
rect 64287 20147 64321 20175
rect 64349 20147 64383 20175
rect 64411 20147 69699 20175
rect 69727 20147 69761 20175
rect 69789 20147 79557 20175
rect 79585 20147 79619 20175
rect 79647 20147 79681 20175
rect 79709 20147 79743 20175
rect 79771 20147 85059 20175
rect 85087 20147 85121 20175
rect 85149 20147 94917 20175
rect 94945 20147 94979 20175
rect 95007 20147 95041 20175
rect 95069 20147 95103 20175
rect 95131 20147 100419 20175
rect 100447 20147 100481 20175
rect 100509 20147 110277 20175
rect 110305 20147 110339 20175
rect 110367 20147 110401 20175
rect 110429 20147 110463 20175
rect 110491 20147 115779 20175
rect 115807 20147 115841 20175
rect 115869 20147 125637 20175
rect 125665 20147 125699 20175
rect 125727 20147 125761 20175
rect 125789 20147 125823 20175
rect 125851 20147 131139 20175
rect 131167 20147 131201 20175
rect 131229 20147 140997 20175
rect 141025 20147 141059 20175
rect 141087 20147 141121 20175
rect 141149 20147 141183 20175
rect 141211 20147 146499 20175
rect 146527 20147 146561 20175
rect 146589 20147 156357 20175
rect 156385 20147 156419 20175
rect 156447 20147 156481 20175
rect 156509 20147 156543 20175
rect 156571 20147 161859 20175
rect 161887 20147 161921 20175
rect 161949 20147 171717 20175
rect 171745 20147 171779 20175
rect 171807 20147 171841 20175
rect 171869 20147 171903 20175
rect 171931 20147 177219 20175
rect 177247 20147 177281 20175
rect 177309 20147 187077 20175
rect 187105 20147 187139 20175
rect 187167 20147 187201 20175
rect 187229 20147 187263 20175
rect 187291 20147 192579 20175
rect 192607 20147 192641 20175
rect 192669 20147 202437 20175
rect 202465 20147 202499 20175
rect 202527 20147 202561 20175
rect 202589 20147 202623 20175
rect 202651 20147 207939 20175
rect 207967 20147 208001 20175
rect 208029 20147 217797 20175
rect 217825 20147 217859 20175
rect 217887 20147 217921 20175
rect 217949 20147 217983 20175
rect 218011 20147 223299 20175
rect 223327 20147 223361 20175
rect 223389 20147 233157 20175
rect 233185 20147 233219 20175
rect 233247 20147 233281 20175
rect 233309 20147 233343 20175
rect 233371 20147 238659 20175
rect 238687 20147 238721 20175
rect 238749 20147 248517 20175
rect 248545 20147 248579 20175
rect 248607 20147 248641 20175
rect 248669 20147 248703 20175
rect 248731 20147 254019 20175
rect 254047 20147 254081 20175
rect 254109 20147 263877 20175
rect 263905 20147 263939 20175
rect 263967 20147 264001 20175
rect 264029 20147 264063 20175
rect 264091 20147 269379 20175
rect 269407 20147 269441 20175
rect 269469 20147 279237 20175
rect 279265 20147 279299 20175
rect 279327 20147 279361 20175
rect 279389 20147 279423 20175
rect 279451 20147 284739 20175
rect 284767 20147 284801 20175
rect 284829 20147 294597 20175
rect 294625 20147 294659 20175
rect 294687 20147 294721 20175
rect 294749 20147 294783 20175
rect 294811 20147 298248 20175
rect 298276 20147 298310 20175
rect 298338 20147 298372 20175
rect 298400 20147 298434 20175
rect 298462 20147 298990 20175
rect -958 20113 298990 20147
rect -958 20085 -430 20113
rect -402 20085 -368 20113
rect -340 20085 -306 20113
rect -278 20085 -244 20113
rect -216 20085 2757 20113
rect 2785 20085 2819 20113
rect 2847 20085 2881 20113
rect 2909 20085 2943 20113
rect 2971 20085 8259 20113
rect 8287 20085 8321 20113
rect 8349 20085 18117 20113
rect 18145 20085 18179 20113
rect 18207 20085 18241 20113
rect 18269 20085 18303 20113
rect 18331 20085 23619 20113
rect 23647 20085 23681 20113
rect 23709 20085 33477 20113
rect 33505 20085 33539 20113
rect 33567 20085 33601 20113
rect 33629 20085 33663 20113
rect 33691 20085 38979 20113
rect 39007 20085 39041 20113
rect 39069 20085 48837 20113
rect 48865 20085 48899 20113
rect 48927 20085 48961 20113
rect 48989 20085 49023 20113
rect 49051 20085 54339 20113
rect 54367 20085 54401 20113
rect 54429 20085 64197 20113
rect 64225 20085 64259 20113
rect 64287 20085 64321 20113
rect 64349 20085 64383 20113
rect 64411 20085 69699 20113
rect 69727 20085 69761 20113
rect 69789 20085 79557 20113
rect 79585 20085 79619 20113
rect 79647 20085 79681 20113
rect 79709 20085 79743 20113
rect 79771 20085 85059 20113
rect 85087 20085 85121 20113
rect 85149 20085 94917 20113
rect 94945 20085 94979 20113
rect 95007 20085 95041 20113
rect 95069 20085 95103 20113
rect 95131 20085 100419 20113
rect 100447 20085 100481 20113
rect 100509 20085 110277 20113
rect 110305 20085 110339 20113
rect 110367 20085 110401 20113
rect 110429 20085 110463 20113
rect 110491 20085 115779 20113
rect 115807 20085 115841 20113
rect 115869 20085 125637 20113
rect 125665 20085 125699 20113
rect 125727 20085 125761 20113
rect 125789 20085 125823 20113
rect 125851 20085 131139 20113
rect 131167 20085 131201 20113
rect 131229 20085 140997 20113
rect 141025 20085 141059 20113
rect 141087 20085 141121 20113
rect 141149 20085 141183 20113
rect 141211 20085 146499 20113
rect 146527 20085 146561 20113
rect 146589 20085 156357 20113
rect 156385 20085 156419 20113
rect 156447 20085 156481 20113
rect 156509 20085 156543 20113
rect 156571 20085 161859 20113
rect 161887 20085 161921 20113
rect 161949 20085 171717 20113
rect 171745 20085 171779 20113
rect 171807 20085 171841 20113
rect 171869 20085 171903 20113
rect 171931 20085 177219 20113
rect 177247 20085 177281 20113
rect 177309 20085 187077 20113
rect 187105 20085 187139 20113
rect 187167 20085 187201 20113
rect 187229 20085 187263 20113
rect 187291 20085 192579 20113
rect 192607 20085 192641 20113
rect 192669 20085 202437 20113
rect 202465 20085 202499 20113
rect 202527 20085 202561 20113
rect 202589 20085 202623 20113
rect 202651 20085 207939 20113
rect 207967 20085 208001 20113
rect 208029 20085 217797 20113
rect 217825 20085 217859 20113
rect 217887 20085 217921 20113
rect 217949 20085 217983 20113
rect 218011 20085 223299 20113
rect 223327 20085 223361 20113
rect 223389 20085 233157 20113
rect 233185 20085 233219 20113
rect 233247 20085 233281 20113
rect 233309 20085 233343 20113
rect 233371 20085 238659 20113
rect 238687 20085 238721 20113
rect 238749 20085 248517 20113
rect 248545 20085 248579 20113
rect 248607 20085 248641 20113
rect 248669 20085 248703 20113
rect 248731 20085 254019 20113
rect 254047 20085 254081 20113
rect 254109 20085 263877 20113
rect 263905 20085 263939 20113
rect 263967 20085 264001 20113
rect 264029 20085 264063 20113
rect 264091 20085 269379 20113
rect 269407 20085 269441 20113
rect 269469 20085 279237 20113
rect 279265 20085 279299 20113
rect 279327 20085 279361 20113
rect 279389 20085 279423 20113
rect 279451 20085 284739 20113
rect 284767 20085 284801 20113
rect 284829 20085 294597 20113
rect 294625 20085 294659 20113
rect 294687 20085 294721 20113
rect 294749 20085 294783 20113
rect 294811 20085 298248 20113
rect 298276 20085 298310 20113
rect 298338 20085 298372 20113
rect 298400 20085 298434 20113
rect 298462 20085 298990 20113
rect -958 20051 298990 20085
rect -958 20023 -430 20051
rect -402 20023 -368 20051
rect -340 20023 -306 20051
rect -278 20023 -244 20051
rect -216 20023 2757 20051
rect 2785 20023 2819 20051
rect 2847 20023 2881 20051
rect 2909 20023 2943 20051
rect 2971 20023 8259 20051
rect 8287 20023 8321 20051
rect 8349 20023 18117 20051
rect 18145 20023 18179 20051
rect 18207 20023 18241 20051
rect 18269 20023 18303 20051
rect 18331 20023 23619 20051
rect 23647 20023 23681 20051
rect 23709 20023 33477 20051
rect 33505 20023 33539 20051
rect 33567 20023 33601 20051
rect 33629 20023 33663 20051
rect 33691 20023 38979 20051
rect 39007 20023 39041 20051
rect 39069 20023 48837 20051
rect 48865 20023 48899 20051
rect 48927 20023 48961 20051
rect 48989 20023 49023 20051
rect 49051 20023 54339 20051
rect 54367 20023 54401 20051
rect 54429 20023 64197 20051
rect 64225 20023 64259 20051
rect 64287 20023 64321 20051
rect 64349 20023 64383 20051
rect 64411 20023 69699 20051
rect 69727 20023 69761 20051
rect 69789 20023 79557 20051
rect 79585 20023 79619 20051
rect 79647 20023 79681 20051
rect 79709 20023 79743 20051
rect 79771 20023 85059 20051
rect 85087 20023 85121 20051
rect 85149 20023 94917 20051
rect 94945 20023 94979 20051
rect 95007 20023 95041 20051
rect 95069 20023 95103 20051
rect 95131 20023 100419 20051
rect 100447 20023 100481 20051
rect 100509 20023 110277 20051
rect 110305 20023 110339 20051
rect 110367 20023 110401 20051
rect 110429 20023 110463 20051
rect 110491 20023 115779 20051
rect 115807 20023 115841 20051
rect 115869 20023 125637 20051
rect 125665 20023 125699 20051
rect 125727 20023 125761 20051
rect 125789 20023 125823 20051
rect 125851 20023 131139 20051
rect 131167 20023 131201 20051
rect 131229 20023 140997 20051
rect 141025 20023 141059 20051
rect 141087 20023 141121 20051
rect 141149 20023 141183 20051
rect 141211 20023 146499 20051
rect 146527 20023 146561 20051
rect 146589 20023 156357 20051
rect 156385 20023 156419 20051
rect 156447 20023 156481 20051
rect 156509 20023 156543 20051
rect 156571 20023 161859 20051
rect 161887 20023 161921 20051
rect 161949 20023 171717 20051
rect 171745 20023 171779 20051
rect 171807 20023 171841 20051
rect 171869 20023 171903 20051
rect 171931 20023 177219 20051
rect 177247 20023 177281 20051
rect 177309 20023 187077 20051
rect 187105 20023 187139 20051
rect 187167 20023 187201 20051
rect 187229 20023 187263 20051
rect 187291 20023 192579 20051
rect 192607 20023 192641 20051
rect 192669 20023 202437 20051
rect 202465 20023 202499 20051
rect 202527 20023 202561 20051
rect 202589 20023 202623 20051
rect 202651 20023 207939 20051
rect 207967 20023 208001 20051
rect 208029 20023 217797 20051
rect 217825 20023 217859 20051
rect 217887 20023 217921 20051
rect 217949 20023 217983 20051
rect 218011 20023 223299 20051
rect 223327 20023 223361 20051
rect 223389 20023 233157 20051
rect 233185 20023 233219 20051
rect 233247 20023 233281 20051
rect 233309 20023 233343 20051
rect 233371 20023 238659 20051
rect 238687 20023 238721 20051
rect 238749 20023 248517 20051
rect 248545 20023 248579 20051
rect 248607 20023 248641 20051
rect 248669 20023 248703 20051
rect 248731 20023 254019 20051
rect 254047 20023 254081 20051
rect 254109 20023 263877 20051
rect 263905 20023 263939 20051
rect 263967 20023 264001 20051
rect 264029 20023 264063 20051
rect 264091 20023 269379 20051
rect 269407 20023 269441 20051
rect 269469 20023 279237 20051
rect 279265 20023 279299 20051
rect 279327 20023 279361 20051
rect 279389 20023 279423 20051
rect 279451 20023 284739 20051
rect 284767 20023 284801 20051
rect 284829 20023 294597 20051
rect 294625 20023 294659 20051
rect 294687 20023 294721 20051
rect 294749 20023 294783 20051
rect 294811 20023 298248 20051
rect 298276 20023 298310 20051
rect 298338 20023 298372 20051
rect 298400 20023 298434 20051
rect 298462 20023 298990 20051
rect -958 19989 298990 20023
rect -958 19961 -430 19989
rect -402 19961 -368 19989
rect -340 19961 -306 19989
rect -278 19961 -244 19989
rect -216 19961 2757 19989
rect 2785 19961 2819 19989
rect 2847 19961 2881 19989
rect 2909 19961 2943 19989
rect 2971 19961 8259 19989
rect 8287 19961 8321 19989
rect 8349 19961 18117 19989
rect 18145 19961 18179 19989
rect 18207 19961 18241 19989
rect 18269 19961 18303 19989
rect 18331 19961 23619 19989
rect 23647 19961 23681 19989
rect 23709 19961 33477 19989
rect 33505 19961 33539 19989
rect 33567 19961 33601 19989
rect 33629 19961 33663 19989
rect 33691 19961 38979 19989
rect 39007 19961 39041 19989
rect 39069 19961 48837 19989
rect 48865 19961 48899 19989
rect 48927 19961 48961 19989
rect 48989 19961 49023 19989
rect 49051 19961 54339 19989
rect 54367 19961 54401 19989
rect 54429 19961 64197 19989
rect 64225 19961 64259 19989
rect 64287 19961 64321 19989
rect 64349 19961 64383 19989
rect 64411 19961 69699 19989
rect 69727 19961 69761 19989
rect 69789 19961 79557 19989
rect 79585 19961 79619 19989
rect 79647 19961 79681 19989
rect 79709 19961 79743 19989
rect 79771 19961 85059 19989
rect 85087 19961 85121 19989
rect 85149 19961 94917 19989
rect 94945 19961 94979 19989
rect 95007 19961 95041 19989
rect 95069 19961 95103 19989
rect 95131 19961 100419 19989
rect 100447 19961 100481 19989
rect 100509 19961 110277 19989
rect 110305 19961 110339 19989
rect 110367 19961 110401 19989
rect 110429 19961 110463 19989
rect 110491 19961 115779 19989
rect 115807 19961 115841 19989
rect 115869 19961 125637 19989
rect 125665 19961 125699 19989
rect 125727 19961 125761 19989
rect 125789 19961 125823 19989
rect 125851 19961 131139 19989
rect 131167 19961 131201 19989
rect 131229 19961 140997 19989
rect 141025 19961 141059 19989
rect 141087 19961 141121 19989
rect 141149 19961 141183 19989
rect 141211 19961 146499 19989
rect 146527 19961 146561 19989
rect 146589 19961 156357 19989
rect 156385 19961 156419 19989
rect 156447 19961 156481 19989
rect 156509 19961 156543 19989
rect 156571 19961 161859 19989
rect 161887 19961 161921 19989
rect 161949 19961 171717 19989
rect 171745 19961 171779 19989
rect 171807 19961 171841 19989
rect 171869 19961 171903 19989
rect 171931 19961 177219 19989
rect 177247 19961 177281 19989
rect 177309 19961 187077 19989
rect 187105 19961 187139 19989
rect 187167 19961 187201 19989
rect 187229 19961 187263 19989
rect 187291 19961 192579 19989
rect 192607 19961 192641 19989
rect 192669 19961 202437 19989
rect 202465 19961 202499 19989
rect 202527 19961 202561 19989
rect 202589 19961 202623 19989
rect 202651 19961 207939 19989
rect 207967 19961 208001 19989
rect 208029 19961 217797 19989
rect 217825 19961 217859 19989
rect 217887 19961 217921 19989
rect 217949 19961 217983 19989
rect 218011 19961 223299 19989
rect 223327 19961 223361 19989
rect 223389 19961 233157 19989
rect 233185 19961 233219 19989
rect 233247 19961 233281 19989
rect 233309 19961 233343 19989
rect 233371 19961 238659 19989
rect 238687 19961 238721 19989
rect 238749 19961 248517 19989
rect 248545 19961 248579 19989
rect 248607 19961 248641 19989
rect 248669 19961 248703 19989
rect 248731 19961 254019 19989
rect 254047 19961 254081 19989
rect 254109 19961 263877 19989
rect 263905 19961 263939 19989
rect 263967 19961 264001 19989
rect 264029 19961 264063 19989
rect 264091 19961 269379 19989
rect 269407 19961 269441 19989
rect 269469 19961 279237 19989
rect 279265 19961 279299 19989
rect 279327 19961 279361 19989
rect 279389 19961 279423 19989
rect 279451 19961 284739 19989
rect 284767 19961 284801 19989
rect 284829 19961 294597 19989
rect 294625 19961 294659 19989
rect 294687 19961 294721 19989
rect 294749 19961 294783 19989
rect 294811 19961 298248 19989
rect 298276 19961 298310 19989
rect 298338 19961 298372 19989
rect 298400 19961 298434 19989
rect 298462 19961 298990 19989
rect -958 19913 298990 19961
rect -958 14175 298990 14223
rect -958 14147 -910 14175
rect -882 14147 -848 14175
rect -820 14147 -786 14175
rect -758 14147 -724 14175
rect -696 14147 4617 14175
rect 4645 14147 4679 14175
rect 4707 14147 4741 14175
rect 4769 14147 4803 14175
rect 4831 14147 15939 14175
rect 15967 14147 16001 14175
rect 16029 14147 19977 14175
rect 20005 14147 20039 14175
rect 20067 14147 20101 14175
rect 20129 14147 20163 14175
rect 20191 14147 31299 14175
rect 31327 14147 31361 14175
rect 31389 14147 35337 14175
rect 35365 14147 35399 14175
rect 35427 14147 35461 14175
rect 35489 14147 35523 14175
rect 35551 14147 46659 14175
rect 46687 14147 46721 14175
rect 46749 14147 50697 14175
rect 50725 14147 50759 14175
rect 50787 14147 50821 14175
rect 50849 14147 50883 14175
rect 50911 14147 62019 14175
rect 62047 14147 62081 14175
rect 62109 14147 66057 14175
rect 66085 14147 66119 14175
rect 66147 14147 66181 14175
rect 66209 14147 66243 14175
rect 66271 14147 77379 14175
rect 77407 14147 77441 14175
rect 77469 14147 81417 14175
rect 81445 14147 81479 14175
rect 81507 14147 81541 14175
rect 81569 14147 81603 14175
rect 81631 14147 92739 14175
rect 92767 14147 92801 14175
rect 92829 14147 96777 14175
rect 96805 14147 96839 14175
rect 96867 14147 96901 14175
rect 96929 14147 96963 14175
rect 96991 14147 108099 14175
rect 108127 14147 108161 14175
rect 108189 14147 112137 14175
rect 112165 14147 112199 14175
rect 112227 14147 112261 14175
rect 112289 14147 112323 14175
rect 112351 14147 123459 14175
rect 123487 14147 123521 14175
rect 123549 14147 127497 14175
rect 127525 14147 127559 14175
rect 127587 14147 127621 14175
rect 127649 14147 127683 14175
rect 127711 14147 138819 14175
rect 138847 14147 138881 14175
rect 138909 14147 142857 14175
rect 142885 14147 142919 14175
rect 142947 14147 142981 14175
rect 143009 14147 143043 14175
rect 143071 14147 154179 14175
rect 154207 14147 154241 14175
rect 154269 14147 158217 14175
rect 158245 14147 158279 14175
rect 158307 14147 158341 14175
rect 158369 14147 158403 14175
rect 158431 14147 169539 14175
rect 169567 14147 169601 14175
rect 169629 14147 173577 14175
rect 173605 14147 173639 14175
rect 173667 14147 173701 14175
rect 173729 14147 173763 14175
rect 173791 14147 184899 14175
rect 184927 14147 184961 14175
rect 184989 14147 188937 14175
rect 188965 14147 188999 14175
rect 189027 14147 189061 14175
rect 189089 14147 189123 14175
rect 189151 14147 200259 14175
rect 200287 14147 200321 14175
rect 200349 14147 204297 14175
rect 204325 14147 204359 14175
rect 204387 14147 204421 14175
rect 204449 14147 204483 14175
rect 204511 14147 215619 14175
rect 215647 14147 215681 14175
rect 215709 14147 219657 14175
rect 219685 14147 219719 14175
rect 219747 14147 219781 14175
rect 219809 14147 219843 14175
rect 219871 14147 230979 14175
rect 231007 14147 231041 14175
rect 231069 14147 235017 14175
rect 235045 14147 235079 14175
rect 235107 14147 235141 14175
rect 235169 14147 235203 14175
rect 235231 14147 246339 14175
rect 246367 14147 246401 14175
rect 246429 14147 250377 14175
rect 250405 14147 250439 14175
rect 250467 14147 250501 14175
rect 250529 14147 250563 14175
rect 250591 14147 261699 14175
rect 261727 14147 261761 14175
rect 261789 14147 265737 14175
rect 265765 14147 265799 14175
rect 265827 14147 265861 14175
rect 265889 14147 265923 14175
rect 265951 14147 277059 14175
rect 277087 14147 277121 14175
rect 277149 14147 281097 14175
rect 281125 14147 281159 14175
rect 281187 14147 281221 14175
rect 281249 14147 281283 14175
rect 281311 14147 296457 14175
rect 296485 14147 296519 14175
rect 296547 14147 296581 14175
rect 296609 14147 296643 14175
rect 296671 14147 298728 14175
rect 298756 14147 298790 14175
rect 298818 14147 298852 14175
rect 298880 14147 298914 14175
rect 298942 14147 298990 14175
rect -958 14113 298990 14147
rect -958 14085 -910 14113
rect -882 14085 -848 14113
rect -820 14085 -786 14113
rect -758 14085 -724 14113
rect -696 14085 4617 14113
rect 4645 14085 4679 14113
rect 4707 14085 4741 14113
rect 4769 14085 4803 14113
rect 4831 14085 15939 14113
rect 15967 14085 16001 14113
rect 16029 14085 19977 14113
rect 20005 14085 20039 14113
rect 20067 14085 20101 14113
rect 20129 14085 20163 14113
rect 20191 14085 31299 14113
rect 31327 14085 31361 14113
rect 31389 14085 35337 14113
rect 35365 14085 35399 14113
rect 35427 14085 35461 14113
rect 35489 14085 35523 14113
rect 35551 14085 46659 14113
rect 46687 14085 46721 14113
rect 46749 14085 50697 14113
rect 50725 14085 50759 14113
rect 50787 14085 50821 14113
rect 50849 14085 50883 14113
rect 50911 14085 62019 14113
rect 62047 14085 62081 14113
rect 62109 14085 66057 14113
rect 66085 14085 66119 14113
rect 66147 14085 66181 14113
rect 66209 14085 66243 14113
rect 66271 14085 77379 14113
rect 77407 14085 77441 14113
rect 77469 14085 81417 14113
rect 81445 14085 81479 14113
rect 81507 14085 81541 14113
rect 81569 14085 81603 14113
rect 81631 14085 92739 14113
rect 92767 14085 92801 14113
rect 92829 14085 96777 14113
rect 96805 14085 96839 14113
rect 96867 14085 96901 14113
rect 96929 14085 96963 14113
rect 96991 14085 108099 14113
rect 108127 14085 108161 14113
rect 108189 14085 112137 14113
rect 112165 14085 112199 14113
rect 112227 14085 112261 14113
rect 112289 14085 112323 14113
rect 112351 14085 123459 14113
rect 123487 14085 123521 14113
rect 123549 14085 127497 14113
rect 127525 14085 127559 14113
rect 127587 14085 127621 14113
rect 127649 14085 127683 14113
rect 127711 14085 138819 14113
rect 138847 14085 138881 14113
rect 138909 14085 142857 14113
rect 142885 14085 142919 14113
rect 142947 14085 142981 14113
rect 143009 14085 143043 14113
rect 143071 14085 154179 14113
rect 154207 14085 154241 14113
rect 154269 14085 158217 14113
rect 158245 14085 158279 14113
rect 158307 14085 158341 14113
rect 158369 14085 158403 14113
rect 158431 14085 169539 14113
rect 169567 14085 169601 14113
rect 169629 14085 173577 14113
rect 173605 14085 173639 14113
rect 173667 14085 173701 14113
rect 173729 14085 173763 14113
rect 173791 14085 184899 14113
rect 184927 14085 184961 14113
rect 184989 14085 188937 14113
rect 188965 14085 188999 14113
rect 189027 14085 189061 14113
rect 189089 14085 189123 14113
rect 189151 14085 200259 14113
rect 200287 14085 200321 14113
rect 200349 14085 204297 14113
rect 204325 14085 204359 14113
rect 204387 14085 204421 14113
rect 204449 14085 204483 14113
rect 204511 14085 215619 14113
rect 215647 14085 215681 14113
rect 215709 14085 219657 14113
rect 219685 14085 219719 14113
rect 219747 14085 219781 14113
rect 219809 14085 219843 14113
rect 219871 14085 230979 14113
rect 231007 14085 231041 14113
rect 231069 14085 235017 14113
rect 235045 14085 235079 14113
rect 235107 14085 235141 14113
rect 235169 14085 235203 14113
rect 235231 14085 246339 14113
rect 246367 14085 246401 14113
rect 246429 14085 250377 14113
rect 250405 14085 250439 14113
rect 250467 14085 250501 14113
rect 250529 14085 250563 14113
rect 250591 14085 261699 14113
rect 261727 14085 261761 14113
rect 261789 14085 265737 14113
rect 265765 14085 265799 14113
rect 265827 14085 265861 14113
rect 265889 14085 265923 14113
rect 265951 14085 277059 14113
rect 277087 14085 277121 14113
rect 277149 14085 281097 14113
rect 281125 14085 281159 14113
rect 281187 14085 281221 14113
rect 281249 14085 281283 14113
rect 281311 14085 296457 14113
rect 296485 14085 296519 14113
rect 296547 14085 296581 14113
rect 296609 14085 296643 14113
rect 296671 14085 298728 14113
rect 298756 14085 298790 14113
rect 298818 14085 298852 14113
rect 298880 14085 298914 14113
rect 298942 14085 298990 14113
rect -958 14051 298990 14085
rect -958 14023 -910 14051
rect -882 14023 -848 14051
rect -820 14023 -786 14051
rect -758 14023 -724 14051
rect -696 14023 4617 14051
rect 4645 14023 4679 14051
rect 4707 14023 4741 14051
rect 4769 14023 4803 14051
rect 4831 14023 15939 14051
rect 15967 14023 16001 14051
rect 16029 14023 19977 14051
rect 20005 14023 20039 14051
rect 20067 14023 20101 14051
rect 20129 14023 20163 14051
rect 20191 14023 31299 14051
rect 31327 14023 31361 14051
rect 31389 14023 35337 14051
rect 35365 14023 35399 14051
rect 35427 14023 35461 14051
rect 35489 14023 35523 14051
rect 35551 14023 46659 14051
rect 46687 14023 46721 14051
rect 46749 14023 50697 14051
rect 50725 14023 50759 14051
rect 50787 14023 50821 14051
rect 50849 14023 50883 14051
rect 50911 14023 62019 14051
rect 62047 14023 62081 14051
rect 62109 14023 66057 14051
rect 66085 14023 66119 14051
rect 66147 14023 66181 14051
rect 66209 14023 66243 14051
rect 66271 14023 77379 14051
rect 77407 14023 77441 14051
rect 77469 14023 81417 14051
rect 81445 14023 81479 14051
rect 81507 14023 81541 14051
rect 81569 14023 81603 14051
rect 81631 14023 92739 14051
rect 92767 14023 92801 14051
rect 92829 14023 96777 14051
rect 96805 14023 96839 14051
rect 96867 14023 96901 14051
rect 96929 14023 96963 14051
rect 96991 14023 108099 14051
rect 108127 14023 108161 14051
rect 108189 14023 112137 14051
rect 112165 14023 112199 14051
rect 112227 14023 112261 14051
rect 112289 14023 112323 14051
rect 112351 14023 123459 14051
rect 123487 14023 123521 14051
rect 123549 14023 127497 14051
rect 127525 14023 127559 14051
rect 127587 14023 127621 14051
rect 127649 14023 127683 14051
rect 127711 14023 138819 14051
rect 138847 14023 138881 14051
rect 138909 14023 142857 14051
rect 142885 14023 142919 14051
rect 142947 14023 142981 14051
rect 143009 14023 143043 14051
rect 143071 14023 154179 14051
rect 154207 14023 154241 14051
rect 154269 14023 158217 14051
rect 158245 14023 158279 14051
rect 158307 14023 158341 14051
rect 158369 14023 158403 14051
rect 158431 14023 169539 14051
rect 169567 14023 169601 14051
rect 169629 14023 173577 14051
rect 173605 14023 173639 14051
rect 173667 14023 173701 14051
rect 173729 14023 173763 14051
rect 173791 14023 184899 14051
rect 184927 14023 184961 14051
rect 184989 14023 188937 14051
rect 188965 14023 188999 14051
rect 189027 14023 189061 14051
rect 189089 14023 189123 14051
rect 189151 14023 200259 14051
rect 200287 14023 200321 14051
rect 200349 14023 204297 14051
rect 204325 14023 204359 14051
rect 204387 14023 204421 14051
rect 204449 14023 204483 14051
rect 204511 14023 215619 14051
rect 215647 14023 215681 14051
rect 215709 14023 219657 14051
rect 219685 14023 219719 14051
rect 219747 14023 219781 14051
rect 219809 14023 219843 14051
rect 219871 14023 230979 14051
rect 231007 14023 231041 14051
rect 231069 14023 235017 14051
rect 235045 14023 235079 14051
rect 235107 14023 235141 14051
rect 235169 14023 235203 14051
rect 235231 14023 246339 14051
rect 246367 14023 246401 14051
rect 246429 14023 250377 14051
rect 250405 14023 250439 14051
rect 250467 14023 250501 14051
rect 250529 14023 250563 14051
rect 250591 14023 261699 14051
rect 261727 14023 261761 14051
rect 261789 14023 265737 14051
rect 265765 14023 265799 14051
rect 265827 14023 265861 14051
rect 265889 14023 265923 14051
rect 265951 14023 277059 14051
rect 277087 14023 277121 14051
rect 277149 14023 281097 14051
rect 281125 14023 281159 14051
rect 281187 14023 281221 14051
rect 281249 14023 281283 14051
rect 281311 14023 296457 14051
rect 296485 14023 296519 14051
rect 296547 14023 296581 14051
rect 296609 14023 296643 14051
rect 296671 14023 298728 14051
rect 298756 14023 298790 14051
rect 298818 14023 298852 14051
rect 298880 14023 298914 14051
rect 298942 14023 298990 14051
rect -958 13989 298990 14023
rect -958 13961 -910 13989
rect -882 13961 -848 13989
rect -820 13961 -786 13989
rect -758 13961 -724 13989
rect -696 13961 4617 13989
rect 4645 13961 4679 13989
rect 4707 13961 4741 13989
rect 4769 13961 4803 13989
rect 4831 13961 15939 13989
rect 15967 13961 16001 13989
rect 16029 13961 19977 13989
rect 20005 13961 20039 13989
rect 20067 13961 20101 13989
rect 20129 13961 20163 13989
rect 20191 13961 31299 13989
rect 31327 13961 31361 13989
rect 31389 13961 35337 13989
rect 35365 13961 35399 13989
rect 35427 13961 35461 13989
rect 35489 13961 35523 13989
rect 35551 13961 46659 13989
rect 46687 13961 46721 13989
rect 46749 13961 50697 13989
rect 50725 13961 50759 13989
rect 50787 13961 50821 13989
rect 50849 13961 50883 13989
rect 50911 13961 62019 13989
rect 62047 13961 62081 13989
rect 62109 13961 66057 13989
rect 66085 13961 66119 13989
rect 66147 13961 66181 13989
rect 66209 13961 66243 13989
rect 66271 13961 77379 13989
rect 77407 13961 77441 13989
rect 77469 13961 81417 13989
rect 81445 13961 81479 13989
rect 81507 13961 81541 13989
rect 81569 13961 81603 13989
rect 81631 13961 92739 13989
rect 92767 13961 92801 13989
rect 92829 13961 96777 13989
rect 96805 13961 96839 13989
rect 96867 13961 96901 13989
rect 96929 13961 96963 13989
rect 96991 13961 108099 13989
rect 108127 13961 108161 13989
rect 108189 13961 112137 13989
rect 112165 13961 112199 13989
rect 112227 13961 112261 13989
rect 112289 13961 112323 13989
rect 112351 13961 123459 13989
rect 123487 13961 123521 13989
rect 123549 13961 127497 13989
rect 127525 13961 127559 13989
rect 127587 13961 127621 13989
rect 127649 13961 127683 13989
rect 127711 13961 138819 13989
rect 138847 13961 138881 13989
rect 138909 13961 142857 13989
rect 142885 13961 142919 13989
rect 142947 13961 142981 13989
rect 143009 13961 143043 13989
rect 143071 13961 154179 13989
rect 154207 13961 154241 13989
rect 154269 13961 158217 13989
rect 158245 13961 158279 13989
rect 158307 13961 158341 13989
rect 158369 13961 158403 13989
rect 158431 13961 169539 13989
rect 169567 13961 169601 13989
rect 169629 13961 173577 13989
rect 173605 13961 173639 13989
rect 173667 13961 173701 13989
rect 173729 13961 173763 13989
rect 173791 13961 184899 13989
rect 184927 13961 184961 13989
rect 184989 13961 188937 13989
rect 188965 13961 188999 13989
rect 189027 13961 189061 13989
rect 189089 13961 189123 13989
rect 189151 13961 200259 13989
rect 200287 13961 200321 13989
rect 200349 13961 204297 13989
rect 204325 13961 204359 13989
rect 204387 13961 204421 13989
rect 204449 13961 204483 13989
rect 204511 13961 215619 13989
rect 215647 13961 215681 13989
rect 215709 13961 219657 13989
rect 219685 13961 219719 13989
rect 219747 13961 219781 13989
rect 219809 13961 219843 13989
rect 219871 13961 230979 13989
rect 231007 13961 231041 13989
rect 231069 13961 235017 13989
rect 235045 13961 235079 13989
rect 235107 13961 235141 13989
rect 235169 13961 235203 13989
rect 235231 13961 246339 13989
rect 246367 13961 246401 13989
rect 246429 13961 250377 13989
rect 250405 13961 250439 13989
rect 250467 13961 250501 13989
rect 250529 13961 250563 13989
rect 250591 13961 261699 13989
rect 261727 13961 261761 13989
rect 261789 13961 265737 13989
rect 265765 13961 265799 13989
rect 265827 13961 265861 13989
rect 265889 13961 265923 13989
rect 265951 13961 277059 13989
rect 277087 13961 277121 13989
rect 277149 13961 281097 13989
rect 281125 13961 281159 13989
rect 281187 13961 281221 13989
rect 281249 13961 281283 13989
rect 281311 13961 296457 13989
rect 296485 13961 296519 13989
rect 296547 13961 296581 13989
rect 296609 13961 296643 13989
rect 296671 13961 298728 13989
rect 298756 13961 298790 13989
rect 298818 13961 298852 13989
rect 298880 13961 298914 13989
rect 298942 13961 298990 13989
rect -958 13913 298990 13961
rect -958 11175 298990 11223
rect -958 11147 -430 11175
rect -402 11147 -368 11175
rect -340 11147 -306 11175
rect -278 11147 -244 11175
rect -216 11147 2757 11175
rect 2785 11147 2819 11175
rect 2847 11147 2881 11175
rect 2909 11147 2943 11175
rect 2971 11147 8259 11175
rect 8287 11147 8321 11175
rect 8349 11147 18117 11175
rect 18145 11147 18179 11175
rect 18207 11147 18241 11175
rect 18269 11147 18303 11175
rect 18331 11147 23619 11175
rect 23647 11147 23681 11175
rect 23709 11147 33477 11175
rect 33505 11147 33539 11175
rect 33567 11147 33601 11175
rect 33629 11147 33663 11175
rect 33691 11147 38979 11175
rect 39007 11147 39041 11175
rect 39069 11147 48837 11175
rect 48865 11147 48899 11175
rect 48927 11147 48961 11175
rect 48989 11147 49023 11175
rect 49051 11147 54339 11175
rect 54367 11147 54401 11175
rect 54429 11147 64197 11175
rect 64225 11147 64259 11175
rect 64287 11147 64321 11175
rect 64349 11147 64383 11175
rect 64411 11147 69699 11175
rect 69727 11147 69761 11175
rect 69789 11147 79557 11175
rect 79585 11147 79619 11175
rect 79647 11147 79681 11175
rect 79709 11147 79743 11175
rect 79771 11147 85059 11175
rect 85087 11147 85121 11175
rect 85149 11147 94917 11175
rect 94945 11147 94979 11175
rect 95007 11147 95041 11175
rect 95069 11147 95103 11175
rect 95131 11147 100419 11175
rect 100447 11147 100481 11175
rect 100509 11147 110277 11175
rect 110305 11147 110339 11175
rect 110367 11147 110401 11175
rect 110429 11147 110463 11175
rect 110491 11147 115779 11175
rect 115807 11147 115841 11175
rect 115869 11147 125637 11175
rect 125665 11147 125699 11175
rect 125727 11147 125761 11175
rect 125789 11147 125823 11175
rect 125851 11147 131139 11175
rect 131167 11147 131201 11175
rect 131229 11147 140997 11175
rect 141025 11147 141059 11175
rect 141087 11147 141121 11175
rect 141149 11147 141183 11175
rect 141211 11147 146499 11175
rect 146527 11147 146561 11175
rect 146589 11147 156357 11175
rect 156385 11147 156419 11175
rect 156447 11147 156481 11175
rect 156509 11147 156543 11175
rect 156571 11147 161859 11175
rect 161887 11147 161921 11175
rect 161949 11147 171717 11175
rect 171745 11147 171779 11175
rect 171807 11147 171841 11175
rect 171869 11147 171903 11175
rect 171931 11147 177219 11175
rect 177247 11147 177281 11175
rect 177309 11147 187077 11175
rect 187105 11147 187139 11175
rect 187167 11147 187201 11175
rect 187229 11147 187263 11175
rect 187291 11147 192579 11175
rect 192607 11147 192641 11175
rect 192669 11147 202437 11175
rect 202465 11147 202499 11175
rect 202527 11147 202561 11175
rect 202589 11147 202623 11175
rect 202651 11147 207939 11175
rect 207967 11147 208001 11175
rect 208029 11147 217797 11175
rect 217825 11147 217859 11175
rect 217887 11147 217921 11175
rect 217949 11147 217983 11175
rect 218011 11147 223299 11175
rect 223327 11147 223361 11175
rect 223389 11147 233157 11175
rect 233185 11147 233219 11175
rect 233247 11147 233281 11175
rect 233309 11147 233343 11175
rect 233371 11147 238659 11175
rect 238687 11147 238721 11175
rect 238749 11147 248517 11175
rect 248545 11147 248579 11175
rect 248607 11147 248641 11175
rect 248669 11147 248703 11175
rect 248731 11147 254019 11175
rect 254047 11147 254081 11175
rect 254109 11147 263877 11175
rect 263905 11147 263939 11175
rect 263967 11147 264001 11175
rect 264029 11147 264063 11175
rect 264091 11147 269379 11175
rect 269407 11147 269441 11175
rect 269469 11147 279237 11175
rect 279265 11147 279299 11175
rect 279327 11147 279361 11175
rect 279389 11147 279423 11175
rect 279451 11147 284739 11175
rect 284767 11147 284801 11175
rect 284829 11147 294597 11175
rect 294625 11147 294659 11175
rect 294687 11147 294721 11175
rect 294749 11147 294783 11175
rect 294811 11147 298248 11175
rect 298276 11147 298310 11175
rect 298338 11147 298372 11175
rect 298400 11147 298434 11175
rect 298462 11147 298990 11175
rect -958 11113 298990 11147
rect -958 11085 -430 11113
rect -402 11085 -368 11113
rect -340 11085 -306 11113
rect -278 11085 -244 11113
rect -216 11085 2757 11113
rect 2785 11085 2819 11113
rect 2847 11085 2881 11113
rect 2909 11085 2943 11113
rect 2971 11085 8259 11113
rect 8287 11085 8321 11113
rect 8349 11085 18117 11113
rect 18145 11085 18179 11113
rect 18207 11085 18241 11113
rect 18269 11085 18303 11113
rect 18331 11085 23619 11113
rect 23647 11085 23681 11113
rect 23709 11085 33477 11113
rect 33505 11085 33539 11113
rect 33567 11085 33601 11113
rect 33629 11085 33663 11113
rect 33691 11085 38979 11113
rect 39007 11085 39041 11113
rect 39069 11085 48837 11113
rect 48865 11085 48899 11113
rect 48927 11085 48961 11113
rect 48989 11085 49023 11113
rect 49051 11085 54339 11113
rect 54367 11085 54401 11113
rect 54429 11085 64197 11113
rect 64225 11085 64259 11113
rect 64287 11085 64321 11113
rect 64349 11085 64383 11113
rect 64411 11085 69699 11113
rect 69727 11085 69761 11113
rect 69789 11085 79557 11113
rect 79585 11085 79619 11113
rect 79647 11085 79681 11113
rect 79709 11085 79743 11113
rect 79771 11085 85059 11113
rect 85087 11085 85121 11113
rect 85149 11085 94917 11113
rect 94945 11085 94979 11113
rect 95007 11085 95041 11113
rect 95069 11085 95103 11113
rect 95131 11085 100419 11113
rect 100447 11085 100481 11113
rect 100509 11085 110277 11113
rect 110305 11085 110339 11113
rect 110367 11085 110401 11113
rect 110429 11085 110463 11113
rect 110491 11085 115779 11113
rect 115807 11085 115841 11113
rect 115869 11085 125637 11113
rect 125665 11085 125699 11113
rect 125727 11085 125761 11113
rect 125789 11085 125823 11113
rect 125851 11085 131139 11113
rect 131167 11085 131201 11113
rect 131229 11085 140997 11113
rect 141025 11085 141059 11113
rect 141087 11085 141121 11113
rect 141149 11085 141183 11113
rect 141211 11085 146499 11113
rect 146527 11085 146561 11113
rect 146589 11085 156357 11113
rect 156385 11085 156419 11113
rect 156447 11085 156481 11113
rect 156509 11085 156543 11113
rect 156571 11085 161859 11113
rect 161887 11085 161921 11113
rect 161949 11085 171717 11113
rect 171745 11085 171779 11113
rect 171807 11085 171841 11113
rect 171869 11085 171903 11113
rect 171931 11085 177219 11113
rect 177247 11085 177281 11113
rect 177309 11085 187077 11113
rect 187105 11085 187139 11113
rect 187167 11085 187201 11113
rect 187229 11085 187263 11113
rect 187291 11085 192579 11113
rect 192607 11085 192641 11113
rect 192669 11085 202437 11113
rect 202465 11085 202499 11113
rect 202527 11085 202561 11113
rect 202589 11085 202623 11113
rect 202651 11085 207939 11113
rect 207967 11085 208001 11113
rect 208029 11085 217797 11113
rect 217825 11085 217859 11113
rect 217887 11085 217921 11113
rect 217949 11085 217983 11113
rect 218011 11085 223299 11113
rect 223327 11085 223361 11113
rect 223389 11085 233157 11113
rect 233185 11085 233219 11113
rect 233247 11085 233281 11113
rect 233309 11085 233343 11113
rect 233371 11085 238659 11113
rect 238687 11085 238721 11113
rect 238749 11085 248517 11113
rect 248545 11085 248579 11113
rect 248607 11085 248641 11113
rect 248669 11085 248703 11113
rect 248731 11085 254019 11113
rect 254047 11085 254081 11113
rect 254109 11085 263877 11113
rect 263905 11085 263939 11113
rect 263967 11085 264001 11113
rect 264029 11085 264063 11113
rect 264091 11085 269379 11113
rect 269407 11085 269441 11113
rect 269469 11085 279237 11113
rect 279265 11085 279299 11113
rect 279327 11085 279361 11113
rect 279389 11085 279423 11113
rect 279451 11085 284739 11113
rect 284767 11085 284801 11113
rect 284829 11085 294597 11113
rect 294625 11085 294659 11113
rect 294687 11085 294721 11113
rect 294749 11085 294783 11113
rect 294811 11085 298248 11113
rect 298276 11085 298310 11113
rect 298338 11085 298372 11113
rect 298400 11085 298434 11113
rect 298462 11085 298990 11113
rect -958 11051 298990 11085
rect -958 11023 -430 11051
rect -402 11023 -368 11051
rect -340 11023 -306 11051
rect -278 11023 -244 11051
rect -216 11023 2757 11051
rect 2785 11023 2819 11051
rect 2847 11023 2881 11051
rect 2909 11023 2943 11051
rect 2971 11023 8259 11051
rect 8287 11023 8321 11051
rect 8349 11023 18117 11051
rect 18145 11023 18179 11051
rect 18207 11023 18241 11051
rect 18269 11023 18303 11051
rect 18331 11023 23619 11051
rect 23647 11023 23681 11051
rect 23709 11023 33477 11051
rect 33505 11023 33539 11051
rect 33567 11023 33601 11051
rect 33629 11023 33663 11051
rect 33691 11023 38979 11051
rect 39007 11023 39041 11051
rect 39069 11023 48837 11051
rect 48865 11023 48899 11051
rect 48927 11023 48961 11051
rect 48989 11023 49023 11051
rect 49051 11023 54339 11051
rect 54367 11023 54401 11051
rect 54429 11023 64197 11051
rect 64225 11023 64259 11051
rect 64287 11023 64321 11051
rect 64349 11023 64383 11051
rect 64411 11023 69699 11051
rect 69727 11023 69761 11051
rect 69789 11023 79557 11051
rect 79585 11023 79619 11051
rect 79647 11023 79681 11051
rect 79709 11023 79743 11051
rect 79771 11023 85059 11051
rect 85087 11023 85121 11051
rect 85149 11023 94917 11051
rect 94945 11023 94979 11051
rect 95007 11023 95041 11051
rect 95069 11023 95103 11051
rect 95131 11023 100419 11051
rect 100447 11023 100481 11051
rect 100509 11023 110277 11051
rect 110305 11023 110339 11051
rect 110367 11023 110401 11051
rect 110429 11023 110463 11051
rect 110491 11023 115779 11051
rect 115807 11023 115841 11051
rect 115869 11023 125637 11051
rect 125665 11023 125699 11051
rect 125727 11023 125761 11051
rect 125789 11023 125823 11051
rect 125851 11023 131139 11051
rect 131167 11023 131201 11051
rect 131229 11023 140997 11051
rect 141025 11023 141059 11051
rect 141087 11023 141121 11051
rect 141149 11023 141183 11051
rect 141211 11023 146499 11051
rect 146527 11023 146561 11051
rect 146589 11023 156357 11051
rect 156385 11023 156419 11051
rect 156447 11023 156481 11051
rect 156509 11023 156543 11051
rect 156571 11023 161859 11051
rect 161887 11023 161921 11051
rect 161949 11023 171717 11051
rect 171745 11023 171779 11051
rect 171807 11023 171841 11051
rect 171869 11023 171903 11051
rect 171931 11023 177219 11051
rect 177247 11023 177281 11051
rect 177309 11023 187077 11051
rect 187105 11023 187139 11051
rect 187167 11023 187201 11051
rect 187229 11023 187263 11051
rect 187291 11023 192579 11051
rect 192607 11023 192641 11051
rect 192669 11023 202437 11051
rect 202465 11023 202499 11051
rect 202527 11023 202561 11051
rect 202589 11023 202623 11051
rect 202651 11023 207939 11051
rect 207967 11023 208001 11051
rect 208029 11023 217797 11051
rect 217825 11023 217859 11051
rect 217887 11023 217921 11051
rect 217949 11023 217983 11051
rect 218011 11023 223299 11051
rect 223327 11023 223361 11051
rect 223389 11023 233157 11051
rect 233185 11023 233219 11051
rect 233247 11023 233281 11051
rect 233309 11023 233343 11051
rect 233371 11023 238659 11051
rect 238687 11023 238721 11051
rect 238749 11023 248517 11051
rect 248545 11023 248579 11051
rect 248607 11023 248641 11051
rect 248669 11023 248703 11051
rect 248731 11023 254019 11051
rect 254047 11023 254081 11051
rect 254109 11023 263877 11051
rect 263905 11023 263939 11051
rect 263967 11023 264001 11051
rect 264029 11023 264063 11051
rect 264091 11023 269379 11051
rect 269407 11023 269441 11051
rect 269469 11023 279237 11051
rect 279265 11023 279299 11051
rect 279327 11023 279361 11051
rect 279389 11023 279423 11051
rect 279451 11023 284739 11051
rect 284767 11023 284801 11051
rect 284829 11023 294597 11051
rect 294625 11023 294659 11051
rect 294687 11023 294721 11051
rect 294749 11023 294783 11051
rect 294811 11023 298248 11051
rect 298276 11023 298310 11051
rect 298338 11023 298372 11051
rect 298400 11023 298434 11051
rect 298462 11023 298990 11051
rect -958 10989 298990 11023
rect -958 10961 -430 10989
rect -402 10961 -368 10989
rect -340 10961 -306 10989
rect -278 10961 -244 10989
rect -216 10961 2757 10989
rect 2785 10961 2819 10989
rect 2847 10961 2881 10989
rect 2909 10961 2943 10989
rect 2971 10961 8259 10989
rect 8287 10961 8321 10989
rect 8349 10961 18117 10989
rect 18145 10961 18179 10989
rect 18207 10961 18241 10989
rect 18269 10961 18303 10989
rect 18331 10961 23619 10989
rect 23647 10961 23681 10989
rect 23709 10961 33477 10989
rect 33505 10961 33539 10989
rect 33567 10961 33601 10989
rect 33629 10961 33663 10989
rect 33691 10961 38979 10989
rect 39007 10961 39041 10989
rect 39069 10961 48837 10989
rect 48865 10961 48899 10989
rect 48927 10961 48961 10989
rect 48989 10961 49023 10989
rect 49051 10961 54339 10989
rect 54367 10961 54401 10989
rect 54429 10961 64197 10989
rect 64225 10961 64259 10989
rect 64287 10961 64321 10989
rect 64349 10961 64383 10989
rect 64411 10961 69699 10989
rect 69727 10961 69761 10989
rect 69789 10961 79557 10989
rect 79585 10961 79619 10989
rect 79647 10961 79681 10989
rect 79709 10961 79743 10989
rect 79771 10961 85059 10989
rect 85087 10961 85121 10989
rect 85149 10961 94917 10989
rect 94945 10961 94979 10989
rect 95007 10961 95041 10989
rect 95069 10961 95103 10989
rect 95131 10961 100419 10989
rect 100447 10961 100481 10989
rect 100509 10961 110277 10989
rect 110305 10961 110339 10989
rect 110367 10961 110401 10989
rect 110429 10961 110463 10989
rect 110491 10961 115779 10989
rect 115807 10961 115841 10989
rect 115869 10961 125637 10989
rect 125665 10961 125699 10989
rect 125727 10961 125761 10989
rect 125789 10961 125823 10989
rect 125851 10961 131139 10989
rect 131167 10961 131201 10989
rect 131229 10961 140997 10989
rect 141025 10961 141059 10989
rect 141087 10961 141121 10989
rect 141149 10961 141183 10989
rect 141211 10961 146499 10989
rect 146527 10961 146561 10989
rect 146589 10961 156357 10989
rect 156385 10961 156419 10989
rect 156447 10961 156481 10989
rect 156509 10961 156543 10989
rect 156571 10961 161859 10989
rect 161887 10961 161921 10989
rect 161949 10961 171717 10989
rect 171745 10961 171779 10989
rect 171807 10961 171841 10989
rect 171869 10961 171903 10989
rect 171931 10961 177219 10989
rect 177247 10961 177281 10989
rect 177309 10961 187077 10989
rect 187105 10961 187139 10989
rect 187167 10961 187201 10989
rect 187229 10961 187263 10989
rect 187291 10961 192579 10989
rect 192607 10961 192641 10989
rect 192669 10961 202437 10989
rect 202465 10961 202499 10989
rect 202527 10961 202561 10989
rect 202589 10961 202623 10989
rect 202651 10961 207939 10989
rect 207967 10961 208001 10989
rect 208029 10961 217797 10989
rect 217825 10961 217859 10989
rect 217887 10961 217921 10989
rect 217949 10961 217983 10989
rect 218011 10961 223299 10989
rect 223327 10961 223361 10989
rect 223389 10961 233157 10989
rect 233185 10961 233219 10989
rect 233247 10961 233281 10989
rect 233309 10961 233343 10989
rect 233371 10961 238659 10989
rect 238687 10961 238721 10989
rect 238749 10961 248517 10989
rect 248545 10961 248579 10989
rect 248607 10961 248641 10989
rect 248669 10961 248703 10989
rect 248731 10961 254019 10989
rect 254047 10961 254081 10989
rect 254109 10961 263877 10989
rect 263905 10961 263939 10989
rect 263967 10961 264001 10989
rect 264029 10961 264063 10989
rect 264091 10961 269379 10989
rect 269407 10961 269441 10989
rect 269469 10961 279237 10989
rect 279265 10961 279299 10989
rect 279327 10961 279361 10989
rect 279389 10961 279423 10989
rect 279451 10961 284739 10989
rect 284767 10961 284801 10989
rect 284829 10961 294597 10989
rect 294625 10961 294659 10989
rect 294687 10961 294721 10989
rect 294749 10961 294783 10989
rect 294811 10961 298248 10989
rect 298276 10961 298310 10989
rect 298338 10961 298372 10989
rect 298400 10961 298434 10989
rect 298462 10961 298990 10989
rect -958 10913 298990 10961
rect -958 5175 298990 5223
rect -958 5147 -910 5175
rect -882 5147 -848 5175
rect -820 5147 -786 5175
rect -758 5147 -724 5175
rect -696 5147 4617 5175
rect 4645 5147 4679 5175
rect 4707 5147 4741 5175
rect 4769 5147 4803 5175
rect 4831 5147 15939 5175
rect 15967 5147 16001 5175
rect 16029 5147 19977 5175
rect 20005 5147 20039 5175
rect 20067 5147 20101 5175
rect 20129 5147 20163 5175
rect 20191 5147 31299 5175
rect 31327 5147 31361 5175
rect 31389 5147 35337 5175
rect 35365 5147 35399 5175
rect 35427 5147 35461 5175
rect 35489 5147 35523 5175
rect 35551 5147 46659 5175
rect 46687 5147 46721 5175
rect 46749 5147 50697 5175
rect 50725 5147 50759 5175
rect 50787 5147 50821 5175
rect 50849 5147 50883 5175
rect 50911 5147 62019 5175
rect 62047 5147 62081 5175
rect 62109 5147 66057 5175
rect 66085 5147 66119 5175
rect 66147 5147 66181 5175
rect 66209 5147 66243 5175
rect 66271 5147 77379 5175
rect 77407 5147 77441 5175
rect 77469 5147 81417 5175
rect 81445 5147 81479 5175
rect 81507 5147 81541 5175
rect 81569 5147 81603 5175
rect 81631 5147 92739 5175
rect 92767 5147 92801 5175
rect 92829 5147 96777 5175
rect 96805 5147 96839 5175
rect 96867 5147 96901 5175
rect 96929 5147 96963 5175
rect 96991 5147 108099 5175
rect 108127 5147 108161 5175
rect 108189 5147 112137 5175
rect 112165 5147 112199 5175
rect 112227 5147 112261 5175
rect 112289 5147 112323 5175
rect 112351 5147 123459 5175
rect 123487 5147 123521 5175
rect 123549 5147 127497 5175
rect 127525 5147 127559 5175
rect 127587 5147 127621 5175
rect 127649 5147 127683 5175
rect 127711 5147 138819 5175
rect 138847 5147 138881 5175
rect 138909 5147 142857 5175
rect 142885 5147 142919 5175
rect 142947 5147 142981 5175
rect 143009 5147 143043 5175
rect 143071 5147 154179 5175
rect 154207 5147 154241 5175
rect 154269 5147 158217 5175
rect 158245 5147 158279 5175
rect 158307 5147 158341 5175
rect 158369 5147 158403 5175
rect 158431 5147 169539 5175
rect 169567 5147 169601 5175
rect 169629 5147 173577 5175
rect 173605 5147 173639 5175
rect 173667 5147 173701 5175
rect 173729 5147 173763 5175
rect 173791 5147 184899 5175
rect 184927 5147 184961 5175
rect 184989 5147 188937 5175
rect 188965 5147 188999 5175
rect 189027 5147 189061 5175
rect 189089 5147 189123 5175
rect 189151 5147 200259 5175
rect 200287 5147 200321 5175
rect 200349 5147 204297 5175
rect 204325 5147 204359 5175
rect 204387 5147 204421 5175
rect 204449 5147 204483 5175
rect 204511 5147 215619 5175
rect 215647 5147 215681 5175
rect 215709 5147 219657 5175
rect 219685 5147 219719 5175
rect 219747 5147 219781 5175
rect 219809 5147 219843 5175
rect 219871 5147 230979 5175
rect 231007 5147 231041 5175
rect 231069 5147 235017 5175
rect 235045 5147 235079 5175
rect 235107 5147 235141 5175
rect 235169 5147 235203 5175
rect 235231 5147 246339 5175
rect 246367 5147 246401 5175
rect 246429 5147 250377 5175
rect 250405 5147 250439 5175
rect 250467 5147 250501 5175
rect 250529 5147 250563 5175
rect 250591 5147 261699 5175
rect 261727 5147 261761 5175
rect 261789 5147 265737 5175
rect 265765 5147 265799 5175
rect 265827 5147 265861 5175
rect 265889 5147 265923 5175
rect 265951 5147 277059 5175
rect 277087 5147 277121 5175
rect 277149 5147 281097 5175
rect 281125 5147 281159 5175
rect 281187 5147 281221 5175
rect 281249 5147 281283 5175
rect 281311 5147 296457 5175
rect 296485 5147 296519 5175
rect 296547 5147 296581 5175
rect 296609 5147 296643 5175
rect 296671 5147 298728 5175
rect 298756 5147 298790 5175
rect 298818 5147 298852 5175
rect 298880 5147 298914 5175
rect 298942 5147 298990 5175
rect -958 5113 298990 5147
rect -958 5085 -910 5113
rect -882 5085 -848 5113
rect -820 5085 -786 5113
rect -758 5085 -724 5113
rect -696 5085 4617 5113
rect 4645 5085 4679 5113
rect 4707 5085 4741 5113
rect 4769 5085 4803 5113
rect 4831 5085 15939 5113
rect 15967 5085 16001 5113
rect 16029 5085 19977 5113
rect 20005 5085 20039 5113
rect 20067 5085 20101 5113
rect 20129 5085 20163 5113
rect 20191 5085 31299 5113
rect 31327 5085 31361 5113
rect 31389 5085 35337 5113
rect 35365 5085 35399 5113
rect 35427 5085 35461 5113
rect 35489 5085 35523 5113
rect 35551 5085 46659 5113
rect 46687 5085 46721 5113
rect 46749 5085 50697 5113
rect 50725 5085 50759 5113
rect 50787 5085 50821 5113
rect 50849 5085 50883 5113
rect 50911 5085 62019 5113
rect 62047 5085 62081 5113
rect 62109 5085 66057 5113
rect 66085 5085 66119 5113
rect 66147 5085 66181 5113
rect 66209 5085 66243 5113
rect 66271 5085 77379 5113
rect 77407 5085 77441 5113
rect 77469 5085 81417 5113
rect 81445 5085 81479 5113
rect 81507 5085 81541 5113
rect 81569 5085 81603 5113
rect 81631 5085 92739 5113
rect 92767 5085 92801 5113
rect 92829 5085 96777 5113
rect 96805 5085 96839 5113
rect 96867 5085 96901 5113
rect 96929 5085 96963 5113
rect 96991 5085 108099 5113
rect 108127 5085 108161 5113
rect 108189 5085 112137 5113
rect 112165 5085 112199 5113
rect 112227 5085 112261 5113
rect 112289 5085 112323 5113
rect 112351 5085 123459 5113
rect 123487 5085 123521 5113
rect 123549 5085 127497 5113
rect 127525 5085 127559 5113
rect 127587 5085 127621 5113
rect 127649 5085 127683 5113
rect 127711 5085 138819 5113
rect 138847 5085 138881 5113
rect 138909 5085 142857 5113
rect 142885 5085 142919 5113
rect 142947 5085 142981 5113
rect 143009 5085 143043 5113
rect 143071 5085 154179 5113
rect 154207 5085 154241 5113
rect 154269 5085 158217 5113
rect 158245 5085 158279 5113
rect 158307 5085 158341 5113
rect 158369 5085 158403 5113
rect 158431 5085 169539 5113
rect 169567 5085 169601 5113
rect 169629 5085 173577 5113
rect 173605 5085 173639 5113
rect 173667 5085 173701 5113
rect 173729 5085 173763 5113
rect 173791 5085 184899 5113
rect 184927 5085 184961 5113
rect 184989 5085 188937 5113
rect 188965 5085 188999 5113
rect 189027 5085 189061 5113
rect 189089 5085 189123 5113
rect 189151 5085 200259 5113
rect 200287 5085 200321 5113
rect 200349 5085 204297 5113
rect 204325 5085 204359 5113
rect 204387 5085 204421 5113
rect 204449 5085 204483 5113
rect 204511 5085 215619 5113
rect 215647 5085 215681 5113
rect 215709 5085 219657 5113
rect 219685 5085 219719 5113
rect 219747 5085 219781 5113
rect 219809 5085 219843 5113
rect 219871 5085 230979 5113
rect 231007 5085 231041 5113
rect 231069 5085 235017 5113
rect 235045 5085 235079 5113
rect 235107 5085 235141 5113
rect 235169 5085 235203 5113
rect 235231 5085 246339 5113
rect 246367 5085 246401 5113
rect 246429 5085 250377 5113
rect 250405 5085 250439 5113
rect 250467 5085 250501 5113
rect 250529 5085 250563 5113
rect 250591 5085 261699 5113
rect 261727 5085 261761 5113
rect 261789 5085 265737 5113
rect 265765 5085 265799 5113
rect 265827 5085 265861 5113
rect 265889 5085 265923 5113
rect 265951 5085 277059 5113
rect 277087 5085 277121 5113
rect 277149 5085 281097 5113
rect 281125 5085 281159 5113
rect 281187 5085 281221 5113
rect 281249 5085 281283 5113
rect 281311 5085 296457 5113
rect 296485 5085 296519 5113
rect 296547 5085 296581 5113
rect 296609 5085 296643 5113
rect 296671 5085 298728 5113
rect 298756 5085 298790 5113
rect 298818 5085 298852 5113
rect 298880 5085 298914 5113
rect 298942 5085 298990 5113
rect -958 5051 298990 5085
rect -958 5023 -910 5051
rect -882 5023 -848 5051
rect -820 5023 -786 5051
rect -758 5023 -724 5051
rect -696 5023 4617 5051
rect 4645 5023 4679 5051
rect 4707 5023 4741 5051
rect 4769 5023 4803 5051
rect 4831 5023 15939 5051
rect 15967 5023 16001 5051
rect 16029 5023 19977 5051
rect 20005 5023 20039 5051
rect 20067 5023 20101 5051
rect 20129 5023 20163 5051
rect 20191 5023 31299 5051
rect 31327 5023 31361 5051
rect 31389 5023 35337 5051
rect 35365 5023 35399 5051
rect 35427 5023 35461 5051
rect 35489 5023 35523 5051
rect 35551 5023 46659 5051
rect 46687 5023 46721 5051
rect 46749 5023 50697 5051
rect 50725 5023 50759 5051
rect 50787 5023 50821 5051
rect 50849 5023 50883 5051
rect 50911 5023 62019 5051
rect 62047 5023 62081 5051
rect 62109 5023 66057 5051
rect 66085 5023 66119 5051
rect 66147 5023 66181 5051
rect 66209 5023 66243 5051
rect 66271 5023 77379 5051
rect 77407 5023 77441 5051
rect 77469 5023 81417 5051
rect 81445 5023 81479 5051
rect 81507 5023 81541 5051
rect 81569 5023 81603 5051
rect 81631 5023 92739 5051
rect 92767 5023 92801 5051
rect 92829 5023 96777 5051
rect 96805 5023 96839 5051
rect 96867 5023 96901 5051
rect 96929 5023 96963 5051
rect 96991 5023 108099 5051
rect 108127 5023 108161 5051
rect 108189 5023 112137 5051
rect 112165 5023 112199 5051
rect 112227 5023 112261 5051
rect 112289 5023 112323 5051
rect 112351 5023 123459 5051
rect 123487 5023 123521 5051
rect 123549 5023 127497 5051
rect 127525 5023 127559 5051
rect 127587 5023 127621 5051
rect 127649 5023 127683 5051
rect 127711 5023 138819 5051
rect 138847 5023 138881 5051
rect 138909 5023 142857 5051
rect 142885 5023 142919 5051
rect 142947 5023 142981 5051
rect 143009 5023 143043 5051
rect 143071 5023 154179 5051
rect 154207 5023 154241 5051
rect 154269 5023 158217 5051
rect 158245 5023 158279 5051
rect 158307 5023 158341 5051
rect 158369 5023 158403 5051
rect 158431 5023 169539 5051
rect 169567 5023 169601 5051
rect 169629 5023 173577 5051
rect 173605 5023 173639 5051
rect 173667 5023 173701 5051
rect 173729 5023 173763 5051
rect 173791 5023 184899 5051
rect 184927 5023 184961 5051
rect 184989 5023 188937 5051
rect 188965 5023 188999 5051
rect 189027 5023 189061 5051
rect 189089 5023 189123 5051
rect 189151 5023 200259 5051
rect 200287 5023 200321 5051
rect 200349 5023 204297 5051
rect 204325 5023 204359 5051
rect 204387 5023 204421 5051
rect 204449 5023 204483 5051
rect 204511 5023 215619 5051
rect 215647 5023 215681 5051
rect 215709 5023 219657 5051
rect 219685 5023 219719 5051
rect 219747 5023 219781 5051
rect 219809 5023 219843 5051
rect 219871 5023 230979 5051
rect 231007 5023 231041 5051
rect 231069 5023 235017 5051
rect 235045 5023 235079 5051
rect 235107 5023 235141 5051
rect 235169 5023 235203 5051
rect 235231 5023 246339 5051
rect 246367 5023 246401 5051
rect 246429 5023 250377 5051
rect 250405 5023 250439 5051
rect 250467 5023 250501 5051
rect 250529 5023 250563 5051
rect 250591 5023 261699 5051
rect 261727 5023 261761 5051
rect 261789 5023 265737 5051
rect 265765 5023 265799 5051
rect 265827 5023 265861 5051
rect 265889 5023 265923 5051
rect 265951 5023 277059 5051
rect 277087 5023 277121 5051
rect 277149 5023 281097 5051
rect 281125 5023 281159 5051
rect 281187 5023 281221 5051
rect 281249 5023 281283 5051
rect 281311 5023 296457 5051
rect 296485 5023 296519 5051
rect 296547 5023 296581 5051
rect 296609 5023 296643 5051
rect 296671 5023 298728 5051
rect 298756 5023 298790 5051
rect 298818 5023 298852 5051
rect 298880 5023 298914 5051
rect 298942 5023 298990 5051
rect -958 4989 298990 5023
rect -958 4961 -910 4989
rect -882 4961 -848 4989
rect -820 4961 -786 4989
rect -758 4961 -724 4989
rect -696 4961 4617 4989
rect 4645 4961 4679 4989
rect 4707 4961 4741 4989
rect 4769 4961 4803 4989
rect 4831 4961 15939 4989
rect 15967 4961 16001 4989
rect 16029 4961 19977 4989
rect 20005 4961 20039 4989
rect 20067 4961 20101 4989
rect 20129 4961 20163 4989
rect 20191 4961 31299 4989
rect 31327 4961 31361 4989
rect 31389 4961 35337 4989
rect 35365 4961 35399 4989
rect 35427 4961 35461 4989
rect 35489 4961 35523 4989
rect 35551 4961 46659 4989
rect 46687 4961 46721 4989
rect 46749 4961 50697 4989
rect 50725 4961 50759 4989
rect 50787 4961 50821 4989
rect 50849 4961 50883 4989
rect 50911 4961 62019 4989
rect 62047 4961 62081 4989
rect 62109 4961 66057 4989
rect 66085 4961 66119 4989
rect 66147 4961 66181 4989
rect 66209 4961 66243 4989
rect 66271 4961 77379 4989
rect 77407 4961 77441 4989
rect 77469 4961 81417 4989
rect 81445 4961 81479 4989
rect 81507 4961 81541 4989
rect 81569 4961 81603 4989
rect 81631 4961 92739 4989
rect 92767 4961 92801 4989
rect 92829 4961 96777 4989
rect 96805 4961 96839 4989
rect 96867 4961 96901 4989
rect 96929 4961 96963 4989
rect 96991 4961 108099 4989
rect 108127 4961 108161 4989
rect 108189 4961 112137 4989
rect 112165 4961 112199 4989
rect 112227 4961 112261 4989
rect 112289 4961 112323 4989
rect 112351 4961 123459 4989
rect 123487 4961 123521 4989
rect 123549 4961 127497 4989
rect 127525 4961 127559 4989
rect 127587 4961 127621 4989
rect 127649 4961 127683 4989
rect 127711 4961 138819 4989
rect 138847 4961 138881 4989
rect 138909 4961 142857 4989
rect 142885 4961 142919 4989
rect 142947 4961 142981 4989
rect 143009 4961 143043 4989
rect 143071 4961 154179 4989
rect 154207 4961 154241 4989
rect 154269 4961 158217 4989
rect 158245 4961 158279 4989
rect 158307 4961 158341 4989
rect 158369 4961 158403 4989
rect 158431 4961 169539 4989
rect 169567 4961 169601 4989
rect 169629 4961 173577 4989
rect 173605 4961 173639 4989
rect 173667 4961 173701 4989
rect 173729 4961 173763 4989
rect 173791 4961 184899 4989
rect 184927 4961 184961 4989
rect 184989 4961 188937 4989
rect 188965 4961 188999 4989
rect 189027 4961 189061 4989
rect 189089 4961 189123 4989
rect 189151 4961 200259 4989
rect 200287 4961 200321 4989
rect 200349 4961 204297 4989
rect 204325 4961 204359 4989
rect 204387 4961 204421 4989
rect 204449 4961 204483 4989
rect 204511 4961 215619 4989
rect 215647 4961 215681 4989
rect 215709 4961 219657 4989
rect 219685 4961 219719 4989
rect 219747 4961 219781 4989
rect 219809 4961 219843 4989
rect 219871 4961 230979 4989
rect 231007 4961 231041 4989
rect 231069 4961 235017 4989
rect 235045 4961 235079 4989
rect 235107 4961 235141 4989
rect 235169 4961 235203 4989
rect 235231 4961 246339 4989
rect 246367 4961 246401 4989
rect 246429 4961 250377 4989
rect 250405 4961 250439 4989
rect 250467 4961 250501 4989
rect 250529 4961 250563 4989
rect 250591 4961 261699 4989
rect 261727 4961 261761 4989
rect 261789 4961 265737 4989
rect 265765 4961 265799 4989
rect 265827 4961 265861 4989
rect 265889 4961 265923 4989
rect 265951 4961 277059 4989
rect 277087 4961 277121 4989
rect 277149 4961 281097 4989
rect 281125 4961 281159 4989
rect 281187 4961 281221 4989
rect 281249 4961 281283 4989
rect 281311 4961 296457 4989
rect 296485 4961 296519 4989
rect 296547 4961 296581 4989
rect 296609 4961 296643 4989
rect 296671 4961 298728 4989
rect 298756 4961 298790 4989
rect 298818 4961 298852 4989
rect 298880 4961 298914 4989
rect 298942 4961 298990 4989
rect -958 4913 298990 4961
rect -958 2175 298990 2223
rect -958 2147 -430 2175
rect -402 2147 -368 2175
rect -340 2147 -306 2175
rect -278 2147 -244 2175
rect -216 2147 2757 2175
rect 2785 2147 2819 2175
rect 2847 2147 2881 2175
rect 2909 2147 2943 2175
rect 2971 2147 18117 2175
rect 18145 2147 18179 2175
rect 18207 2147 18241 2175
rect 18269 2147 18303 2175
rect 18331 2147 33477 2175
rect 33505 2147 33539 2175
rect 33567 2147 33601 2175
rect 33629 2147 33663 2175
rect 33691 2147 48837 2175
rect 48865 2147 48899 2175
rect 48927 2147 48961 2175
rect 48989 2147 49023 2175
rect 49051 2147 64197 2175
rect 64225 2147 64259 2175
rect 64287 2147 64321 2175
rect 64349 2147 64383 2175
rect 64411 2147 79557 2175
rect 79585 2147 79619 2175
rect 79647 2147 79681 2175
rect 79709 2147 79743 2175
rect 79771 2147 94917 2175
rect 94945 2147 94979 2175
rect 95007 2147 95041 2175
rect 95069 2147 95103 2175
rect 95131 2147 110277 2175
rect 110305 2147 110339 2175
rect 110367 2147 110401 2175
rect 110429 2147 110463 2175
rect 110491 2147 125637 2175
rect 125665 2147 125699 2175
rect 125727 2147 125761 2175
rect 125789 2147 125823 2175
rect 125851 2147 140997 2175
rect 141025 2147 141059 2175
rect 141087 2147 141121 2175
rect 141149 2147 141183 2175
rect 141211 2147 156357 2175
rect 156385 2147 156419 2175
rect 156447 2147 156481 2175
rect 156509 2147 156543 2175
rect 156571 2147 171717 2175
rect 171745 2147 171779 2175
rect 171807 2147 171841 2175
rect 171869 2147 171903 2175
rect 171931 2147 187077 2175
rect 187105 2147 187139 2175
rect 187167 2147 187201 2175
rect 187229 2147 187263 2175
rect 187291 2147 202437 2175
rect 202465 2147 202499 2175
rect 202527 2147 202561 2175
rect 202589 2147 202623 2175
rect 202651 2147 217797 2175
rect 217825 2147 217859 2175
rect 217887 2147 217921 2175
rect 217949 2147 217983 2175
rect 218011 2147 233157 2175
rect 233185 2147 233219 2175
rect 233247 2147 233281 2175
rect 233309 2147 233343 2175
rect 233371 2147 248517 2175
rect 248545 2147 248579 2175
rect 248607 2147 248641 2175
rect 248669 2147 248703 2175
rect 248731 2147 263877 2175
rect 263905 2147 263939 2175
rect 263967 2147 264001 2175
rect 264029 2147 264063 2175
rect 264091 2147 279237 2175
rect 279265 2147 279299 2175
rect 279327 2147 279361 2175
rect 279389 2147 279423 2175
rect 279451 2147 294597 2175
rect 294625 2147 294659 2175
rect 294687 2147 294721 2175
rect 294749 2147 294783 2175
rect 294811 2147 298248 2175
rect 298276 2147 298310 2175
rect 298338 2147 298372 2175
rect 298400 2147 298434 2175
rect 298462 2147 298990 2175
rect -958 2113 298990 2147
rect -958 2085 -430 2113
rect -402 2085 -368 2113
rect -340 2085 -306 2113
rect -278 2085 -244 2113
rect -216 2085 2757 2113
rect 2785 2085 2819 2113
rect 2847 2085 2881 2113
rect 2909 2085 2943 2113
rect 2971 2085 18117 2113
rect 18145 2085 18179 2113
rect 18207 2085 18241 2113
rect 18269 2085 18303 2113
rect 18331 2085 33477 2113
rect 33505 2085 33539 2113
rect 33567 2085 33601 2113
rect 33629 2085 33663 2113
rect 33691 2085 48837 2113
rect 48865 2085 48899 2113
rect 48927 2085 48961 2113
rect 48989 2085 49023 2113
rect 49051 2085 64197 2113
rect 64225 2085 64259 2113
rect 64287 2085 64321 2113
rect 64349 2085 64383 2113
rect 64411 2085 79557 2113
rect 79585 2085 79619 2113
rect 79647 2085 79681 2113
rect 79709 2085 79743 2113
rect 79771 2085 94917 2113
rect 94945 2085 94979 2113
rect 95007 2085 95041 2113
rect 95069 2085 95103 2113
rect 95131 2085 110277 2113
rect 110305 2085 110339 2113
rect 110367 2085 110401 2113
rect 110429 2085 110463 2113
rect 110491 2085 125637 2113
rect 125665 2085 125699 2113
rect 125727 2085 125761 2113
rect 125789 2085 125823 2113
rect 125851 2085 140997 2113
rect 141025 2085 141059 2113
rect 141087 2085 141121 2113
rect 141149 2085 141183 2113
rect 141211 2085 156357 2113
rect 156385 2085 156419 2113
rect 156447 2085 156481 2113
rect 156509 2085 156543 2113
rect 156571 2085 171717 2113
rect 171745 2085 171779 2113
rect 171807 2085 171841 2113
rect 171869 2085 171903 2113
rect 171931 2085 187077 2113
rect 187105 2085 187139 2113
rect 187167 2085 187201 2113
rect 187229 2085 187263 2113
rect 187291 2085 202437 2113
rect 202465 2085 202499 2113
rect 202527 2085 202561 2113
rect 202589 2085 202623 2113
rect 202651 2085 217797 2113
rect 217825 2085 217859 2113
rect 217887 2085 217921 2113
rect 217949 2085 217983 2113
rect 218011 2085 233157 2113
rect 233185 2085 233219 2113
rect 233247 2085 233281 2113
rect 233309 2085 233343 2113
rect 233371 2085 248517 2113
rect 248545 2085 248579 2113
rect 248607 2085 248641 2113
rect 248669 2085 248703 2113
rect 248731 2085 263877 2113
rect 263905 2085 263939 2113
rect 263967 2085 264001 2113
rect 264029 2085 264063 2113
rect 264091 2085 279237 2113
rect 279265 2085 279299 2113
rect 279327 2085 279361 2113
rect 279389 2085 279423 2113
rect 279451 2085 294597 2113
rect 294625 2085 294659 2113
rect 294687 2085 294721 2113
rect 294749 2085 294783 2113
rect 294811 2085 298248 2113
rect 298276 2085 298310 2113
rect 298338 2085 298372 2113
rect 298400 2085 298434 2113
rect 298462 2085 298990 2113
rect -958 2051 298990 2085
rect -958 2023 -430 2051
rect -402 2023 -368 2051
rect -340 2023 -306 2051
rect -278 2023 -244 2051
rect -216 2023 2757 2051
rect 2785 2023 2819 2051
rect 2847 2023 2881 2051
rect 2909 2023 2943 2051
rect 2971 2023 18117 2051
rect 18145 2023 18179 2051
rect 18207 2023 18241 2051
rect 18269 2023 18303 2051
rect 18331 2023 33477 2051
rect 33505 2023 33539 2051
rect 33567 2023 33601 2051
rect 33629 2023 33663 2051
rect 33691 2023 48837 2051
rect 48865 2023 48899 2051
rect 48927 2023 48961 2051
rect 48989 2023 49023 2051
rect 49051 2023 64197 2051
rect 64225 2023 64259 2051
rect 64287 2023 64321 2051
rect 64349 2023 64383 2051
rect 64411 2023 79557 2051
rect 79585 2023 79619 2051
rect 79647 2023 79681 2051
rect 79709 2023 79743 2051
rect 79771 2023 94917 2051
rect 94945 2023 94979 2051
rect 95007 2023 95041 2051
rect 95069 2023 95103 2051
rect 95131 2023 110277 2051
rect 110305 2023 110339 2051
rect 110367 2023 110401 2051
rect 110429 2023 110463 2051
rect 110491 2023 125637 2051
rect 125665 2023 125699 2051
rect 125727 2023 125761 2051
rect 125789 2023 125823 2051
rect 125851 2023 140997 2051
rect 141025 2023 141059 2051
rect 141087 2023 141121 2051
rect 141149 2023 141183 2051
rect 141211 2023 156357 2051
rect 156385 2023 156419 2051
rect 156447 2023 156481 2051
rect 156509 2023 156543 2051
rect 156571 2023 171717 2051
rect 171745 2023 171779 2051
rect 171807 2023 171841 2051
rect 171869 2023 171903 2051
rect 171931 2023 187077 2051
rect 187105 2023 187139 2051
rect 187167 2023 187201 2051
rect 187229 2023 187263 2051
rect 187291 2023 202437 2051
rect 202465 2023 202499 2051
rect 202527 2023 202561 2051
rect 202589 2023 202623 2051
rect 202651 2023 217797 2051
rect 217825 2023 217859 2051
rect 217887 2023 217921 2051
rect 217949 2023 217983 2051
rect 218011 2023 233157 2051
rect 233185 2023 233219 2051
rect 233247 2023 233281 2051
rect 233309 2023 233343 2051
rect 233371 2023 248517 2051
rect 248545 2023 248579 2051
rect 248607 2023 248641 2051
rect 248669 2023 248703 2051
rect 248731 2023 263877 2051
rect 263905 2023 263939 2051
rect 263967 2023 264001 2051
rect 264029 2023 264063 2051
rect 264091 2023 279237 2051
rect 279265 2023 279299 2051
rect 279327 2023 279361 2051
rect 279389 2023 279423 2051
rect 279451 2023 294597 2051
rect 294625 2023 294659 2051
rect 294687 2023 294721 2051
rect 294749 2023 294783 2051
rect 294811 2023 298248 2051
rect 298276 2023 298310 2051
rect 298338 2023 298372 2051
rect 298400 2023 298434 2051
rect 298462 2023 298990 2051
rect -958 1989 298990 2023
rect -958 1961 -430 1989
rect -402 1961 -368 1989
rect -340 1961 -306 1989
rect -278 1961 -244 1989
rect -216 1961 2757 1989
rect 2785 1961 2819 1989
rect 2847 1961 2881 1989
rect 2909 1961 2943 1989
rect 2971 1961 18117 1989
rect 18145 1961 18179 1989
rect 18207 1961 18241 1989
rect 18269 1961 18303 1989
rect 18331 1961 33477 1989
rect 33505 1961 33539 1989
rect 33567 1961 33601 1989
rect 33629 1961 33663 1989
rect 33691 1961 48837 1989
rect 48865 1961 48899 1989
rect 48927 1961 48961 1989
rect 48989 1961 49023 1989
rect 49051 1961 64197 1989
rect 64225 1961 64259 1989
rect 64287 1961 64321 1989
rect 64349 1961 64383 1989
rect 64411 1961 79557 1989
rect 79585 1961 79619 1989
rect 79647 1961 79681 1989
rect 79709 1961 79743 1989
rect 79771 1961 94917 1989
rect 94945 1961 94979 1989
rect 95007 1961 95041 1989
rect 95069 1961 95103 1989
rect 95131 1961 110277 1989
rect 110305 1961 110339 1989
rect 110367 1961 110401 1989
rect 110429 1961 110463 1989
rect 110491 1961 125637 1989
rect 125665 1961 125699 1989
rect 125727 1961 125761 1989
rect 125789 1961 125823 1989
rect 125851 1961 140997 1989
rect 141025 1961 141059 1989
rect 141087 1961 141121 1989
rect 141149 1961 141183 1989
rect 141211 1961 156357 1989
rect 156385 1961 156419 1989
rect 156447 1961 156481 1989
rect 156509 1961 156543 1989
rect 156571 1961 171717 1989
rect 171745 1961 171779 1989
rect 171807 1961 171841 1989
rect 171869 1961 171903 1989
rect 171931 1961 187077 1989
rect 187105 1961 187139 1989
rect 187167 1961 187201 1989
rect 187229 1961 187263 1989
rect 187291 1961 202437 1989
rect 202465 1961 202499 1989
rect 202527 1961 202561 1989
rect 202589 1961 202623 1989
rect 202651 1961 217797 1989
rect 217825 1961 217859 1989
rect 217887 1961 217921 1989
rect 217949 1961 217983 1989
rect 218011 1961 233157 1989
rect 233185 1961 233219 1989
rect 233247 1961 233281 1989
rect 233309 1961 233343 1989
rect 233371 1961 248517 1989
rect 248545 1961 248579 1989
rect 248607 1961 248641 1989
rect 248669 1961 248703 1989
rect 248731 1961 263877 1989
rect 263905 1961 263939 1989
rect 263967 1961 264001 1989
rect 264029 1961 264063 1989
rect 264091 1961 279237 1989
rect 279265 1961 279299 1989
rect 279327 1961 279361 1989
rect 279389 1961 279423 1989
rect 279451 1961 294597 1989
rect 294625 1961 294659 1989
rect 294687 1961 294721 1989
rect 294749 1961 294783 1989
rect 294811 1961 298248 1989
rect 298276 1961 298310 1989
rect 298338 1961 298372 1989
rect 298400 1961 298434 1989
rect 298462 1961 298990 1989
rect -958 1913 298990 1961
rect -478 -80 298510 -32
rect -478 -108 -430 -80
rect -402 -108 -368 -80
rect -340 -108 -306 -80
rect -278 -108 -244 -80
rect -216 -108 2757 -80
rect 2785 -108 2819 -80
rect 2847 -108 2881 -80
rect 2909 -108 2943 -80
rect 2971 -108 18117 -80
rect 18145 -108 18179 -80
rect 18207 -108 18241 -80
rect 18269 -108 18303 -80
rect 18331 -108 33477 -80
rect 33505 -108 33539 -80
rect 33567 -108 33601 -80
rect 33629 -108 33663 -80
rect 33691 -108 48837 -80
rect 48865 -108 48899 -80
rect 48927 -108 48961 -80
rect 48989 -108 49023 -80
rect 49051 -108 64197 -80
rect 64225 -108 64259 -80
rect 64287 -108 64321 -80
rect 64349 -108 64383 -80
rect 64411 -108 79557 -80
rect 79585 -108 79619 -80
rect 79647 -108 79681 -80
rect 79709 -108 79743 -80
rect 79771 -108 94917 -80
rect 94945 -108 94979 -80
rect 95007 -108 95041 -80
rect 95069 -108 95103 -80
rect 95131 -108 110277 -80
rect 110305 -108 110339 -80
rect 110367 -108 110401 -80
rect 110429 -108 110463 -80
rect 110491 -108 125637 -80
rect 125665 -108 125699 -80
rect 125727 -108 125761 -80
rect 125789 -108 125823 -80
rect 125851 -108 140997 -80
rect 141025 -108 141059 -80
rect 141087 -108 141121 -80
rect 141149 -108 141183 -80
rect 141211 -108 156357 -80
rect 156385 -108 156419 -80
rect 156447 -108 156481 -80
rect 156509 -108 156543 -80
rect 156571 -108 171717 -80
rect 171745 -108 171779 -80
rect 171807 -108 171841 -80
rect 171869 -108 171903 -80
rect 171931 -108 187077 -80
rect 187105 -108 187139 -80
rect 187167 -108 187201 -80
rect 187229 -108 187263 -80
rect 187291 -108 202437 -80
rect 202465 -108 202499 -80
rect 202527 -108 202561 -80
rect 202589 -108 202623 -80
rect 202651 -108 217797 -80
rect 217825 -108 217859 -80
rect 217887 -108 217921 -80
rect 217949 -108 217983 -80
rect 218011 -108 233157 -80
rect 233185 -108 233219 -80
rect 233247 -108 233281 -80
rect 233309 -108 233343 -80
rect 233371 -108 248517 -80
rect 248545 -108 248579 -80
rect 248607 -108 248641 -80
rect 248669 -108 248703 -80
rect 248731 -108 263877 -80
rect 263905 -108 263939 -80
rect 263967 -108 264001 -80
rect 264029 -108 264063 -80
rect 264091 -108 279237 -80
rect 279265 -108 279299 -80
rect 279327 -108 279361 -80
rect 279389 -108 279423 -80
rect 279451 -108 294597 -80
rect 294625 -108 294659 -80
rect 294687 -108 294721 -80
rect 294749 -108 294783 -80
rect 294811 -108 298248 -80
rect 298276 -108 298310 -80
rect 298338 -108 298372 -80
rect 298400 -108 298434 -80
rect 298462 -108 298510 -80
rect -478 -142 298510 -108
rect -478 -170 -430 -142
rect -402 -170 -368 -142
rect -340 -170 -306 -142
rect -278 -170 -244 -142
rect -216 -170 2757 -142
rect 2785 -170 2819 -142
rect 2847 -170 2881 -142
rect 2909 -170 2943 -142
rect 2971 -170 18117 -142
rect 18145 -170 18179 -142
rect 18207 -170 18241 -142
rect 18269 -170 18303 -142
rect 18331 -170 33477 -142
rect 33505 -170 33539 -142
rect 33567 -170 33601 -142
rect 33629 -170 33663 -142
rect 33691 -170 48837 -142
rect 48865 -170 48899 -142
rect 48927 -170 48961 -142
rect 48989 -170 49023 -142
rect 49051 -170 64197 -142
rect 64225 -170 64259 -142
rect 64287 -170 64321 -142
rect 64349 -170 64383 -142
rect 64411 -170 79557 -142
rect 79585 -170 79619 -142
rect 79647 -170 79681 -142
rect 79709 -170 79743 -142
rect 79771 -170 94917 -142
rect 94945 -170 94979 -142
rect 95007 -170 95041 -142
rect 95069 -170 95103 -142
rect 95131 -170 110277 -142
rect 110305 -170 110339 -142
rect 110367 -170 110401 -142
rect 110429 -170 110463 -142
rect 110491 -170 125637 -142
rect 125665 -170 125699 -142
rect 125727 -170 125761 -142
rect 125789 -170 125823 -142
rect 125851 -170 140997 -142
rect 141025 -170 141059 -142
rect 141087 -170 141121 -142
rect 141149 -170 141183 -142
rect 141211 -170 156357 -142
rect 156385 -170 156419 -142
rect 156447 -170 156481 -142
rect 156509 -170 156543 -142
rect 156571 -170 171717 -142
rect 171745 -170 171779 -142
rect 171807 -170 171841 -142
rect 171869 -170 171903 -142
rect 171931 -170 187077 -142
rect 187105 -170 187139 -142
rect 187167 -170 187201 -142
rect 187229 -170 187263 -142
rect 187291 -170 202437 -142
rect 202465 -170 202499 -142
rect 202527 -170 202561 -142
rect 202589 -170 202623 -142
rect 202651 -170 217797 -142
rect 217825 -170 217859 -142
rect 217887 -170 217921 -142
rect 217949 -170 217983 -142
rect 218011 -170 233157 -142
rect 233185 -170 233219 -142
rect 233247 -170 233281 -142
rect 233309 -170 233343 -142
rect 233371 -170 248517 -142
rect 248545 -170 248579 -142
rect 248607 -170 248641 -142
rect 248669 -170 248703 -142
rect 248731 -170 263877 -142
rect 263905 -170 263939 -142
rect 263967 -170 264001 -142
rect 264029 -170 264063 -142
rect 264091 -170 279237 -142
rect 279265 -170 279299 -142
rect 279327 -170 279361 -142
rect 279389 -170 279423 -142
rect 279451 -170 294597 -142
rect 294625 -170 294659 -142
rect 294687 -170 294721 -142
rect 294749 -170 294783 -142
rect 294811 -170 298248 -142
rect 298276 -170 298310 -142
rect 298338 -170 298372 -142
rect 298400 -170 298434 -142
rect 298462 -170 298510 -142
rect -478 -204 298510 -170
rect -478 -232 -430 -204
rect -402 -232 -368 -204
rect -340 -232 -306 -204
rect -278 -232 -244 -204
rect -216 -232 2757 -204
rect 2785 -232 2819 -204
rect 2847 -232 2881 -204
rect 2909 -232 2943 -204
rect 2971 -232 18117 -204
rect 18145 -232 18179 -204
rect 18207 -232 18241 -204
rect 18269 -232 18303 -204
rect 18331 -232 33477 -204
rect 33505 -232 33539 -204
rect 33567 -232 33601 -204
rect 33629 -232 33663 -204
rect 33691 -232 48837 -204
rect 48865 -232 48899 -204
rect 48927 -232 48961 -204
rect 48989 -232 49023 -204
rect 49051 -232 64197 -204
rect 64225 -232 64259 -204
rect 64287 -232 64321 -204
rect 64349 -232 64383 -204
rect 64411 -232 79557 -204
rect 79585 -232 79619 -204
rect 79647 -232 79681 -204
rect 79709 -232 79743 -204
rect 79771 -232 94917 -204
rect 94945 -232 94979 -204
rect 95007 -232 95041 -204
rect 95069 -232 95103 -204
rect 95131 -232 110277 -204
rect 110305 -232 110339 -204
rect 110367 -232 110401 -204
rect 110429 -232 110463 -204
rect 110491 -232 125637 -204
rect 125665 -232 125699 -204
rect 125727 -232 125761 -204
rect 125789 -232 125823 -204
rect 125851 -232 140997 -204
rect 141025 -232 141059 -204
rect 141087 -232 141121 -204
rect 141149 -232 141183 -204
rect 141211 -232 156357 -204
rect 156385 -232 156419 -204
rect 156447 -232 156481 -204
rect 156509 -232 156543 -204
rect 156571 -232 171717 -204
rect 171745 -232 171779 -204
rect 171807 -232 171841 -204
rect 171869 -232 171903 -204
rect 171931 -232 187077 -204
rect 187105 -232 187139 -204
rect 187167 -232 187201 -204
rect 187229 -232 187263 -204
rect 187291 -232 202437 -204
rect 202465 -232 202499 -204
rect 202527 -232 202561 -204
rect 202589 -232 202623 -204
rect 202651 -232 217797 -204
rect 217825 -232 217859 -204
rect 217887 -232 217921 -204
rect 217949 -232 217983 -204
rect 218011 -232 233157 -204
rect 233185 -232 233219 -204
rect 233247 -232 233281 -204
rect 233309 -232 233343 -204
rect 233371 -232 248517 -204
rect 248545 -232 248579 -204
rect 248607 -232 248641 -204
rect 248669 -232 248703 -204
rect 248731 -232 263877 -204
rect 263905 -232 263939 -204
rect 263967 -232 264001 -204
rect 264029 -232 264063 -204
rect 264091 -232 279237 -204
rect 279265 -232 279299 -204
rect 279327 -232 279361 -204
rect 279389 -232 279423 -204
rect 279451 -232 294597 -204
rect 294625 -232 294659 -204
rect 294687 -232 294721 -204
rect 294749 -232 294783 -204
rect 294811 -232 298248 -204
rect 298276 -232 298310 -204
rect 298338 -232 298372 -204
rect 298400 -232 298434 -204
rect 298462 -232 298510 -204
rect -478 -266 298510 -232
rect -478 -294 -430 -266
rect -402 -294 -368 -266
rect -340 -294 -306 -266
rect -278 -294 -244 -266
rect -216 -294 2757 -266
rect 2785 -294 2819 -266
rect 2847 -294 2881 -266
rect 2909 -294 2943 -266
rect 2971 -294 18117 -266
rect 18145 -294 18179 -266
rect 18207 -294 18241 -266
rect 18269 -294 18303 -266
rect 18331 -294 33477 -266
rect 33505 -294 33539 -266
rect 33567 -294 33601 -266
rect 33629 -294 33663 -266
rect 33691 -294 48837 -266
rect 48865 -294 48899 -266
rect 48927 -294 48961 -266
rect 48989 -294 49023 -266
rect 49051 -294 64197 -266
rect 64225 -294 64259 -266
rect 64287 -294 64321 -266
rect 64349 -294 64383 -266
rect 64411 -294 79557 -266
rect 79585 -294 79619 -266
rect 79647 -294 79681 -266
rect 79709 -294 79743 -266
rect 79771 -294 94917 -266
rect 94945 -294 94979 -266
rect 95007 -294 95041 -266
rect 95069 -294 95103 -266
rect 95131 -294 110277 -266
rect 110305 -294 110339 -266
rect 110367 -294 110401 -266
rect 110429 -294 110463 -266
rect 110491 -294 125637 -266
rect 125665 -294 125699 -266
rect 125727 -294 125761 -266
rect 125789 -294 125823 -266
rect 125851 -294 140997 -266
rect 141025 -294 141059 -266
rect 141087 -294 141121 -266
rect 141149 -294 141183 -266
rect 141211 -294 156357 -266
rect 156385 -294 156419 -266
rect 156447 -294 156481 -266
rect 156509 -294 156543 -266
rect 156571 -294 171717 -266
rect 171745 -294 171779 -266
rect 171807 -294 171841 -266
rect 171869 -294 171903 -266
rect 171931 -294 187077 -266
rect 187105 -294 187139 -266
rect 187167 -294 187201 -266
rect 187229 -294 187263 -266
rect 187291 -294 202437 -266
rect 202465 -294 202499 -266
rect 202527 -294 202561 -266
rect 202589 -294 202623 -266
rect 202651 -294 217797 -266
rect 217825 -294 217859 -266
rect 217887 -294 217921 -266
rect 217949 -294 217983 -266
rect 218011 -294 233157 -266
rect 233185 -294 233219 -266
rect 233247 -294 233281 -266
rect 233309 -294 233343 -266
rect 233371 -294 248517 -266
rect 248545 -294 248579 -266
rect 248607 -294 248641 -266
rect 248669 -294 248703 -266
rect 248731 -294 263877 -266
rect 263905 -294 263939 -266
rect 263967 -294 264001 -266
rect 264029 -294 264063 -266
rect 264091 -294 279237 -266
rect 279265 -294 279299 -266
rect 279327 -294 279361 -266
rect 279389 -294 279423 -266
rect 279451 -294 294597 -266
rect 294625 -294 294659 -266
rect 294687 -294 294721 -266
rect 294749 -294 294783 -266
rect 294811 -294 298248 -266
rect 298276 -294 298310 -266
rect 298338 -294 298372 -266
rect 298400 -294 298434 -266
rect 298462 -294 298510 -266
rect -478 -342 298510 -294
rect -958 -560 298990 -512
rect -958 -588 -910 -560
rect -882 -588 -848 -560
rect -820 -588 -786 -560
rect -758 -588 -724 -560
rect -696 -588 4617 -560
rect 4645 -588 4679 -560
rect 4707 -588 4741 -560
rect 4769 -588 4803 -560
rect 4831 -588 19977 -560
rect 20005 -588 20039 -560
rect 20067 -588 20101 -560
rect 20129 -588 20163 -560
rect 20191 -588 35337 -560
rect 35365 -588 35399 -560
rect 35427 -588 35461 -560
rect 35489 -588 35523 -560
rect 35551 -588 50697 -560
rect 50725 -588 50759 -560
rect 50787 -588 50821 -560
rect 50849 -588 50883 -560
rect 50911 -588 66057 -560
rect 66085 -588 66119 -560
rect 66147 -588 66181 -560
rect 66209 -588 66243 -560
rect 66271 -588 81417 -560
rect 81445 -588 81479 -560
rect 81507 -588 81541 -560
rect 81569 -588 81603 -560
rect 81631 -588 96777 -560
rect 96805 -588 96839 -560
rect 96867 -588 96901 -560
rect 96929 -588 96963 -560
rect 96991 -588 112137 -560
rect 112165 -588 112199 -560
rect 112227 -588 112261 -560
rect 112289 -588 112323 -560
rect 112351 -588 127497 -560
rect 127525 -588 127559 -560
rect 127587 -588 127621 -560
rect 127649 -588 127683 -560
rect 127711 -588 142857 -560
rect 142885 -588 142919 -560
rect 142947 -588 142981 -560
rect 143009 -588 143043 -560
rect 143071 -588 158217 -560
rect 158245 -588 158279 -560
rect 158307 -588 158341 -560
rect 158369 -588 158403 -560
rect 158431 -588 173577 -560
rect 173605 -588 173639 -560
rect 173667 -588 173701 -560
rect 173729 -588 173763 -560
rect 173791 -588 188937 -560
rect 188965 -588 188999 -560
rect 189027 -588 189061 -560
rect 189089 -588 189123 -560
rect 189151 -588 204297 -560
rect 204325 -588 204359 -560
rect 204387 -588 204421 -560
rect 204449 -588 204483 -560
rect 204511 -588 219657 -560
rect 219685 -588 219719 -560
rect 219747 -588 219781 -560
rect 219809 -588 219843 -560
rect 219871 -588 235017 -560
rect 235045 -588 235079 -560
rect 235107 -588 235141 -560
rect 235169 -588 235203 -560
rect 235231 -588 250377 -560
rect 250405 -588 250439 -560
rect 250467 -588 250501 -560
rect 250529 -588 250563 -560
rect 250591 -588 265737 -560
rect 265765 -588 265799 -560
rect 265827 -588 265861 -560
rect 265889 -588 265923 -560
rect 265951 -588 281097 -560
rect 281125 -588 281159 -560
rect 281187 -588 281221 -560
rect 281249 -588 281283 -560
rect 281311 -588 296457 -560
rect 296485 -588 296519 -560
rect 296547 -588 296581 -560
rect 296609 -588 296643 -560
rect 296671 -588 298728 -560
rect 298756 -588 298790 -560
rect 298818 -588 298852 -560
rect 298880 -588 298914 -560
rect 298942 -588 298990 -560
rect -958 -622 298990 -588
rect -958 -650 -910 -622
rect -882 -650 -848 -622
rect -820 -650 -786 -622
rect -758 -650 -724 -622
rect -696 -650 4617 -622
rect 4645 -650 4679 -622
rect 4707 -650 4741 -622
rect 4769 -650 4803 -622
rect 4831 -650 19977 -622
rect 20005 -650 20039 -622
rect 20067 -650 20101 -622
rect 20129 -650 20163 -622
rect 20191 -650 35337 -622
rect 35365 -650 35399 -622
rect 35427 -650 35461 -622
rect 35489 -650 35523 -622
rect 35551 -650 50697 -622
rect 50725 -650 50759 -622
rect 50787 -650 50821 -622
rect 50849 -650 50883 -622
rect 50911 -650 66057 -622
rect 66085 -650 66119 -622
rect 66147 -650 66181 -622
rect 66209 -650 66243 -622
rect 66271 -650 81417 -622
rect 81445 -650 81479 -622
rect 81507 -650 81541 -622
rect 81569 -650 81603 -622
rect 81631 -650 96777 -622
rect 96805 -650 96839 -622
rect 96867 -650 96901 -622
rect 96929 -650 96963 -622
rect 96991 -650 112137 -622
rect 112165 -650 112199 -622
rect 112227 -650 112261 -622
rect 112289 -650 112323 -622
rect 112351 -650 127497 -622
rect 127525 -650 127559 -622
rect 127587 -650 127621 -622
rect 127649 -650 127683 -622
rect 127711 -650 142857 -622
rect 142885 -650 142919 -622
rect 142947 -650 142981 -622
rect 143009 -650 143043 -622
rect 143071 -650 158217 -622
rect 158245 -650 158279 -622
rect 158307 -650 158341 -622
rect 158369 -650 158403 -622
rect 158431 -650 173577 -622
rect 173605 -650 173639 -622
rect 173667 -650 173701 -622
rect 173729 -650 173763 -622
rect 173791 -650 188937 -622
rect 188965 -650 188999 -622
rect 189027 -650 189061 -622
rect 189089 -650 189123 -622
rect 189151 -650 204297 -622
rect 204325 -650 204359 -622
rect 204387 -650 204421 -622
rect 204449 -650 204483 -622
rect 204511 -650 219657 -622
rect 219685 -650 219719 -622
rect 219747 -650 219781 -622
rect 219809 -650 219843 -622
rect 219871 -650 235017 -622
rect 235045 -650 235079 -622
rect 235107 -650 235141 -622
rect 235169 -650 235203 -622
rect 235231 -650 250377 -622
rect 250405 -650 250439 -622
rect 250467 -650 250501 -622
rect 250529 -650 250563 -622
rect 250591 -650 265737 -622
rect 265765 -650 265799 -622
rect 265827 -650 265861 -622
rect 265889 -650 265923 -622
rect 265951 -650 281097 -622
rect 281125 -650 281159 -622
rect 281187 -650 281221 -622
rect 281249 -650 281283 -622
rect 281311 -650 296457 -622
rect 296485 -650 296519 -622
rect 296547 -650 296581 -622
rect 296609 -650 296643 -622
rect 296671 -650 298728 -622
rect 298756 -650 298790 -622
rect 298818 -650 298852 -622
rect 298880 -650 298914 -622
rect 298942 -650 298990 -622
rect -958 -684 298990 -650
rect -958 -712 -910 -684
rect -882 -712 -848 -684
rect -820 -712 -786 -684
rect -758 -712 -724 -684
rect -696 -712 4617 -684
rect 4645 -712 4679 -684
rect 4707 -712 4741 -684
rect 4769 -712 4803 -684
rect 4831 -712 19977 -684
rect 20005 -712 20039 -684
rect 20067 -712 20101 -684
rect 20129 -712 20163 -684
rect 20191 -712 35337 -684
rect 35365 -712 35399 -684
rect 35427 -712 35461 -684
rect 35489 -712 35523 -684
rect 35551 -712 50697 -684
rect 50725 -712 50759 -684
rect 50787 -712 50821 -684
rect 50849 -712 50883 -684
rect 50911 -712 66057 -684
rect 66085 -712 66119 -684
rect 66147 -712 66181 -684
rect 66209 -712 66243 -684
rect 66271 -712 81417 -684
rect 81445 -712 81479 -684
rect 81507 -712 81541 -684
rect 81569 -712 81603 -684
rect 81631 -712 96777 -684
rect 96805 -712 96839 -684
rect 96867 -712 96901 -684
rect 96929 -712 96963 -684
rect 96991 -712 112137 -684
rect 112165 -712 112199 -684
rect 112227 -712 112261 -684
rect 112289 -712 112323 -684
rect 112351 -712 127497 -684
rect 127525 -712 127559 -684
rect 127587 -712 127621 -684
rect 127649 -712 127683 -684
rect 127711 -712 142857 -684
rect 142885 -712 142919 -684
rect 142947 -712 142981 -684
rect 143009 -712 143043 -684
rect 143071 -712 158217 -684
rect 158245 -712 158279 -684
rect 158307 -712 158341 -684
rect 158369 -712 158403 -684
rect 158431 -712 173577 -684
rect 173605 -712 173639 -684
rect 173667 -712 173701 -684
rect 173729 -712 173763 -684
rect 173791 -712 188937 -684
rect 188965 -712 188999 -684
rect 189027 -712 189061 -684
rect 189089 -712 189123 -684
rect 189151 -712 204297 -684
rect 204325 -712 204359 -684
rect 204387 -712 204421 -684
rect 204449 -712 204483 -684
rect 204511 -712 219657 -684
rect 219685 -712 219719 -684
rect 219747 -712 219781 -684
rect 219809 -712 219843 -684
rect 219871 -712 235017 -684
rect 235045 -712 235079 -684
rect 235107 -712 235141 -684
rect 235169 -712 235203 -684
rect 235231 -712 250377 -684
rect 250405 -712 250439 -684
rect 250467 -712 250501 -684
rect 250529 -712 250563 -684
rect 250591 -712 265737 -684
rect 265765 -712 265799 -684
rect 265827 -712 265861 -684
rect 265889 -712 265923 -684
rect 265951 -712 281097 -684
rect 281125 -712 281159 -684
rect 281187 -712 281221 -684
rect 281249 -712 281283 -684
rect 281311 -712 296457 -684
rect 296485 -712 296519 -684
rect 296547 -712 296581 -684
rect 296609 -712 296643 -684
rect 296671 -712 298728 -684
rect 298756 -712 298790 -684
rect 298818 -712 298852 -684
rect 298880 -712 298914 -684
rect 298942 -712 298990 -684
rect -958 -746 298990 -712
rect -958 -774 -910 -746
rect -882 -774 -848 -746
rect -820 -774 -786 -746
rect -758 -774 -724 -746
rect -696 -774 4617 -746
rect 4645 -774 4679 -746
rect 4707 -774 4741 -746
rect 4769 -774 4803 -746
rect 4831 -774 19977 -746
rect 20005 -774 20039 -746
rect 20067 -774 20101 -746
rect 20129 -774 20163 -746
rect 20191 -774 35337 -746
rect 35365 -774 35399 -746
rect 35427 -774 35461 -746
rect 35489 -774 35523 -746
rect 35551 -774 50697 -746
rect 50725 -774 50759 -746
rect 50787 -774 50821 -746
rect 50849 -774 50883 -746
rect 50911 -774 66057 -746
rect 66085 -774 66119 -746
rect 66147 -774 66181 -746
rect 66209 -774 66243 -746
rect 66271 -774 81417 -746
rect 81445 -774 81479 -746
rect 81507 -774 81541 -746
rect 81569 -774 81603 -746
rect 81631 -774 96777 -746
rect 96805 -774 96839 -746
rect 96867 -774 96901 -746
rect 96929 -774 96963 -746
rect 96991 -774 112137 -746
rect 112165 -774 112199 -746
rect 112227 -774 112261 -746
rect 112289 -774 112323 -746
rect 112351 -774 127497 -746
rect 127525 -774 127559 -746
rect 127587 -774 127621 -746
rect 127649 -774 127683 -746
rect 127711 -774 142857 -746
rect 142885 -774 142919 -746
rect 142947 -774 142981 -746
rect 143009 -774 143043 -746
rect 143071 -774 158217 -746
rect 158245 -774 158279 -746
rect 158307 -774 158341 -746
rect 158369 -774 158403 -746
rect 158431 -774 173577 -746
rect 173605 -774 173639 -746
rect 173667 -774 173701 -746
rect 173729 -774 173763 -746
rect 173791 -774 188937 -746
rect 188965 -774 188999 -746
rect 189027 -774 189061 -746
rect 189089 -774 189123 -746
rect 189151 -774 204297 -746
rect 204325 -774 204359 -746
rect 204387 -774 204421 -746
rect 204449 -774 204483 -746
rect 204511 -774 219657 -746
rect 219685 -774 219719 -746
rect 219747 -774 219781 -746
rect 219809 -774 219843 -746
rect 219871 -774 235017 -746
rect 235045 -774 235079 -746
rect 235107 -774 235141 -746
rect 235169 -774 235203 -746
rect 235231 -774 250377 -746
rect 250405 -774 250439 -746
rect 250467 -774 250501 -746
rect 250529 -774 250563 -746
rect 250591 -774 265737 -746
rect 265765 -774 265799 -746
rect 265827 -774 265861 -746
rect 265889 -774 265923 -746
rect 265951 -774 281097 -746
rect 281125 -774 281159 -746
rect 281187 -774 281221 -746
rect 281249 -774 281283 -746
rect 281311 -774 296457 -746
rect 296485 -774 296519 -746
rect 296547 -774 296581 -746
rect 296609 -774 296643 -746
rect 296671 -774 298728 -746
rect 298756 -774 298790 -746
rect 298818 -774 298852 -746
rect 298880 -774 298914 -746
rect 298942 -774 298990 -746
rect -958 -822 298990 -774
use user_proj_example  mprj
timestamp 0
transform 1 0 6000 0 1 1500
box 0 0 280000 174078
<< labels >>
flabel metal3 s 297780 3556 298500 3668 0 FreeSans 448 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 297780 201796 298500 201908 0 FreeSans 448 0 0 0 io_in[10]
port 1 nsew signal input
flabel metal3 s 297780 221620 298500 221732 0 FreeSans 448 0 0 0 io_in[11]
port 2 nsew signal input
flabel metal3 s 297780 241444 298500 241556 0 FreeSans 448 0 0 0 io_in[12]
port 3 nsew signal input
flabel metal3 s 297780 261268 298500 261380 0 FreeSans 448 0 0 0 io_in[13]
port 4 nsew signal input
flabel metal3 s 297780 281092 298500 281204 0 FreeSans 448 0 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 292348 297780 292460 298500 0 FreeSans 448 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 259252 297780 259364 298500 0 FreeSans 448 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 226156 297780 226268 298500 0 FreeSans 448 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 193060 297780 193172 298500 0 FreeSans 448 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 159964 297780 160076 298500 0 FreeSans 448 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 297780 23380 298500 23492 0 FreeSans 448 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 126868 297780 126980 298500 0 FreeSans 448 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 93772 297780 93884 298500 0 FreeSans 448 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 60676 297780 60788 298500 0 FreeSans 448 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 27580 297780 27692 298500 0 FreeSans 448 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s -480 293580 240 293692 0 FreeSans 448 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal3 s -480 272412 240 272524 0 FreeSans 448 0 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s -480 251244 240 251356 0 FreeSans 448 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s -480 230076 240 230188 0 FreeSans 448 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s -480 208908 240 209020 0 FreeSans 448 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal3 s -480 187740 240 187852 0 FreeSans 448 0 0 0 io_in[29]
port 21 nsew signal input
flabel metal3 s 297780 43204 298500 43316 0 FreeSans 448 0 0 0 io_in[2]
port 22 nsew signal input
flabel metal3 s -480 166572 240 166684 0 FreeSans 448 0 0 0 io_in[30]
port 23 nsew signal input
flabel metal3 s -480 145404 240 145516 0 FreeSans 448 0 0 0 io_in[31]
port 24 nsew signal input
flabel metal3 s -480 124236 240 124348 0 FreeSans 448 0 0 0 io_in[32]
port 25 nsew signal input
flabel metal3 s -480 103068 240 103180 0 FreeSans 448 0 0 0 io_in[33]
port 26 nsew signal input
flabel metal3 s -480 81900 240 82012 0 FreeSans 448 0 0 0 io_in[34]
port 27 nsew signal input
flabel metal3 s -480 60732 240 60844 0 FreeSans 448 0 0 0 io_in[35]
port 28 nsew signal input
flabel metal3 s -480 39564 240 39676 0 FreeSans 448 0 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s -480 18396 240 18508 0 FreeSans 448 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 297780 63028 298500 63140 0 FreeSans 448 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal3 s 297780 82852 298500 82964 0 FreeSans 448 0 0 0 io_in[4]
port 32 nsew signal input
flabel metal3 s 297780 102676 298500 102788 0 FreeSans 448 0 0 0 io_in[5]
port 33 nsew signal input
flabel metal3 s 297780 122500 298500 122612 0 FreeSans 448 0 0 0 io_in[6]
port 34 nsew signal input
flabel metal3 s 297780 142324 298500 142436 0 FreeSans 448 0 0 0 io_in[7]
port 35 nsew signal input
flabel metal3 s 297780 162148 298500 162260 0 FreeSans 448 0 0 0 io_in[8]
port 36 nsew signal input
flabel metal3 s 297780 181972 298500 182084 0 FreeSans 448 0 0 0 io_in[9]
port 37 nsew signal input
flabel metal3 s 297780 16772 298500 16884 0 FreeSans 448 0 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal3 s 297780 215012 298500 215124 0 FreeSans 448 0 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal3 s 297780 234836 298500 234948 0 FreeSans 448 0 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal3 s 297780 254660 298500 254772 0 FreeSans 448 0 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal3 s 297780 274484 298500 274596 0 FreeSans 448 0 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal3 s 297780 294308 298500 294420 0 FreeSans 448 0 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 270284 297780 270396 298500 0 FreeSans 448 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 237188 297780 237300 298500 0 FreeSans 448 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 204092 297780 204204 298500 0 FreeSans 448 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 170996 297780 171108 298500 0 FreeSans 448 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 137900 297780 138012 298500 0 FreeSans 448 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal3 s 297780 36596 298500 36708 0 FreeSans 448 0 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 104804 297780 104916 298500 0 FreeSans 448 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 71708 297780 71820 298500 0 FreeSans 448 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 38612 297780 38724 298500 0 FreeSans 448 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 5516 297780 5628 298500 0 FreeSans 448 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal3 s -480 279468 240 279580 0 FreeSans 448 0 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal3 s -480 258300 240 258412 0 FreeSans 448 0 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal3 s -480 237132 240 237244 0 FreeSans 448 0 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal3 s -480 215964 240 216076 0 FreeSans 448 0 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal3 s -480 194796 240 194908 0 FreeSans 448 0 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal3 s -480 173628 240 173740 0 FreeSans 448 0 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal3 s 297780 56420 298500 56532 0 FreeSans 448 0 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal3 s -480 152460 240 152572 0 FreeSans 448 0 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal3 s -480 131292 240 131404 0 FreeSans 448 0 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal3 s -480 110124 240 110236 0 FreeSans 448 0 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal3 s -480 88956 240 89068 0 FreeSans 448 0 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal3 s -480 67788 240 67900 0 FreeSans 448 0 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal3 s -480 46620 240 46732 0 FreeSans 448 0 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal3 s -480 25452 240 25564 0 FreeSans 448 0 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal3 s -480 4284 240 4396 0 FreeSans 448 0 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal3 s 297780 76244 298500 76356 0 FreeSans 448 0 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal3 s 297780 96068 298500 96180 0 FreeSans 448 0 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal3 s 297780 115892 298500 116004 0 FreeSans 448 0 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal3 s 297780 135716 298500 135828 0 FreeSans 448 0 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal3 s 297780 155540 298500 155652 0 FreeSans 448 0 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal3 s 297780 175364 298500 175476 0 FreeSans 448 0 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal3 s 297780 195188 298500 195300 0 FreeSans 448 0 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal3 s 297780 10164 298500 10276 0 FreeSans 448 0 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal3 s 297780 208404 298500 208516 0 FreeSans 448 0 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal3 s 297780 228228 298500 228340 0 FreeSans 448 0 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal3 s 297780 248052 298500 248164 0 FreeSans 448 0 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal3 s 297780 267876 298500 267988 0 FreeSans 448 0 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal3 s 297780 287700 298500 287812 0 FreeSans 448 0 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 281316 297780 281428 298500 0 FreeSans 448 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 248220 297780 248332 298500 0 FreeSans 448 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 215124 297780 215236 298500 0 FreeSans 448 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 182028 297780 182140 298500 0 FreeSans 448 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 148932 297780 149044 298500 0 FreeSans 448 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal3 s 297780 29988 298500 30100 0 FreeSans 448 0 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 115836 297780 115948 298500 0 FreeSans 448 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 82740 297780 82852 298500 0 FreeSans 448 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 49644 297780 49756 298500 0 FreeSans 448 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 16548 297780 16660 298500 0 FreeSans 448 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal3 s -480 286524 240 286636 0 FreeSans 448 0 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal3 s -480 265356 240 265468 0 FreeSans 448 0 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal3 s -480 244188 240 244300 0 FreeSans 448 0 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal3 s -480 223020 240 223132 0 FreeSans 448 0 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal3 s -480 201852 240 201964 0 FreeSans 448 0 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal3 s -480 180684 240 180796 0 FreeSans 448 0 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal3 s 297780 49812 298500 49924 0 FreeSans 448 0 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal3 s -480 159516 240 159628 0 FreeSans 448 0 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal3 s -480 138348 240 138460 0 FreeSans 448 0 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal3 s -480 117180 240 117292 0 FreeSans 448 0 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal3 s -480 96012 240 96124 0 FreeSans 448 0 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal3 s -480 74844 240 74956 0 FreeSans 448 0 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal3 s -480 53676 240 53788 0 FreeSans 448 0 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal3 s -480 32508 240 32620 0 FreeSans 448 0 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal3 s -480 11340 240 11452 0 FreeSans 448 0 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal3 s 297780 69636 298500 69748 0 FreeSans 448 0 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal3 s 297780 89460 298500 89572 0 FreeSans 448 0 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal3 s 297780 109284 298500 109396 0 FreeSans 448 0 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal3 s 297780 129108 298500 129220 0 FreeSans 448 0 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal3 s 297780 148932 298500 149044 0 FreeSans 448 0 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal3 s 297780 168756 298500 168868 0 FreeSans 448 0 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal3 s 297780 188580 298500 188692 0 FreeSans 448 0 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal2 s 106596 -480 106708 240 0 FreeSans 448 90 0 0 la_data_in[0]
port 114 nsew signal input
flabel metal2 s 135156 -480 135268 240 0 FreeSans 448 90 0 0 la_data_in[10]
port 115 nsew signal input
flabel metal2 s 138012 -480 138124 240 0 FreeSans 448 90 0 0 la_data_in[11]
port 116 nsew signal input
flabel metal2 s 140868 -480 140980 240 0 FreeSans 448 90 0 0 la_data_in[12]
port 117 nsew signal input
flabel metal2 s 143724 -480 143836 240 0 FreeSans 448 90 0 0 la_data_in[13]
port 118 nsew signal input
flabel metal2 s 146580 -480 146692 240 0 FreeSans 448 90 0 0 la_data_in[14]
port 119 nsew signal input
flabel metal2 s 149436 -480 149548 240 0 FreeSans 448 90 0 0 la_data_in[15]
port 120 nsew signal input
flabel metal2 s 152292 -480 152404 240 0 FreeSans 448 90 0 0 la_data_in[16]
port 121 nsew signal input
flabel metal2 s 155148 -480 155260 240 0 FreeSans 448 90 0 0 la_data_in[17]
port 122 nsew signal input
flabel metal2 s 158004 -480 158116 240 0 FreeSans 448 90 0 0 la_data_in[18]
port 123 nsew signal input
flabel metal2 s 160860 -480 160972 240 0 FreeSans 448 90 0 0 la_data_in[19]
port 124 nsew signal input
flabel metal2 s 109452 -480 109564 240 0 FreeSans 448 90 0 0 la_data_in[1]
port 125 nsew signal input
flabel metal2 s 163716 -480 163828 240 0 FreeSans 448 90 0 0 la_data_in[20]
port 126 nsew signal input
flabel metal2 s 166572 -480 166684 240 0 FreeSans 448 90 0 0 la_data_in[21]
port 127 nsew signal input
flabel metal2 s 169428 -480 169540 240 0 FreeSans 448 90 0 0 la_data_in[22]
port 128 nsew signal input
flabel metal2 s 172284 -480 172396 240 0 FreeSans 448 90 0 0 la_data_in[23]
port 129 nsew signal input
flabel metal2 s 175140 -480 175252 240 0 FreeSans 448 90 0 0 la_data_in[24]
port 130 nsew signal input
flabel metal2 s 177996 -480 178108 240 0 FreeSans 448 90 0 0 la_data_in[25]
port 131 nsew signal input
flabel metal2 s 180852 -480 180964 240 0 FreeSans 448 90 0 0 la_data_in[26]
port 132 nsew signal input
flabel metal2 s 183708 -480 183820 240 0 FreeSans 448 90 0 0 la_data_in[27]
port 133 nsew signal input
flabel metal2 s 186564 -480 186676 240 0 FreeSans 448 90 0 0 la_data_in[28]
port 134 nsew signal input
flabel metal2 s 189420 -480 189532 240 0 FreeSans 448 90 0 0 la_data_in[29]
port 135 nsew signal input
flabel metal2 s 112308 -480 112420 240 0 FreeSans 448 90 0 0 la_data_in[2]
port 136 nsew signal input
flabel metal2 s 192276 -480 192388 240 0 FreeSans 448 90 0 0 la_data_in[30]
port 137 nsew signal input
flabel metal2 s 195132 -480 195244 240 0 FreeSans 448 90 0 0 la_data_in[31]
port 138 nsew signal input
flabel metal2 s 197988 -480 198100 240 0 FreeSans 448 90 0 0 la_data_in[32]
port 139 nsew signal input
flabel metal2 s 200844 -480 200956 240 0 FreeSans 448 90 0 0 la_data_in[33]
port 140 nsew signal input
flabel metal2 s 203700 -480 203812 240 0 FreeSans 448 90 0 0 la_data_in[34]
port 141 nsew signal input
flabel metal2 s 206556 -480 206668 240 0 FreeSans 448 90 0 0 la_data_in[35]
port 142 nsew signal input
flabel metal2 s 209412 -480 209524 240 0 FreeSans 448 90 0 0 la_data_in[36]
port 143 nsew signal input
flabel metal2 s 212268 -480 212380 240 0 FreeSans 448 90 0 0 la_data_in[37]
port 144 nsew signal input
flabel metal2 s 215124 -480 215236 240 0 FreeSans 448 90 0 0 la_data_in[38]
port 145 nsew signal input
flabel metal2 s 217980 -480 218092 240 0 FreeSans 448 90 0 0 la_data_in[39]
port 146 nsew signal input
flabel metal2 s 115164 -480 115276 240 0 FreeSans 448 90 0 0 la_data_in[3]
port 147 nsew signal input
flabel metal2 s 220836 -480 220948 240 0 FreeSans 448 90 0 0 la_data_in[40]
port 148 nsew signal input
flabel metal2 s 223692 -480 223804 240 0 FreeSans 448 90 0 0 la_data_in[41]
port 149 nsew signal input
flabel metal2 s 226548 -480 226660 240 0 FreeSans 448 90 0 0 la_data_in[42]
port 150 nsew signal input
flabel metal2 s 229404 -480 229516 240 0 FreeSans 448 90 0 0 la_data_in[43]
port 151 nsew signal input
flabel metal2 s 232260 -480 232372 240 0 FreeSans 448 90 0 0 la_data_in[44]
port 152 nsew signal input
flabel metal2 s 235116 -480 235228 240 0 FreeSans 448 90 0 0 la_data_in[45]
port 153 nsew signal input
flabel metal2 s 237972 -480 238084 240 0 FreeSans 448 90 0 0 la_data_in[46]
port 154 nsew signal input
flabel metal2 s 240828 -480 240940 240 0 FreeSans 448 90 0 0 la_data_in[47]
port 155 nsew signal input
flabel metal2 s 243684 -480 243796 240 0 FreeSans 448 90 0 0 la_data_in[48]
port 156 nsew signal input
flabel metal2 s 246540 -480 246652 240 0 FreeSans 448 90 0 0 la_data_in[49]
port 157 nsew signal input
flabel metal2 s 118020 -480 118132 240 0 FreeSans 448 90 0 0 la_data_in[4]
port 158 nsew signal input
flabel metal2 s 249396 -480 249508 240 0 FreeSans 448 90 0 0 la_data_in[50]
port 159 nsew signal input
flabel metal2 s 252252 -480 252364 240 0 FreeSans 448 90 0 0 la_data_in[51]
port 160 nsew signal input
flabel metal2 s 255108 -480 255220 240 0 FreeSans 448 90 0 0 la_data_in[52]
port 161 nsew signal input
flabel metal2 s 257964 -480 258076 240 0 FreeSans 448 90 0 0 la_data_in[53]
port 162 nsew signal input
flabel metal2 s 260820 -480 260932 240 0 FreeSans 448 90 0 0 la_data_in[54]
port 163 nsew signal input
flabel metal2 s 263676 -480 263788 240 0 FreeSans 448 90 0 0 la_data_in[55]
port 164 nsew signal input
flabel metal2 s 266532 -480 266644 240 0 FreeSans 448 90 0 0 la_data_in[56]
port 165 nsew signal input
flabel metal2 s 269388 -480 269500 240 0 FreeSans 448 90 0 0 la_data_in[57]
port 166 nsew signal input
flabel metal2 s 272244 -480 272356 240 0 FreeSans 448 90 0 0 la_data_in[58]
port 167 nsew signal input
flabel metal2 s 275100 -480 275212 240 0 FreeSans 448 90 0 0 la_data_in[59]
port 168 nsew signal input
flabel metal2 s 120876 -480 120988 240 0 FreeSans 448 90 0 0 la_data_in[5]
port 169 nsew signal input
flabel metal2 s 277956 -480 278068 240 0 FreeSans 448 90 0 0 la_data_in[60]
port 170 nsew signal input
flabel metal2 s 280812 -480 280924 240 0 FreeSans 448 90 0 0 la_data_in[61]
port 171 nsew signal input
flabel metal2 s 283668 -480 283780 240 0 FreeSans 448 90 0 0 la_data_in[62]
port 172 nsew signal input
flabel metal2 s 286524 -480 286636 240 0 FreeSans 448 90 0 0 la_data_in[63]
port 173 nsew signal input
flabel metal2 s 123732 -480 123844 240 0 FreeSans 448 90 0 0 la_data_in[6]
port 174 nsew signal input
flabel metal2 s 126588 -480 126700 240 0 FreeSans 448 90 0 0 la_data_in[7]
port 175 nsew signal input
flabel metal2 s 129444 -480 129556 240 0 FreeSans 448 90 0 0 la_data_in[8]
port 176 nsew signal input
flabel metal2 s 132300 -480 132412 240 0 FreeSans 448 90 0 0 la_data_in[9]
port 177 nsew signal input
flabel metal2 s 107548 -480 107660 240 0 FreeSans 448 90 0 0 la_data_out[0]
port 178 nsew signal tristate
flabel metal2 s 136108 -480 136220 240 0 FreeSans 448 90 0 0 la_data_out[10]
port 179 nsew signal tristate
flabel metal2 s 138964 -480 139076 240 0 FreeSans 448 90 0 0 la_data_out[11]
port 180 nsew signal tristate
flabel metal2 s 141820 -480 141932 240 0 FreeSans 448 90 0 0 la_data_out[12]
port 181 nsew signal tristate
flabel metal2 s 144676 -480 144788 240 0 FreeSans 448 90 0 0 la_data_out[13]
port 182 nsew signal tristate
flabel metal2 s 147532 -480 147644 240 0 FreeSans 448 90 0 0 la_data_out[14]
port 183 nsew signal tristate
flabel metal2 s 150388 -480 150500 240 0 FreeSans 448 90 0 0 la_data_out[15]
port 184 nsew signal tristate
flabel metal2 s 153244 -480 153356 240 0 FreeSans 448 90 0 0 la_data_out[16]
port 185 nsew signal tristate
flabel metal2 s 156100 -480 156212 240 0 FreeSans 448 90 0 0 la_data_out[17]
port 186 nsew signal tristate
flabel metal2 s 158956 -480 159068 240 0 FreeSans 448 90 0 0 la_data_out[18]
port 187 nsew signal tristate
flabel metal2 s 161812 -480 161924 240 0 FreeSans 448 90 0 0 la_data_out[19]
port 188 nsew signal tristate
flabel metal2 s 110404 -480 110516 240 0 FreeSans 448 90 0 0 la_data_out[1]
port 189 nsew signal tristate
flabel metal2 s 164668 -480 164780 240 0 FreeSans 448 90 0 0 la_data_out[20]
port 190 nsew signal tristate
flabel metal2 s 167524 -480 167636 240 0 FreeSans 448 90 0 0 la_data_out[21]
port 191 nsew signal tristate
flabel metal2 s 170380 -480 170492 240 0 FreeSans 448 90 0 0 la_data_out[22]
port 192 nsew signal tristate
flabel metal2 s 173236 -480 173348 240 0 FreeSans 448 90 0 0 la_data_out[23]
port 193 nsew signal tristate
flabel metal2 s 176092 -480 176204 240 0 FreeSans 448 90 0 0 la_data_out[24]
port 194 nsew signal tristate
flabel metal2 s 178948 -480 179060 240 0 FreeSans 448 90 0 0 la_data_out[25]
port 195 nsew signal tristate
flabel metal2 s 181804 -480 181916 240 0 FreeSans 448 90 0 0 la_data_out[26]
port 196 nsew signal tristate
flabel metal2 s 184660 -480 184772 240 0 FreeSans 448 90 0 0 la_data_out[27]
port 197 nsew signal tristate
flabel metal2 s 187516 -480 187628 240 0 FreeSans 448 90 0 0 la_data_out[28]
port 198 nsew signal tristate
flabel metal2 s 190372 -480 190484 240 0 FreeSans 448 90 0 0 la_data_out[29]
port 199 nsew signal tristate
flabel metal2 s 113260 -480 113372 240 0 FreeSans 448 90 0 0 la_data_out[2]
port 200 nsew signal tristate
flabel metal2 s 193228 -480 193340 240 0 FreeSans 448 90 0 0 la_data_out[30]
port 201 nsew signal tristate
flabel metal2 s 196084 -480 196196 240 0 FreeSans 448 90 0 0 la_data_out[31]
port 202 nsew signal tristate
flabel metal2 s 198940 -480 199052 240 0 FreeSans 448 90 0 0 la_data_out[32]
port 203 nsew signal tristate
flabel metal2 s 201796 -480 201908 240 0 FreeSans 448 90 0 0 la_data_out[33]
port 204 nsew signal tristate
flabel metal2 s 204652 -480 204764 240 0 FreeSans 448 90 0 0 la_data_out[34]
port 205 nsew signal tristate
flabel metal2 s 207508 -480 207620 240 0 FreeSans 448 90 0 0 la_data_out[35]
port 206 nsew signal tristate
flabel metal2 s 210364 -480 210476 240 0 FreeSans 448 90 0 0 la_data_out[36]
port 207 nsew signal tristate
flabel metal2 s 213220 -480 213332 240 0 FreeSans 448 90 0 0 la_data_out[37]
port 208 nsew signal tristate
flabel metal2 s 216076 -480 216188 240 0 FreeSans 448 90 0 0 la_data_out[38]
port 209 nsew signal tristate
flabel metal2 s 218932 -480 219044 240 0 FreeSans 448 90 0 0 la_data_out[39]
port 210 nsew signal tristate
flabel metal2 s 116116 -480 116228 240 0 FreeSans 448 90 0 0 la_data_out[3]
port 211 nsew signal tristate
flabel metal2 s 221788 -480 221900 240 0 FreeSans 448 90 0 0 la_data_out[40]
port 212 nsew signal tristate
flabel metal2 s 224644 -480 224756 240 0 FreeSans 448 90 0 0 la_data_out[41]
port 213 nsew signal tristate
flabel metal2 s 227500 -480 227612 240 0 FreeSans 448 90 0 0 la_data_out[42]
port 214 nsew signal tristate
flabel metal2 s 230356 -480 230468 240 0 FreeSans 448 90 0 0 la_data_out[43]
port 215 nsew signal tristate
flabel metal2 s 233212 -480 233324 240 0 FreeSans 448 90 0 0 la_data_out[44]
port 216 nsew signal tristate
flabel metal2 s 236068 -480 236180 240 0 FreeSans 448 90 0 0 la_data_out[45]
port 217 nsew signal tristate
flabel metal2 s 238924 -480 239036 240 0 FreeSans 448 90 0 0 la_data_out[46]
port 218 nsew signal tristate
flabel metal2 s 241780 -480 241892 240 0 FreeSans 448 90 0 0 la_data_out[47]
port 219 nsew signal tristate
flabel metal2 s 244636 -480 244748 240 0 FreeSans 448 90 0 0 la_data_out[48]
port 220 nsew signal tristate
flabel metal2 s 247492 -480 247604 240 0 FreeSans 448 90 0 0 la_data_out[49]
port 221 nsew signal tristate
flabel metal2 s 118972 -480 119084 240 0 FreeSans 448 90 0 0 la_data_out[4]
port 222 nsew signal tristate
flabel metal2 s 250348 -480 250460 240 0 FreeSans 448 90 0 0 la_data_out[50]
port 223 nsew signal tristate
flabel metal2 s 253204 -480 253316 240 0 FreeSans 448 90 0 0 la_data_out[51]
port 224 nsew signal tristate
flabel metal2 s 256060 -480 256172 240 0 FreeSans 448 90 0 0 la_data_out[52]
port 225 nsew signal tristate
flabel metal2 s 258916 -480 259028 240 0 FreeSans 448 90 0 0 la_data_out[53]
port 226 nsew signal tristate
flabel metal2 s 261772 -480 261884 240 0 FreeSans 448 90 0 0 la_data_out[54]
port 227 nsew signal tristate
flabel metal2 s 264628 -480 264740 240 0 FreeSans 448 90 0 0 la_data_out[55]
port 228 nsew signal tristate
flabel metal2 s 267484 -480 267596 240 0 FreeSans 448 90 0 0 la_data_out[56]
port 229 nsew signal tristate
flabel metal2 s 270340 -480 270452 240 0 FreeSans 448 90 0 0 la_data_out[57]
port 230 nsew signal tristate
flabel metal2 s 273196 -480 273308 240 0 FreeSans 448 90 0 0 la_data_out[58]
port 231 nsew signal tristate
flabel metal2 s 276052 -480 276164 240 0 FreeSans 448 90 0 0 la_data_out[59]
port 232 nsew signal tristate
flabel metal2 s 121828 -480 121940 240 0 FreeSans 448 90 0 0 la_data_out[5]
port 233 nsew signal tristate
flabel metal2 s 278908 -480 279020 240 0 FreeSans 448 90 0 0 la_data_out[60]
port 234 nsew signal tristate
flabel metal2 s 281764 -480 281876 240 0 FreeSans 448 90 0 0 la_data_out[61]
port 235 nsew signal tristate
flabel metal2 s 284620 -480 284732 240 0 FreeSans 448 90 0 0 la_data_out[62]
port 236 nsew signal tristate
flabel metal2 s 287476 -480 287588 240 0 FreeSans 448 90 0 0 la_data_out[63]
port 237 nsew signal tristate
flabel metal2 s 124684 -480 124796 240 0 FreeSans 448 90 0 0 la_data_out[6]
port 238 nsew signal tristate
flabel metal2 s 127540 -480 127652 240 0 FreeSans 448 90 0 0 la_data_out[7]
port 239 nsew signal tristate
flabel metal2 s 130396 -480 130508 240 0 FreeSans 448 90 0 0 la_data_out[8]
port 240 nsew signal tristate
flabel metal2 s 133252 -480 133364 240 0 FreeSans 448 90 0 0 la_data_out[9]
port 241 nsew signal tristate
flabel metal2 s 108500 -480 108612 240 0 FreeSans 448 90 0 0 la_oenb[0]
port 242 nsew signal input
flabel metal2 s 137060 -480 137172 240 0 FreeSans 448 90 0 0 la_oenb[10]
port 243 nsew signal input
flabel metal2 s 139916 -480 140028 240 0 FreeSans 448 90 0 0 la_oenb[11]
port 244 nsew signal input
flabel metal2 s 142772 -480 142884 240 0 FreeSans 448 90 0 0 la_oenb[12]
port 245 nsew signal input
flabel metal2 s 145628 -480 145740 240 0 FreeSans 448 90 0 0 la_oenb[13]
port 246 nsew signal input
flabel metal2 s 148484 -480 148596 240 0 FreeSans 448 90 0 0 la_oenb[14]
port 247 nsew signal input
flabel metal2 s 151340 -480 151452 240 0 FreeSans 448 90 0 0 la_oenb[15]
port 248 nsew signal input
flabel metal2 s 154196 -480 154308 240 0 FreeSans 448 90 0 0 la_oenb[16]
port 249 nsew signal input
flabel metal2 s 157052 -480 157164 240 0 FreeSans 448 90 0 0 la_oenb[17]
port 250 nsew signal input
flabel metal2 s 159908 -480 160020 240 0 FreeSans 448 90 0 0 la_oenb[18]
port 251 nsew signal input
flabel metal2 s 162764 -480 162876 240 0 FreeSans 448 90 0 0 la_oenb[19]
port 252 nsew signal input
flabel metal2 s 111356 -480 111468 240 0 FreeSans 448 90 0 0 la_oenb[1]
port 253 nsew signal input
flabel metal2 s 165620 -480 165732 240 0 FreeSans 448 90 0 0 la_oenb[20]
port 254 nsew signal input
flabel metal2 s 168476 -480 168588 240 0 FreeSans 448 90 0 0 la_oenb[21]
port 255 nsew signal input
flabel metal2 s 171332 -480 171444 240 0 FreeSans 448 90 0 0 la_oenb[22]
port 256 nsew signal input
flabel metal2 s 174188 -480 174300 240 0 FreeSans 448 90 0 0 la_oenb[23]
port 257 nsew signal input
flabel metal2 s 177044 -480 177156 240 0 FreeSans 448 90 0 0 la_oenb[24]
port 258 nsew signal input
flabel metal2 s 179900 -480 180012 240 0 FreeSans 448 90 0 0 la_oenb[25]
port 259 nsew signal input
flabel metal2 s 182756 -480 182868 240 0 FreeSans 448 90 0 0 la_oenb[26]
port 260 nsew signal input
flabel metal2 s 185612 -480 185724 240 0 FreeSans 448 90 0 0 la_oenb[27]
port 261 nsew signal input
flabel metal2 s 188468 -480 188580 240 0 FreeSans 448 90 0 0 la_oenb[28]
port 262 nsew signal input
flabel metal2 s 191324 -480 191436 240 0 FreeSans 448 90 0 0 la_oenb[29]
port 263 nsew signal input
flabel metal2 s 114212 -480 114324 240 0 FreeSans 448 90 0 0 la_oenb[2]
port 264 nsew signal input
flabel metal2 s 194180 -480 194292 240 0 FreeSans 448 90 0 0 la_oenb[30]
port 265 nsew signal input
flabel metal2 s 197036 -480 197148 240 0 FreeSans 448 90 0 0 la_oenb[31]
port 266 nsew signal input
flabel metal2 s 199892 -480 200004 240 0 FreeSans 448 90 0 0 la_oenb[32]
port 267 nsew signal input
flabel metal2 s 202748 -480 202860 240 0 FreeSans 448 90 0 0 la_oenb[33]
port 268 nsew signal input
flabel metal2 s 205604 -480 205716 240 0 FreeSans 448 90 0 0 la_oenb[34]
port 269 nsew signal input
flabel metal2 s 208460 -480 208572 240 0 FreeSans 448 90 0 0 la_oenb[35]
port 270 nsew signal input
flabel metal2 s 211316 -480 211428 240 0 FreeSans 448 90 0 0 la_oenb[36]
port 271 nsew signal input
flabel metal2 s 214172 -480 214284 240 0 FreeSans 448 90 0 0 la_oenb[37]
port 272 nsew signal input
flabel metal2 s 217028 -480 217140 240 0 FreeSans 448 90 0 0 la_oenb[38]
port 273 nsew signal input
flabel metal2 s 219884 -480 219996 240 0 FreeSans 448 90 0 0 la_oenb[39]
port 274 nsew signal input
flabel metal2 s 117068 -480 117180 240 0 FreeSans 448 90 0 0 la_oenb[3]
port 275 nsew signal input
flabel metal2 s 222740 -480 222852 240 0 FreeSans 448 90 0 0 la_oenb[40]
port 276 nsew signal input
flabel metal2 s 225596 -480 225708 240 0 FreeSans 448 90 0 0 la_oenb[41]
port 277 nsew signal input
flabel metal2 s 228452 -480 228564 240 0 FreeSans 448 90 0 0 la_oenb[42]
port 278 nsew signal input
flabel metal2 s 231308 -480 231420 240 0 FreeSans 448 90 0 0 la_oenb[43]
port 279 nsew signal input
flabel metal2 s 234164 -480 234276 240 0 FreeSans 448 90 0 0 la_oenb[44]
port 280 nsew signal input
flabel metal2 s 237020 -480 237132 240 0 FreeSans 448 90 0 0 la_oenb[45]
port 281 nsew signal input
flabel metal2 s 239876 -480 239988 240 0 FreeSans 448 90 0 0 la_oenb[46]
port 282 nsew signal input
flabel metal2 s 242732 -480 242844 240 0 FreeSans 448 90 0 0 la_oenb[47]
port 283 nsew signal input
flabel metal2 s 245588 -480 245700 240 0 FreeSans 448 90 0 0 la_oenb[48]
port 284 nsew signal input
flabel metal2 s 248444 -480 248556 240 0 FreeSans 448 90 0 0 la_oenb[49]
port 285 nsew signal input
flabel metal2 s 119924 -480 120036 240 0 FreeSans 448 90 0 0 la_oenb[4]
port 286 nsew signal input
flabel metal2 s 251300 -480 251412 240 0 FreeSans 448 90 0 0 la_oenb[50]
port 287 nsew signal input
flabel metal2 s 254156 -480 254268 240 0 FreeSans 448 90 0 0 la_oenb[51]
port 288 nsew signal input
flabel metal2 s 257012 -480 257124 240 0 FreeSans 448 90 0 0 la_oenb[52]
port 289 nsew signal input
flabel metal2 s 259868 -480 259980 240 0 FreeSans 448 90 0 0 la_oenb[53]
port 290 nsew signal input
flabel metal2 s 262724 -480 262836 240 0 FreeSans 448 90 0 0 la_oenb[54]
port 291 nsew signal input
flabel metal2 s 265580 -480 265692 240 0 FreeSans 448 90 0 0 la_oenb[55]
port 292 nsew signal input
flabel metal2 s 268436 -480 268548 240 0 FreeSans 448 90 0 0 la_oenb[56]
port 293 nsew signal input
flabel metal2 s 271292 -480 271404 240 0 FreeSans 448 90 0 0 la_oenb[57]
port 294 nsew signal input
flabel metal2 s 274148 -480 274260 240 0 FreeSans 448 90 0 0 la_oenb[58]
port 295 nsew signal input
flabel metal2 s 277004 -480 277116 240 0 FreeSans 448 90 0 0 la_oenb[59]
port 296 nsew signal input
flabel metal2 s 122780 -480 122892 240 0 FreeSans 448 90 0 0 la_oenb[5]
port 297 nsew signal input
flabel metal2 s 279860 -480 279972 240 0 FreeSans 448 90 0 0 la_oenb[60]
port 298 nsew signal input
flabel metal2 s 282716 -480 282828 240 0 FreeSans 448 90 0 0 la_oenb[61]
port 299 nsew signal input
flabel metal2 s 285572 -480 285684 240 0 FreeSans 448 90 0 0 la_oenb[62]
port 300 nsew signal input
flabel metal2 s 288428 -480 288540 240 0 FreeSans 448 90 0 0 la_oenb[63]
port 301 nsew signal input
flabel metal2 s 125636 -480 125748 240 0 FreeSans 448 90 0 0 la_oenb[6]
port 302 nsew signal input
flabel metal2 s 128492 -480 128604 240 0 FreeSans 448 90 0 0 la_oenb[7]
port 303 nsew signal input
flabel metal2 s 131348 -480 131460 240 0 FreeSans 448 90 0 0 la_oenb[8]
port 304 nsew signal input
flabel metal2 s 134204 -480 134316 240 0 FreeSans 448 90 0 0 la_oenb[9]
port 305 nsew signal input
flabel metal2 s 289380 -480 289492 240 0 FreeSans 448 90 0 0 user_clock2
port 306 nsew signal input
flabel metal2 s 290332 -480 290444 240 0 FreeSans 448 90 0 0 user_irq[0]
port 307 nsew signal tristate
flabel metal2 s 291284 -480 291396 240 0 FreeSans 448 90 0 0 user_irq[1]
port 308 nsew signal tristate
flabel metal2 s 292236 -480 292348 240 0 FreeSans 448 90 0 0 user_irq[2]
port 309 nsew signal tristate
flabel metal4 s -478 -342 -168 298654 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -478 -342 298510 -32 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -478 298344 298510 298654 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 298200 -342 298510 298654 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 2709 -822 3019 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 18069 -822 18379 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 33429 -822 33739 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 48789 -822 49099 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 64149 -822 64459 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 79509 -822 79819 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 94869 -822 95179 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 110229 -822 110539 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 125589 -822 125899 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 140949 -822 141259 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 156309 -822 156619 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 171669 -822 171979 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 187029 -822 187339 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 202389 -822 202699 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 217749 -822 218059 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 233109 -822 233419 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 248469 -822 248779 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 263829 -822 264139 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 279189 -822 279499 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 294549 -822 294859 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 1913 298990 2223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 10913 298990 11223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 19913 298990 20223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 28913 298990 29223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 37913 298990 38223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 46913 298990 47223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 55913 298990 56223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 64913 298990 65223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 73913 298990 74223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 82913 298990 83223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 91913 298990 92223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 100913 298990 101223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 109913 298990 110223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 118913 298990 119223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 127913 298990 128223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 136913 298990 137223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 145913 298990 146223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 154913 298990 155223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 163913 298990 164223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 172913 298990 173223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 181913 298990 182223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 190913 298990 191223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 199913 298990 200223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 208913 298990 209223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 217913 298990 218223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 226913 298990 227223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 235913 298990 236223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 244913 298990 245223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 253913 298990 254223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 262913 298990 263223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 271913 298990 272223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 280913 298990 281223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 289913 298990 290223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s -958 -822 -648 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 -822 298990 -512 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 298824 298990 299134 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 298680 -822 298990 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 4569 -822 4879 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 19929 -822 20239 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 35289 -822 35599 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 50649 -822 50959 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 66009 -822 66319 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 81369 -822 81679 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 96729 -822 97039 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 112089 -822 112399 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 127449 -822 127759 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 142809 -822 143119 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 158169 -822 158479 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 173529 -822 173839 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 188889 -822 189199 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 204249 -822 204559 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 219609 -822 219919 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 234969 -822 235279 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 250329 -822 250639 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 265689 -822 265999 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 281049 -822 281359 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 296409 -822 296719 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 4913 298990 5223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 13913 298990 14223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 22913 298990 23223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 31913 298990 32223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 40913 298990 41223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 49913 298990 50223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 58913 298990 59223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 67913 298990 68223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 76913 298990 77223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 85913 298990 86223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 94913 298990 95223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 103913 298990 104223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 112913 298990 113223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 121913 298990 122223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 130913 298990 131223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 139913 298990 140223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 148913 298990 149223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 157913 298990 158223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 166913 298990 167223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 175913 298990 176223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 184913 298990 185223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 193913 298990 194223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 202913 298990 203223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 211913 298990 212223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 220913 298990 221223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 229913 298990 230223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 238913 298990 239223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 247913 298990 248223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 256913 298990 257223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 265913 298990 266223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 274913 298990 275223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 283913 298990 284223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 292913 298990 293223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal2 s 5684 -480 5796 240 0 FreeSans 448 90 0 0 wb_clk_i
port 312 nsew signal input
flabel metal2 s 6636 -480 6748 240 0 FreeSans 448 90 0 0 wb_rst_i
port 313 nsew signal input
flabel metal2 s 7588 -480 7700 240 0 FreeSans 448 90 0 0 wbs_ack_o
port 314 nsew signal tristate
flabel metal2 s 11396 -480 11508 240 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 315 nsew signal input
flabel metal2 s 43764 -480 43876 240 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 316 nsew signal input
flabel metal2 s 46620 -480 46732 240 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 317 nsew signal input
flabel metal2 s 49476 -480 49588 240 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 318 nsew signal input
flabel metal2 s 52332 -480 52444 240 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 319 nsew signal input
flabel metal2 s 55188 -480 55300 240 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 320 nsew signal input
flabel metal2 s 58044 -480 58156 240 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 321 nsew signal input
flabel metal2 s 60900 -480 61012 240 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 322 nsew signal input
flabel metal2 s 63756 -480 63868 240 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 323 nsew signal input
flabel metal2 s 66612 -480 66724 240 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 324 nsew signal input
flabel metal2 s 69468 -480 69580 240 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 325 nsew signal input
flabel metal2 s 15204 -480 15316 240 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 326 nsew signal input
flabel metal2 s 72324 -480 72436 240 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 327 nsew signal input
flabel metal2 s 75180 -480 75292 240 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 328 nsew signal input
flabel metal2 s 78036 -480 78148 240 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 329 nsew signal input
flabel metal2 s 80892 -480 81004 240 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 330 nsew signal input
flabel metal2 s 83748 -480 83860 240 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 331 nsew signal input
flabel metal2 s 86604 -480 86716 240 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 332 nsew signal input
flabel metal2 s 89460 -480 89572 240 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 333 nsew signal input
flabel metal2 s 92316 -480 92428 240 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 334 nsew signal input
flabel metal2 s 95172 -480 95284 240 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 335 nsew signal input
flabel metal2 s 98028 -480 98140 240 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 336 nsew signal input
flabel metal2 s 19012 -480 19124 240 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 337 nsew signal input
flabel metal2 s 100884 -480 100996 240 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 338 nsew signal input
flabel metal2 s 103740 -480 103852 240 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 339 nsew signal input
flabel metal2 s 22820 -480 22932 240 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 340 nsew signal input
flabel metal2 s 26628 -480 26740 240 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 341 nsew signal input
flabel metal2 s 29484 -480 29596 240 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 342 nsew signal input
flabel metal2 s 32340 -480 32452 240 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 343 nsew signal input
flabel metal2 s 35196 -480 35308 240 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 344 nsew signal input
flabel metal2 s 38052 -480 38164 240 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 345 nsew signal input
flabel metal2 s 40908 -480 41020 240 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 346 nsew signal input
flabel metal2 s 8540 -480 8652 240 0 FreeSans 448 90 0 0 wbs_cyc_i
port 347 nsew signal input
flabel metal2 s 12348 -480 12460 240 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 348 nsew signal input
flabel metal2 s 44716 -480 44828 240 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 349 nsew signal input
flabel metal2 s 47572 -480 47684 240 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 350 nsew signal input
flabel metal2 s 50428 -480 50540 240 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 351 nsew signal input
flabel metal2 s 53284 -480 53396 240 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 352 nsew signal input
flabel metal2 s 56140 -480 56252 240 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 353 nsew signal input
flabel metal2 s 58996 -480 59108 240 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 354 nsew signal input
flabel metal2 s 61852 -480 61964 240 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 355 nsew signal input
flabel metal2 s 64708 -480 64820 240 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 356 nsew signal input
flabel metal2 s 67564 -480 67676 240 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 357 nsew signal input
flabel metal2 s 70420 -480 70532 240 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 358 nsew signal input
flabel metal2 s 16156 -480 16268 240 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 359 nsew signal input
flabel metal2 s 73276 -480 73388 240 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 360 nsew signal input
flabel metal2 s 76132 -480 76244 240 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 361 nsew signal input
flabel metal2 s 78988 -480 79100 240 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 362 nsew signal input
flabel metal2 s 81844 -480 81956 240 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 363 nsew signal input
flabel metal2 s 84700 -480 84812 240 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 364 nsew signal input
flabel metal2 s 87556 -480 87668 240 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 365 nsew signal input
flabel metal2 s 90412 -480 90524 240 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 366 nsew signal input
flabel metal2 s 93268 -480 93380 240 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 367 nsew signal input
flabel metal2 s 96124 -480 96236 240 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 368 nsew signal input
flabel metal2 s 98980 -480 99092 240 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 369 nsew signal input
flabel metal2 s 19964 -480 20076 240 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 370 nsew signal input
flabel metal2 s 101836 -480 101948 240 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 371 nsew signal input
flabel metal2 s 104692 -480 104804 240 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 372 nsew signal input
flabel metal2 s 23772 -480 23884 240 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 373 nsew signal input
flabel metal2 s 27580 -480 27692 240 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 374 nsew signal input
flabel metal2 s 30436 -480 30548 240 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 375 nsew signal input
flabel metal2 s 33292 -480 33404 240 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 376 nsew signal input
flabel metal2 s 36148 -480 36260 240 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 377 nsew signal input
flabel metal2 s 39004 -480 39116 240 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 378 nsew signal input
flabel metal2 s 41860 -480 41972 240 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 379 nsew signal input
flabel metal2 s 13300 -480 13412 240 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 380 nsew signal tristate
flabel metal2 s 45668 -480 45780 240 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 381 nsew signal tristate
flabel metal2 s 48524 -480 48636 240 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 382 nsew signal tristate
flabel metal2 s 51380 -480 51492 240 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 383 nsew signal tristate
flabel metal2 s 54236 -480 54348 240 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 384 nsew signal tristate
flabel metal2 s 57092 -480 57204 240 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 385 nsew signal tristate
flabel metal2 s 59948 -480 60060 240 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 386 nsew signal tristate
flabel metal2 s 62804 -480 62916 240 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 387 nsew signal tristate
flabel metal2 s 65660 -480 65772 240 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 388 nsew signal tristate
flabel metal2 s 68516 -480 68628 240 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 389 nsew signal tristate
flabel metal2 s 71372 -480 71484 240 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 390 nsew signal tristate
flabel metal2 s 17108 -480 17220 240 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 391 nsew signal tristate
flabel metal2 s 74228 -480 74340 240 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 392 nsew signal tristate
flabel metal2 s 77084 -480 77196 240 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 393 nsew signal tristate
flabel metal2 s 79940 -480 80052 240 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 394 nsew signal tristate
flabel metal2 s 82796 -480 82908 240 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 395 nsew signal tristate
flabel metal2 s 85652 -480 85764 240 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 396 nsew signal tristate
flabel metal2 s 88508 -480 88620 240 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 397 nsew signal tristate
flabel metal2 s 91364 -480 91476 240 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 398 nsew signal tristate
flabel metal2 s 94220 -480 94332 240 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 399 nsew signal tristate
flabel metal2 s 97076 -480 97188 240 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 400 nsew signal tristate
flabel metal2 s 99932 -480 100044 240 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 401 nsew signal tristate
flabel metal2 s 20916 -480 21028 240 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 402 nsew signal tristate
flabel metal2 s 102788 -480 102900 240 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 403 nsew signal tristate
flabel metal2 s 105644 -480 105756 240 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 404 nsew signal tristate
flabel metal2 s 24724 -480 24836 240 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 405 nsew signal tristate
flabel metal2 s 28532 -480 28644 240 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 406 nsew signal tristate
flabel metal2 s 31388 -480 31500 240 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 407 nsew signal tristate
flabel metal2 s 34244 -480 34356 240 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 408 nsew signal tristate
flabel metal2 s 37100 -480 37212 240 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 409 nsew signal tristate
flabel metal2 s 39956 -480 40068 240 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 410 nsew signal tristate
flabel metal2 s 42812 -480 42924 240 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 411 nsew signal tristate
flabel metal2 s 14252 -480 14364 240 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 412 nsew signal input
flabel metal2 s 18060 -480 18172 240 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 413 nsew signal input
flabel metal2 s 21868 -480 21980 240 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 414 nsew signal input
flabel metal2 s 25676 -480 25788 240 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 415 nsew signal input
flabel metal2 s 9492 -480 9604 240 0 FreeSans 448 90 0 0 wbs_stb_i
port 416 nsew signal input
flabel metal2 s 10444 -480 10556 240 0 FreeSans 448 90 0 0 wbs_we_i
port 417 nsew signal input
rlabel via4 284815 173161 284815 173161 0 vdd
rlabel via4 281297 176161 281297 176161 0 vss
rlabel metal4 295652 4732 295652 4732 0 io_in[0]
rlabel metal3 289779 27636 289779 27636 0 io_in[1]
rlabel metal3 289779 49476 289779 49476 0 io_in[2]
rlabel metal3 1995 166684 1995 166684 0 io_in[30]
rlabel metal3 1995 145516 1995 145516 0 io_in[31]
rlabel metal3 1995 124292 1995 124292 0 io_in[32]
rlabel metal3 1659 103180 1659 103180 0 io_in[33]
rlabel metal3 1155 82012 1155 82012 0 io_in[34]
rlabel metal3 1799 60844 1799 60844 0 io_in[35]
rlabel metal3 1995 39676 1995 39676 0 io_in[36]
rlabel metal3 1799 18452 1799 18452 0 io_in[37]
rlabel metal3 286895 71316 286895 71316 0 io_in[3]
rlabel metal3 286895 93156 286895 93156 0 io_in[4]
rlabel metal3 286867 114996 286867 114996 0 io_in[5]
rlabel metal3 286895 136836 286895 136836 0 io_in[6]
rlabel metal3 286895 158676 286895 158676 0 io_in[7]
rlabel metal3 295701 16828 295701 16828 0 io_oeb[0]
rlabel metal3 295701 36596 295701 36596 0 io_oeb[1]
rlabel metal3 286839 64036 286839 64036 0 io_oeb[2]
rlabel metal3 1995 152572 1995 152572 0 io_oeb[30]
rlabel metal3 1659 131404 1659 131404 0 io_oeb[31]
rlabel metal3 1155 110236 1155 110236 0 io_oeb[32]
rlabel metal3 1351 89012 1351 89012 0 io_oeb[33]
rlabel metal3 1995 67900 1995 67900 0 io_oeb[34]
rlabel metal3 1995 46732 1995 46732 0 io_oeb[35]
rlabel metal3 1351 25564 1351 25564 0 io_oeb[36]
rlabel metal3 1799 4396 1799 4396 0 io_oeb[37]
rlabel metal3 286839 85876 286839 85876 0 io_oeb[3]
rlabel metal3 286839 107716 286839 107716 0 io_oeb[4]
rlabel metal3 286839 129556 286839 129556 0 io_oeb[5]
rlabel metal3 286839 151396 286839 151396 0 io_oeb[6]
rlabel metal3 286839 173236 286839 173236 0 io_oeb[7]
rlabel metal3 289779 13076 289779 13076 0 io_out[0]
rlabel metal4 293188 32452 293188 32452 0 io_out[1]
rlabel metal3 296541 49924 296541 49924 0 io_out[2]
rlabel metal3 1995 159572 1995 159572 0 io_out[30]
rlabel metal3 1995 138460 1995 138460 0 io_out[31]
rlabel metal3 1659 117292 1659 117292 0 io_out[32]
rlabel metal3 1155 96124 1155 96124 0 io_out[33]
rlabel metal3 1995 74956 1995 74956 0 io_out[34]
rlabel metal3 1799 53732 1799 53732 0 io_out[35]
rlabel metal3 1799 32620 1799 32620 0 io_out[36]
rlabel metal3 1155 11452 1155 11452 0 io_out[37]
rlabel metal3 286867 78596 286867 78596 0 io_out[3]
rlabel metal3 286867 100436 286867 100436 0 io_out[4]
rlabel metal3 286951 122276 286951 122276 0 io_out[5]
rlabel metal3 286867 144116 286867 144116 0 io_out[6]
rlabel metal3 286867 165956 286867 165956 0 io_out[7]
rlabel metal2 145908 777 145908 777 0 user_irq[0]
rlabel metal2 202244 812 202244 812 0 user_irq[1]
rlabel metal2 257908 833 257908 833 0 user_irq[2]
rlabel metal2 5852 140 5852 140 0 wb_clk_i
rlabel metal2 6580 168 6580 168 0 wb_rst_i
<< properties >>
string FIXED_BBOX 0 0 298020 298020
<< end >>
